module iCache(
  input         clock,
  input         reset,
  output        fromFetch_req_ready,
  input         fromFetch_req_valid,
  input  [63:0] fromFetch_req_bits,
  input         fromFetch_resp_ready,
  output        fromFetch_resp_valid,
  output [31:0] fromFetch_resp_bits,
  output        updateAllCachelines_ready,
  input         updateAllCachelines_fired,
  output        cachelinesUpdatesResp_ready,
  input         cachelinesUpdatesResp_fired,
  output [31:0] lowLevelMem_ARADDR,
  output        lowLevelMem_ARVALID,
  input         lowLevelMem_ARREADY,
  input  [63:0] lowLevelMem_RDATA,
  input         lowLevelMem_RLAST,
  input         lowLevelMem_RVALID,
  output        lowLevelMem_RREADY,
  output        debug_probe_arvalid_internal,
  output        debug_probe_cacheMissed,
  output        debug_probe_rready_signal,
  output        debug_probe_cacheFill_valid,
  output        debug_probe_axi_arvalid,
  output        debug_probe_axi_arready,
  output        debug_probe_req_valid,
  output [63:0] debug_probe_req_pc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [511:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] cache_address; // @[ICache.scala 83:21]
  wire [31:0] cache_instruction; // @[ICache.scala 83:21]
  wire [19:0] cache_tag; // @[ICache.scala 83:21]
  wire  cache_tag_valid; // @[ICache.scala 83:21]
  wire [5:0] cache_write_line_index; // @[ICache.scala 83:21]
  wire [511:0] cache_write_block; // @[ICache.scala 83:21]
  wire [19:0] cache_write_tag; // @[ICache.scala 83:21]
  wire  cache_write_in; // @[ICache.scala 83:21]
  wire  cache_invalidate_all; // @[ICache.scala 83:21]
  wire  cache_clock; // @[ICache.scala 83:21]
  wire  cache_reset; // @[ICache.scala 83:21]
  reg  commitFence; // @[ICache.scala 68:28]
  reg  requests_0_valid; // @[ICache.scala 75:25]
  reg [63:0] requests_0_address; // @[ICache.scala 75:25]
  reg  requests_1_valid; // @[ICache.scala 75:25]
  reg [63:0] requests_1_address; // @[ICache.scala 75:25]
  reg  requests_2_valid; // @[ICache.scala 75:25]
  reg [63:0] requests_2_address; // @[ICache.scala 75:25]
  reg  results_0_valid; // @[ICache.scala 85:24]
  reg [63:0] results_0_address; // @[ICache.scala 85:24]
  reg [31:0] results_0_instruction; // @[ICache.scala 85:24]
  reg [19:0] results_0_tag; // @[ICache.scala 85:24]
  reg  results_0_tagValid; // @[ICache.scala 85:24]
  reg  results_1_valid; // @[ICache.scala 85:24]
  reg [63:0] results_1_address; // @[ICache.scala 85:24]
  reg [31:0] results_1_instruction; // @[ICache.scala 85:24]
  reg [19:0] results_1_tag; // @[ICache.scala 85:24]
  reg  results_1_tagValid; // @[ICache.scala 85:24]
  reg  cacheFill_valid; // @[ICache.scala 99:26]
  reg [511:0] cacheFill_block; // @[ICache.scala 99:26]
  wire [51:0] _GEN_68 = {{32'd0}, results_0_tag}; // @[ICache.scala 106:96]
  wire  cacheMissed = ~(results_0_tagValid & results_0_address[63:12] == _GEN_68) & results_0_valid; // @[ICache.scala 106:119]
  reg  arvalid; // @[ICache.scala 107:33]
  reg  rready; // @[ICache.scala 107:33]
  wire [511:0] _cacheFill_block_T_1 = {lowLevelMem_RDATA,cacheFill_block[511:64]}; // @[Cat.scala 33:92]
  wire  _arvalid_T = ~rready; // @[ICache.scala 111:46]
  wire  _arvalid_T_2 = ~cacheFill_valid; // @[ICache.scala 111:57]
  wire  _arvalid_T_4 = lowLevelMem_ARVALID & lowLevelMem_ARREADY; // @[ICache.scala 112:49]
  wire  _rready_T_2 = lowLevelMem_RLAST & lowLevelMem_RREADY & lowLevelMem_RVALID; // @[ICache.scala 116:68]
  wire  _GEN_3 = _arvalid_T_2 & _rready_T_2; // @[ICache.scala 118:{26,44} 119:32]
  wire  _cacheStalled_T = ~fromFetch_resp_ready; // @[ICache.scala 140:62]
  wire  cacheStalled = cacheMissed | fromFetch_resp_valid & ~fromFetch_resp_ready; // @[ICache.scala 140:34]
  wire  _T_4 = ~cacheMissed; // @[ICache.scala 141:9]
  wire [19:0] _GEN_7 = results_1_valid ? results_1_tag : cache_tag; // @[ICache.scala 142:{35,51} 147:25]
  wire  _T_9 = cacheMissed & cacheFill_valid; // @[ICache.scala 150:26]
  wire [31:0] _GEN_10 = 4'h1 == results_0_address[5:2] ? cacheFill_block[63:32] : cacheFill_block[31:0]; // @[ICache.scala 151:{31,31}]
  wire [31:0] _GEN_11 = 4'h2 == results_0_address[5:2] ? cacheFill_block[95:64] : _GEN_10; // @[ICache.scala 151:{31,31}]
  wire [31:0] _GEN_12 = 4'h3 == results_0_address[5:2] ? cacheFill_block[127:96] : _GEN_11; // @[ICache.scala 151:{31,31}]
  wire [31:0] _GEN_13 = 4'h4 == results_0_address[5:2] ? cacheFill_block[159:128] : _GEN_12; // @[ICache.scala 151:{31,31}]
  wire [31:0] _GEN_14 = 4'h5 == results_0_address[5:2] ? cacheFill_block[191:160] : _GEN_13; // @[ICache.scala 151:{31,31}]
  wire [31:0] _GEN_15 = 4'h6 == results_0_address[5:2] ? cacheFill_block[223:192] : _GEN_14; // @[ICache.scala 151:{31,31}]
  wire [31:0] _GEN_16 = 4'h7 == results_0_address[5:2] ? cacheFill_block[255:224] : _GEN_15; // @[ICache.scala 151:{31,31}]
  wire [31:0] _GEN_17 = 4'h8 == results_0_address[5:2] ? cacheFill_block[287:256] : _GEN_16; // @[ICache.scala 151:{31,31}]
  wire [31:0] _GEN_18 = 4'h9 == results_0_address[5:2] ? cacheFill_block[319:288] : _GEN_17; // @[ICache.scala 151:{31,31}]
  wire [31:0] _GEN_19 = 4'ha == results_0_address[5:2] ? cacheFill_block[351:320] : _GEN_18; // @[ICache.scala 151:{31,31}]
  wire [31:0] _GEN_20 = 4'hb == results_0_address[5:2] ? cacheFill_block[383:352] : _GEN_19; // @[ICache.scala 151:{31,31}]
  wire [31:0] _GEN_21 = 4'hc == results_0_address[5:2] ? cacheFill_block[415:384] : _GEN_20; // @[ICache.scala 151:{31,31}]
  wire [31:0] _GEN_22 = 4'hd == results_0_address[5:2] ? cacheFill_block[447:416] : _GEN_21; // @[ICache.scala 151:{31,31}]
  wire [31:0] _GEN_23 = 4'he == results_0_address[5:2] ? cacheFill_block[479:448] : _GEN_22; // @[ICache.scala 151:{31,31}]
  wire [20:0] _GEN_26 = cacheMissed & cacheFill_valid ? results_0_address[32:12] : {{1'd0}, results_0_tag}; // @[ICache.scala 150:46 152:23 85:24]
  wire  _GEN_27 = cacheMissed & cacheFill_valid | results_0_tagValid; // @[ICache.scala 150:46 153:28 85:24]
  wire [20:0] _GEN_31 = ~cacheMissed & (fromFetch_resp_ready | commitFence) | ~results_0_valid ? {{1'd0}, _GEN_7} :
    _GEN_26; // @[ICache.scala 141:89]
  wire  _T_10 = ~results_1_valid; // @[ICache.scala 156:8]
  wire [31:0] _GEN_34 = 4'h1 == results_1_address[5:2] ? cacheFill_block[63:32] : cacheFill_block[31:0]; // @[ICache.scala 163:{35,35}]
  wire [31:0] _GEN_35 = 4'h2 == results_1_address[5:2] ? cacheFill_block[95:64] : _GEN_34; // @[ICache.scala 163:{35,35}]
  wire [31:0] _GEN_36 = 4'h3 == results_1_address[5:2] ? cacheFill_block[127:96] : _GEN_35; // @[ICache.scala 163:{35,35}]
  wire [31:0] _GEN_37 = 4'h4 == results_1_address[5:2] ? cacheFill_block[159:128] : _GEN_36; // @[ICache.scala 163:{35,35}]
  wire [31:0] _GEN_38 = 4'h5 == results_1_address[5:2] ? cacheFill_block[191:160] : _GEN_37; // @[ICache.scala 163:{35,35}]
  wire [31:0] _GEN_39 = 4'h6 == results_1_address[5:2] ? cacheFill_block[223:192] : _GEN_38; // @[ICache.scala 163:{35,35}]
  wire [31:0] _GEN_40 = 4'h7 == results_1_address[5:2] ? cacheFill_block[255:224] : _GEN_39; // @[ICache.scala 163:{35,35}]
  wire [31:0] _GEN_41 = 4'h8 == results_1_address[5:2] ? cacheFill_block[287:256] : _GEN_40; // @[ICache.scala 163:{35,35}]
  wire [31:0] _GEN_42 = 4'h9 == results_1_address[5:2] ? cacheFill_block[319:288] : _GEN_41; // @[ICache.scala 163:{35,35}]
  wire [31:0] _GEN_43 = 4'ha == results_1_address[5:2] ? cacheFill_block[351:320] : _GEN_42; // @[ICache.scala 163:{35,35}]
  wire [31:0] _GEN_44 = 4'hb == results_1_address[5:2] ? cacheFill_block[383:352] : _GEN_43; // @[ICache.scala 163:{35,35}]
  wire [31:0] _GEN_45 = 4'hc == results_1_address[5:2] ? cacheFill_block[415:384] : _GEN_44; // @[ICache.scala 163:{35,35}]
  wire [31:0] _GEN_46 = 4'hd == results_1_address[5:2] ? cacheFill_block[447:416] : _GEN_45; // @[ICache.scala 163:{35,35}]
  wire [31:0] _GEN_47 = 4'he == results_1_address[5:2] ? cacheFill_block[479:448] : _GEN_46; // @[ICache.scala 163:{35,35}]
  wire  _T_16 = ~cacheStalled; // @[ICache.scala 166:14]
  wire [20:0] _GEN_51 = _T_9 & results_0_address[31:6] == results_1_address[31:6] ? results_0_address[32:12] : {{1'd0},
    results_1_tag}; // @[ICache.scala 162:157 164:27 85:24]
  wire  _GEN_52 = _T_9 & results_0_address[31:6] == results_1_address[31:6] | results_1_tagValid; // @[ICache.scala 162:157 165:32 85:24]
  wire [20:0] _GEN_57 = ~results_1_valid ? {{1'd0}, cache_tag} : _GEN_51; // @[ICache.scala 156:34 160:27]
  wire  _GEN_59 = _T_10 & (_T_16 & requests_0_valid); // @[ICache.scala 170:34 172:31 174:31]
  wire  _requests_0_valid_T = fromFetch_req_ready & fromFetch_req_valid; // @[ICache.scala 180:52]
  wire  _T_23 = ~requests_1_valid; // @[ICache.scala 185:8]
  wire  _fromFetch_req_ready_T_1 = ~commitFence; // @[ICache.scala 194:55]
  wire  _commitFence_T_3 = requests_0_valid | requests_1_valid | requests_2_valid | results_0_valid | results_1_valid; // @[ICache.scala 200:74]
  wire [20:0] _GEN_69 = reset ? 21'h0 : _GEN_31; // @[ICache.scala 85:{24,24}]
  wire [20:0] _GEN_70 = reset ? 21'h0 : _GEN_57; // @[ICache.scala 85:{24,24}]
  iCacheRegisters #(.offset_width (4), .line_width(6)) cache ( // @[ICache.scala 83:21]
    .address(cache_address),
    .instruction(cache_instruction),
    .tag(cache_tag),
    .tag_valid(cache_tag_valid),
    .write_line_index(cache_write_line_index),
    .write_block(cache_write_block),
    .write_tag(cache_write_tag),
    .write_in(cache_write_in),
    .invalidate_all(cache_invalidate_all),
    .clock(cache_clock),
    .reset(cache_reset)
  );
  assign fromFetch_req_ready = _T_23 & ~commitFence; // @[ICache.scala 194:52]
  assign fromFetch_resp_valid = _T_4 & results_0_valid; // @[ICache.scala 192:40]
  assign fromFetch_resp_bits = results_0_instruction; // @[ICache.scala 193:23]
  assign updateAllCachelines_ready = ~commitFence; // @[ICache.scala 202:32]
  assign cachelinesUpdatesResp_ready = ~_commitFence_T_3 & commitFence; // @[ICache.scala 203:96]
  assign lowLevelMem_ARADDR = {results_0_address[31:6],6'h0}; // @[Cat.scala 33:92]
  assign lowLevelMem_ARVALID = arvalid; // @[ICache.scala 216:23]
  assign lowLevelMem_RREADY = rready; // @[ICache.scala 221:22]
  assign debug_probe_arvalid_internal = arvalid; // @[ICache.scala 123:32]
  assign debug_probe_cacheMissed = ~(results_0_tagValid & results_0_address[63:12] == _GEN_68) & results_0_valid; // @[ICache.scala 106:119]
  assign debug_probe_rready_signal = rready; // @[ICache.scala 125:32]
  assign debug_probe_cacheFill_valid = cacheFill_valid; // @[ICache.scala 126:32]
  assign debug_probe_axi_arvalid = lowLevelMem_ARVALID; // @[ICache.scala 127:32]
  assign debug_probe_axi_arready = lowLevelMem_ARREADY; // @[ICache.scala 128:32]
  assign debug_probe_req_valid = fromFetch_req_valid; // @[ICache.scala 129:32]
  assign debug_probe_req_pc = fromFetch_req_bits; // @[ICache.scala 130:32]
  assign cache_address = requests_0_address[31:0]; // @[ICache.scala 196:20]
  assign cache_write_line_index = results_0_address[11:6]; // @[ICache.scala 135:29]
  assign cache_write_block = cacheFill_block; // @[ICache.scala 133:24]
  assign cache_write_tag = results_0_address[31:12]; // @[ICache.scala 136:22]
  assign cache_write_in = cacheFill_valid; // @[ICache.scala 134:21]
  assign cache_invalidate_all = cachelinesUpdatesResp_fired; // @[ICache.scala 204:27]
  assign cache_clock = clock; // @[ICache.scala 137:18]
  assign cache_reset = reset; // @[ICache.scala 138:18]
  always @(posedge clock) begin
    if (reset) begin // @[ICache.scala 68:28]
      commitFence <= 1'h0; // @[ICache.scala 68:28]
    end else if (_fromFetch_req_ready_T_1) begin // @[ICache.scala 197:22]
      commitFence <= updateAllCachelines_fired; // @[ICache.scala 198:17]
    end else begin
      commitFence <= requests_0_valid | requests_1_valid | requests_2_valid | results_0_valid | results_1_valid | ~
        cachelinesUpdatesResp_fired; // @[ICache.scala 200:17]
    end
    if (reset) begin // @[ICache.scala 75:25]
      requests_0_valid <= 1'h0; // @[ICache.scala 75:25]
    end else if (_T_16 & _T_10 | ~requests_0_valid) begin // @[ICache.scala 177:78]
      if (requests_1_valid) begin // @[ICache.scala 178:36]
        requests_0_valid <= requests_1_valid; // @[ICache.scala 178:53]
      end else begin
        requests_0_valid <= fromFetch_req_ready & fromFetch_req_valid; // @[ICache.scala 180:28]
      end
    end
    if (reset) begin // @[ICache.scala 75:25]
      requests_0_address <= 64'h0; // @[ICache.scala 75:25]
    end else if (_T_16 & _T_10 | ~requests_0_valid) begin // @[ICache.scala 177:78]
      if (requests_1_valid) begin // @[ICache.scala 178:36]
        requests_0_address <= requests_1_address; // @[ICache.scala 178:53]
      end else begin
        requests_0_address <= fromFetch_req_bits; // @[ICache.scala 181:30]
      end
    end
    if (reset) begin // @[ICache.scala 75:25]
      requests_1_valid <= 1'h0; // @[ICache.scala 75:25]
    end else if (~requests_1_valid) begin // @[ICache.scala 185:35]
      requests_1_valid <= (cacheStalled | results_1_valid) & _requests_0_valid_T & requests_0_valid; // @[ICache.scala 186:30]
    end else begin
      requests_1_valid <= cacheStalled | results_1_valid; // @[ICache.scala 189:30]
    end
    if (reset) begin // @[ICache.scala 75:25]
      requests_1_address <= 64'h0; // @[ICache.scala 75:25]
    end else if (~requests_1_valid) begin // @[ICache.scala 185:35]
      requests_1_address <= fromFetch_req_bits; // @[ICache.scala 187:32]
    end
    if (reset) begin // @[ICache.scala 75:25]
      requests_2_valid <= 1'h0; // @[ICache.scala 75:25]
    end else begin
      requests_2_valid <= _GEN_59;
    end
    if (reset) begin // @[ICache.scala 75:25]
      requests_2_address <= 64'h0; // @[ICache.scala 75:25]
    end else if (_T_10) begin // @[ICache.scala 170:34]
      requests_2_address <= requests_0_address; // @[ICache.scala 171:25]
    end
    if (reset) begin // @[ICache.scala 85:24]
      results_0_valid <= 1'h0; // @[ICache.scala 85:24]
    end else if (~cacheMissed & (fromFetch_resp_ready | commitFence) | ~results_0_valid) begin // @[ICache.scala 141:89]
      if (results_1_valid) begin // @[ICache.scala 142:35]
        results_0_valid <= results_1_valid; // @[ICache.scala 142:51]
      end else begin
        results_0_valid <= requests_2_valid; // @[ICache.scala 144:27]
      end
    end
    if (reset) begin // @[ICache.scala 85:24]
      results_0_address <= 64'h0; // @[ICache.scala 85:24]
    end else if (~cacheMissed & (fromFetch_resp_ready | commitFence) | ~results_0_valid) begin // @[ICache.scala 141:89]
      if (results_1_valid) begin // @[ICache.scala 142:35]
        results_0_address <= results_1_address; // @[ICache.scala 142:51]
      end else begin
        results_0_address <= requests_2_address; // @[ICache.scala 145:29]
      end
    end
    if (reset) begin // @[ICache.scala 85:24]
      results_0_instruction <= 32'h0; // @[ICache.scala 85:24]
    end else if (~cacheMissed & (fromFetch_resp_ready | commitFence) | ~results_0_valid) begin // @[ICache.scala 141:89]
      if (results_1_valid) begin // @[ICache.scala 142:35]
        results_0_instruction <= results_1_instruction; // @[ICache.scala 142:51]
      end else begin
        results_0_instruction <= cache_instruction; // @[ICache.scala 146:33]
      end
    end else if (cacheMissed & cacheFill_valid) begin // @[ICache.scala 150:46]
      if (4'hf == results_0_address[5:2]) begin // @[ICache.scala 151:31]
        results_0_instruction <= cacheFill_block[511:480]; // @[ICache.scala 151:31]
      end else begin
        results_0_instruction <= _GEN_23;
      end
    end
    results_0_tag <= _GEN_69[19:0]; // @[ICache.scala 85:{24,24}]
    if (reset) begin // @[ICache.scala 85:24]
      results_0_tagValid <= 1'h0; // @[ICache.scala 85:24]
    end else if (~cacheMissed & (fromFetch_resp_ready | commitFence) | ~results_0_valid) begin // @[ICache.scala 141:89]
      if (results_1_valid) begin // @[ICache.scala 142:35]
        results_0_tagValid <= results_1_tagValid; // @[ICache.scala 142:51]
      end else begin
        results_0_tagValid <= cache_tag_valid; // @[ICache.scala 148:30]
      end
    end else begin
      results_0_tagValid <= _GEN_27;
    end
    if (reset) begin // @[ICache.scala 85:24]
      results_1_valid <= 1'h0; // @[ICache.scala 85:24]
    end else if (~results_1_valid) begin // @[ICache.scala 156:34]
      results_1_valid <= requests_2_valid & results_0_valid & (cacheMissed | _cacheStalled_T); // @[ICache.scala 157:29]
    end else if (!(_T_9 & results_0_address[31:6] == results_1_address[31:6])) begin // @[ICache.scala 162:157]
      if (~cacheStalled) begin // @[ICache.scala 166:29]
        results_1_valid <= 1'h0; // @[ICache.scala 167:29]
      end
    end
    if (reset) begin // @[ICache.scala 85:24]
      results_1_address <= 64'h0; // @[ICache.scala 85:24]
    end else if (~results_1_valid) begin // @[ICache.scala 156:34]
      results_1_address <= requests_2_address; // @[ICache.scala 158:31]
    end
    if (reset) begin // @[ICache.scala 85:24]
      results_1_instruction <= 32'h0; // @[ICache.scala 85:24]
    end else if (~results_1_valid) begin // @[ICache.scala 156:34]
      results_1_instruction <= cache_instruction; // @[ICache.scala 159:35]
    end else if (_T_9 & results_0_address[31:6] == results_1_address[31:6]) begin // @[ICache.scala 162:157]
      if (4'hf == results_1_address[5:2]) begin // @[ICache.scala 163:35]
        results_1_instruction <= cacheFill_block[511:480]; // @[ICache.scala 163:35]
      end else begin
        results_1_instruction <= _GEN_47;
      end
    end
    results_1_tag <= _GEN_70[19:0]; // @[ICache.scala 85:{24,24}]
    if (reset) begin // @[ICache.scala 85:24]
      results_1_tagValid <= 1'h0; // @[ICache.scala 85:24]
    end else if (~results_1_valid) begin // @[ICache.scala 156:34]
      results_1_tagValid <= cache_tag_valid; // @[ICache.scala 161:32]
    end else begin
      results_1_tagValid <= _GEN_52;
    end
    if (reset) begin // @[ICache.scala 99:26]
      cacheFill_valid <= 1'h0; // @[ICache.scala 99:26]
    end else begin
      cacheFill_valid <= _GEN_3;
    end
    if (reset) begin // @[ICache.scala 99:26]
      cacheFill_block <= 512'h0; // @[ICache.scala 99:26]
    end else if (lowLevelMem_RREADY & lowLevelMem_RVALID) begin // @[ICache.scala 109:50]
      cacheFill_block <= _cacheFill_block_T_1; // @[ICache.scala 109:68]
    end
    if (reset) begin // @[ICache.scala 107:33]
      arvalid <= 1'h0; // @[ICache.scala 107:33]
    end else if (~arvalid) begin // @[ICache.scala 111:18]
      arvalid <= cacheMissed & ~rready & ~cacheFill_valid; // @[ICache.scala 111:28]
    end else begin
      arvalid <= ~(lowLevelMem_ARVALID & lowLevelMem_ARREADY); // @[ICache.scala 112:24]
    end
    if (reset) begin // @[ICache.scala 107:33]
      rready <= 1'h0; // @[ICache.scala 107:33]
    end else if (_arvalid_T) begin // @[ICache.scala 115:17]
      rready <= _arvalid_T_4; // @[ICache.scala 115:26]
    end else begin
      rready <= ~(lowLevelMem_RLAST & lowLevelMem_RREADY & lowLevelMem_RVALID); // @[ICache.scala 116:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  commitFence = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  requests_0_valid = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  requests_0_address = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  requests_1_valid = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  requests_1_address = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  requests_2_valid = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  requests_2_address = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  results_0_valid = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  results_0_address = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  results_0_instruction = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  results_0_tag = _RAND_10[19:0];
  _RAND_11 = {1{`RANDOM}};
  results_0_tagValid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  results_1_valid = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  results_1_address = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  results_1_instruction = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  results_1_tag = _RAND_15[19:0];
  _RAND_16 = {1{`RANDOM}};
  results_1_tagValid = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  cacheFill_valid = _RAND_17[0:0];
  _RAND_18 = {16{`RANDOM}};
  cacheFill_block = _RAND_18[511:0];
  _RAND_19 = {1{`RANDOM}};
  arvalid = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  rready = _RAND_20[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module shiftReg(
  input   clock,
  input   reset,
  input   in,
  input   en,
  output  output_0,
  output  output_1,
  output  output_2,
  output  output_3,
  output  output_4
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  shiftregs_0; // @[fetch.scala 92:56]
  reg  shiftregs_1; // @[fetch.scala 92:56]
  reg  shiftregs_2; // @[fetch.scala 92:56]
  reg  shiftregs_3; // @[fetch.scala 92:56]
  reg  shiftregs_4; // @[fetch.scala 92:56]
  assign output_0 = shiftregs_0; // @[fetch.scala 101:54]
  assign output_1 = shiftregs_1; // @[fetch.scala 101:54]
  assign output_2 = shiftregs_2; // @[fetch.scala 101:54]
  assign output_3 = shiftregs_3; // @[fetch.scala 101:54]
  assign output_4 = shiftregs_4; // @[fetch.scala 101:54]
  always @(posedge clock) begin
    if (reset) begin // @[fetch.scala 92:56]
      shiftregs_0 <= 1'h0; // @[fetch.scala 92:56]
    end else if (en) begin // @[fetch.scala 94:14]
      shiftregs_0 <= in; // @[fetch.scala 95:20]
    end
    if (reset) begin // @[fetch.scala 92:56]
      shiftregs_1 <= 1'h0; // @[fetch.scala 92:56]
    end else if (en) begin // @[fetch.scala 94:14]
      shiftregs_1 <= shiftregs_0; // @[fetch.scala 97:22]
    end
    if (reset) begin // @[fetch.scala 92:56]
      shiftregs_2 <= 1'h0; // @[fetch.scala 92:56]
    end else if (en) begin // @[fetch.scala 94:14]
      shiftregs_2 <= shiftregs_1; // @[fetch.scala 97:22]
    end
    if (reset) begin // @[fetch.scala 92:56]
      shiftregs_3 <= 1'h0; // @[fetch.scala 92:56]
    end else if (en) begin // @[fetch.scala 94:14]
      shiftregs_3 <= shiftregs_2; // @[fetch.scala 97:22]
    end
    if (reset) begin // @[fetch.scala 92:56]
      shiftregs_4 <= 1'h0; // @[fetch.scala 92:56]
    end else if (en) begin // @[fetch.scala 94:14]
      shiftregs_4 <= shiftregs_3; // @[fetch.scala 97:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shiftregs_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  shiftregs_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  shiftregs_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  shiftregs_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  shiftregs_4 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module updateShiftReg(
  input   clock,
  input   reset,
  input   in,
  input   en,
  output  output_0,
  output  output_1,
  output  output_2,
  output  output_3,
  output  output_4,
  input   updateVals_0,
  input   updateVals_1,
  input   updateVals_2,
  input   updateVals_3,
  input   updateVals_4,
  input   update
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  shiftregs_0; // @[fetch.scala 92:56]
  reg  shiftregs_1; // @[fetch.scala 92:56]
  reg  shiftregs_2; // @[fetch.scala 92:56]
  reg  shiftregs_3; // @[fetch.scala 92:56]
  reg  shiftregs_4; // @[fetch.scala 92:56]
  assign output_0 = shiftregs_0; // @[fetch.scala 101:54]
  assign output_1 = shiftregs_1; // @[fetch.scala 101:54]
  assign output_2 = shiftregs_2; // @[fetch.scala 101:54]
  assign output_3 = shiftregs_3; // @[fetch.scala 101:54]
  assign output_4 = shiftregs_4; // @[fetch.scala 101:54]
  always @(posedge clock) begin
    if (reset) begin // @[fetch.scala 92:56]
      shiftregs_0 <= 1'h0; // @[fetch.scala 92:56]
    end else if (update) begin // @[fetch.scala 108:17]
      shiftregs_0 <= updateVals_0; // @[fetch.scala 109:48]
    end else if (en) begin // @[fetch.scala 94:14]
      shiftregs_0 <= in; // @[fetch.scala 95:20]
    end
    if (reset) begin // @[fetch.scala 92:56]
      shiftregs_1 <= 1'h0; // @[fetch.scala 92:56]
    end else if (update) begin // @[fetch.scala 108:17]
      shiftregs_1 <= updateVals_1; // @[fetch.scala 109:48]
    end else if (en) begin // @[fetch.scala 94:14]
      shiftregs_1 <= shiftregs_0; // @[fetch.scala 97:22]
    end
    if (reset) begin // @[fetch.scala 92:56]
      shiftregs_2 <= 1'h0; // @[fetch.scala 92:56]
    end else if (update) begin // @[fetch.scala 108:17]
      shiftregs_2 <= updateVals_2; // @[fetch.scala 109:48]
    end else if (en) begin // @[fetch.scala 94:14]
      shiftregs_2 <= shiftregs_1; // @[fetch.scala 97:22]
    end
    if (reset) begin // @[fetch.scala 92:56]
      shiftregs_3 <= 1'h0; // @[fetch.scala 92:56]
    end else if (update) begin // @[fetch.scala 108:17]
      shiftregs_3 <= updateVals_3; // @[fetch.scala 109:48]
    end else if (en) begin // @[fetch.scala 94:14]
      shiftregs_3 <= shiftregs_2; // @[fetch.scala 97:22]
    end
    if (reset) begin // @[fetch.scala 92:56]
      shiftregs_4 <= 1'h0; // @[fetch.scala 92:56]
    end else if (update) begin // @[fetch.scala 108:17]
      shiftregs_4 <= updateVals_4; // @[fetch.scala 109:48]
    end else if (en) begin // @[fetch.scala 94:14]
      shiftregs_4 <= shiftregs_3; // @[fetch.scala 97:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shiftregs_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  shiftregs_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  shiftregs_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  shiftregs_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  shiftregs_4 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module gshare_predictor(
  input         clock,
  input         reset,
  input         io_branchres_fired,
  input         io_branchres_branchTaken,
  input  [63:0] io_branchres_pc,
  input  [63:0] io_branchres_pcAfterBrnach,
  input  [63:0] io_curr_pc,
  output [63:0] io_next_pc,
  input         requestSent,
  input         mispredicted
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
`endif // RANDOMIZE_REG_INIT
  wire  correct_history_clock; // @[fetch.scala 123:31]
  wire  correct_history_reset; // @[fetch.scala 123:31]
  wire  correct_history_in; // @[fetch.scala 123:31]
  wire  correct_history_en; // @[fetch.scala 123:31]
  wire  correct_history_output_0; // @[fetch.scala 123:31]
  wire  correct_history_output_1; // @[fetch.scala 123:31]
  wire  correct_history_output_2; // @[fetch.scala 123:31]
  wire  correct_history_output_3; // @[fetch.scala 123:31]
  wire  correct_history_output_4; // @[fetch.scala 123:31]
  wire  predicted_history_clock; // @[fetch.scala 124:33]
  wire  predicted_history_reset; // @[fetch.scala 124:33]
  wire  predicted_history_in; // @[fetch.scala 124:33]
  wire  predicted_history_en; // @[fetch.scala 124:33]
  wire  predicted_history_output_0; // @[fetch.scala 124:33]
  wire  predicted_history_output_1; // @[fetch.scala 124:33]
  wire  predicted_history_output_2; // @[fetch.scala 124:33]
  wire  predicted_history_output_3; // @[fetch.scala 124:33]
  wire  predicted_history_output_4; // @[fetch.scala 124:33]
  wire  predicted_history_updateVals_0; // @[fetch.scala 124:33]
  wire  predicted_history_updateVals_1; // @[fetch.scala 124:33]
  wire  predicted_history_updateVals_2; // @[fetch.scala 124:33]
  wire  predicted_history_updateVals_3; // @[fetch.scala 124:33]
  wire  predicted_history_updateVals_4; // @[fetch.scala 124:33]
  wire  predicted_history_update; // @[fetch.scala 124:33]
  reg [63:0] btb [0:255]; // @[fetch.scala 148:16]
  wire  btb_io_next_pc_MPORT_en; // @[fetch.scala 148:16]
  wire [7:0] btb_io_next_pc_MPORT_addr; // @[fetch.scala 148:16]
  wire [63:0] btb_io_next_pc_MPORT_data; // @[fetch.scala 148:16]
  wire [63:0] btb_MPORT_1_data; // @[fetch.scala 148:16]
  wire [7:0] btb_MPORT_1_addr; // @[fetch.scala 148:16]
  wire  btb_MPORT_1_mask; // @[fetch.scala 148:16]
  wire  btb_MPORT_1_en; // @[fetch.scala 148:16]
  reg [1:0] counters [0:2047]; // @[fetch.scala 149:21]
  wire  counters_MPORT_2_en; // @[fetch.scala 149:21]
  wire [10:0] counters_MPORT_2_addr; // @[fetch.scala 149:21]
  wire [1:0] counters_MPORT_2_data; // @[fetch.scala 149:21]
  wire  counters_MPORT_4_en; // @[fetch.scala 149:21]
  wire [10:0] counters_MPORT_4_addr; // @[fetch.scala 149:21]
  wire [1:0] counters_MPORT_4_data; // @[fetch.scala 149:21]
  wire  counters_MPORT_5_en; // @[fetch.scala 149:21]
  wire [10:0] counters_MPORT_5_addr; // @[fetch.scala 149:21]
  wire [1:0] counters_MPORT_5_data; // @[fetch.scala 149:21]
  wire  counters_MPORT_7_en; // @[fetch.scala 149:21]
  wire [10:0] counters_MPORT_7_addr; // @[fetch.scala 149:21]
  wire [1:0] counters_MPORT_7_data; // @[fetch.scala 149:21]
  wire  counters_prediction_MPORT_en; // @[fetch.scala 149:21]
  wire [10:0] counters_prediction_MPORT_addr; // @[fetch.scala 149:21]
  wire [1:0] counters_prediction_MPORT_data; // @[fetch.scala 149:21]
  wire [1:0] counters_MPORT_3_data; // @[fetch.scala 149:21]
  wire [10:0] counters_MPORT_3_addr; // @[fetch.scala 149:21]
  wire  counters_MPORT_3_mask; // @[fetch.scala 149:21]
  wire  counters_MPORT_3_en; // @[fetch.scala 149:21]
  wire [1:0] counters_MPORT_6_data; // @[fetch.scala 149:21]
  wire [10:0] counters_MPORT_6_addr; // @[fetch.scala 149:21]
  wire  counters_MPORT_6_mask; // @[fetch.scala 149:21]
  wire  counters_MPORT_6_en; // @[fetch.scala 149:21]
  reg [53:0] tag_store [0:255]; // @[fetch.scala 151:22]
  wire  tag_store_btb_hit_MPORT_en; // @[fetch.scala 151:22]
  wire [7:0] tag_store_btb_hit_MPORT_addr; // @[fetch.scala 151:22]
  wire [53:0] tag_store_btb_hit_MPORT_data; // @[fetch.scala 151:22]
  wire [53:0] tag_store_MPORT_data; // @[fetch.scala 151:22]
  wire [7:0] tag_store_MPORT_addr; // @[fetch.scala 151:22]
  wire  tag_store_MPORT_mask; // @[fetch.scala 151:22]
  wire  tag_store_MPORT_en; // @[fetch.scala 151:22]
  wire [4:0] _counterIndex_pred_T_2 = {predicted_history_output_4,predicted_history_output_3,predicted_history_output_2,
    predicted_history_output_1,predicted_history_output_0}; // @[fetch.scala 133:178]
  wire [4:0] _counterIndex_pred_T_14 = {_counterIndex_pred_T_2[0],_counterIndex_pred_T_2[1],_counterIndex_pred_T_2[2],
    _counterIndex_pred_T_2[3],_counterIndex_pred_T_2[4]}; // @[Cat.scala 33:92]
  wire [4:0] _counterIndex_pred_T_15 = io_curr_pc[6:2] ^ _counterIndex_pred_T_14; // @[fetch.scala 133:143]
  wire [4:0] _counterIndex_train_T_2 = {correct_history_output_4,correct_history_output_3,correct_history_output_2,
    correct_history_output_1,correct_history_output_0}; // @[fetch.scala 134:187]
  wire [4:0] _counterIndex_train_T_14 = {_counterIndex_train_T_2[0],_counterIndex_train_T_2[1],_counterIndex_train_T_2[2
    ],_counterIndex_train_T_2[3],_counterIndex_train_T_2[4]}; // @[Cat.scala 33:92]
  wire [4:0] _counterIndex_train_T_15 = io_branchres_pc[6:2] ^ _counterIndex_train_T_14; // @[fetch.scala 134:154]
  wire [7:0] btb_addr = io_curr_pc[9:2]; // @[fetch.scala 142:28]
  wire [53:0] tag = io_curr_pc[63:10]; // @[fetch.scala 143:23]
  wire [7:0] result_addr = io_branchres_pc[9:2]; // @[fetch.scala 144:36]
  reg  valid_bits_0; // @[fetch.scala 150:27]
  reg  valid_bits_1; // @[fetch.scala 150:27]
  reg  valid_bits_2; // @[fetch.scala 150:27]
  reg  valid_bits_3; // @[fetch.scala 150:27]
  reg  valid_bits_4; // @[fetch.scala 150:27]
  reg  valid_bits_5; // @[fetch.scala 150:27]
  reg  valid_bits_6; // @[fetch.scala 150:27]
  reg  valid_bits_7; // @[fetch.scala 150:27]
  reg  valid_bits_8; // @[fetch.scala 150:27]
  reg  valid_bits_9; // @[fetch.scala 150:27]
  reg  valid_bits_10; // @[fetch.scala 150:27]
  reg  valid_bits_11; // @[fetch.scala 150:27]
  reg  valid_bits_12; // @[fetch.scala 150:27]
  reg  valid_bits_13; // @[fetch.scala 150:27]
  reg  valid_bits_14; // @[fetch.scala 150:27]
  reg  valid_bits_15; // @[fetch.scala 150:27]
  reg  valid_bits_16; // @[fetch.scala 150:27]
  reg  valid_bits_17; // @[fetch.scala 150:27]
  reg  valid_bits_18; // @[fetch.scala 150:27]
  reg  valid_bits_19; // @[fetch.scala 150:27]
  reg  valid_bits_20; // @[fetch.scala 150:27]
  reg  valid_bits_21; // @[fetch.scala 150:27]
  reg  valid_bits_22; // @[fetch.scala 150:27]
  reg  valid_bits_23; // @[fetch.scala 150:27]
  reg  valid_bits_24; // @[fetch.scala 150:27]
  reg  valid_bits_25; // @[fetch.scala 150:27]
  reg  valid_bits_26; // @[fetch.scala 150:27]
  reg  valid_bits_27; // @[fetch.scala 150:27]
  reg  valid_bits_28; // @[fetch.scala 150:27]
  reg  valid_bits_29; // @[fetch.scala 150:27]
  reg  valid_bits_30; // @[fetch.scala 150:27]
  reg  valid_bits_31; // @[fetch.scala 150:27]
  reg  valid_bits_32; // @[fetch.scala 150:27]
  reg  valid_bits_33; // @[fetch.scala 150:27]
  reg  valid_bits_34; // @[fetch.scala 150:27]
  reg  valid_bits_35; // @[fetch.scala 150:27]
  reg  valid_bits_36; // @[fetch.scala 150:27]
  reg  valid_bits_37; // @[fetch.scala 150:27]
  reg  valid_bits_38; // @[fetch.scala 150:27]
  reg  valid_bits_39; // @[fetch.scala 150:27]
  reg  valid_bits_40; // @[fetch.scala 150:27]
  reg  valid_bits_41; // @[fetch.scala 150:27]
  reg  valid_bits_42; // @[fetch.scala 150:27]
  reg  valid_bits_43; // @[fetch.scala 150:27]
  reg  valid_bits_44; // @[fetch.scala 150:27]
  reg  valid_bits_45; // @[fetch.scala 150:27]
  reg  valid_bits_46; // @[fetch.scala 150:27]
  reg  valid_bits_47; // @[fetch.scala 150:27]
  reg  valid_bits_48; // @[fetch.scala 150:27]
  reg  valid_bits_49; // @[fetch.scala 150:27]
  reg  valid_bits_50; // @[fetch.scala 150:27]
  reg  valid_bits_51; // @[fetch.scala 150:27]
  reg  valid_bits_52; // @[fetch.scala 150:27]
  reg  valid_bits_53; // @[fetch.scala 150:27]
  reg  valid_bits_54; // @[fetch.scala 150:27]
  reg  valid_bits_55; // @[fetch.scala 150:27]
  reg  valid_bits_56; // @[fetch.scala 150:27]
  reg  valid_bits_57; // @[fetch.scala 150:27]
  reg  valid_bits_58; // @[fetch.scala 150:27]
  reg  valid_bits_59; // @[fetch.scala 150:27]
  reg  valid_bits_60; // @[fetch.scala 150:27]
  reg  valid_bits_61; // @[fetch.scala 150:27]
  reg  valid_bits_62; // @[fetch.scala 150:27]
  reg  valid_bits_63; // @[fetch.scala 150:27]
  reg  valid_bits_64; // @[fetch.scala 150:27]
  reg  valid_bits_65; // @[fetch.scala 150:27]
  reg  valid_bits_66; // @[fetch.scala 150:27]
  reg  valid_bits_67; // @[fetch.scala 150:27]
  reg  valid_bits_68; // @[fetch.scala 150:27]
  reg  valid_bits_69; // @[fetch.scala 150:27]
  reg  valid_bits_70; // @[fetch.scala 150:27]
  reg  valid_bits_71; // @[fetch.scala 150:27]
  reg  valid_bits_72; // @[fetch.scala 150:27]
  reg  valid_bits_73; // @[fetch.scala 150:27]
  reg  valid_bits_74; // @[fetch.scala 150:27]
  reg  valid_bits_75; // @[fetch.scala 150:27]
  reg  valid_bits_76; // @[fetch.scala 150:27]
  reg  valid_bits_77; // @[fetch.scala 150:27]
  reg  valid_bits_78; // @[fetch.scala 150:27]
  reg  valid_bits_79; // @[fetch.scala 150:27]
  reg  valid_bits_80; // @[fetch.scala 150:27]
  reg  valid_bits_81; // @[fetch.scala 150:27]
  reg  valid_bits_82; // @[fetch.scala 150:27]
  reg  valid_bits_83; // @[fetch.scala 150:27]
  reg  valid_bits_84; // @[fetch.scala 150:27]
  reg  valid_bits_85; // @[fetch.scala 150:27]
  reg  valid_bits_86; // @[fetch.scala 150:27]
  reg  valid_bits_87; // @[fetch.scala 150:27]
  reg  valid_bits_88; // @[fetch.scala 150:27]
  reg  valid_bits_89; // @[fetch.scala 150:27]
  reg  valid_bits_90; // @[fetch.scala 150:27]
  reg  valid_bits_91; // @[fetch.scala 150:27]
  reg  valid_bits_92; // @[fetch.scala 150:27]
  reg  valid_bits_93; // @[fetch.scala 150:27]
  reg  valid_bits_94; // @[fetch.scala 150:27]
  reg  valid_bits_95; // @[fetch.scala 150:27]
  reg  valid_bits_96; // @[fetch.scala 150:27]
  reg  valid_bits_97; // @[fetch.scala 150:27]
  reg  valid_bits_98; // @[fetch.scala 150:27]
  reg  valid_bits_99; // @[fetch.scala 150:27]
  reg  valid_bits_100; // @[fetch.scala 150:27]
  reg  valid_bits_101; // @[fetch.scala 150:27]
  reg  valid_bits_102; // @[fetch.scala 150:27]
  reg  valid_bits_103; // @[fetch.scala 150:27]
  reg  valid_bits_104; // @[fetch.scala 150:27]
  reg  valid_bits_105; // @[fetch.scala 150:27]
  reg  valid_bits_106; // @[fetch.scala 150:27]
  reg  valid_bits_107; // @[fetch.scala 150:27]
  reg  valid_bits_108; // @[fetch.scala 150:27]
  reg  valid_bits_109; // @[fetch.scala 150:27]
  reg  valid_bits_110; // @[fetch.scala 150:27]
  reg  valid_bits_111; // @[fetch.scala 150:27]
  reg  valid_bits_112; // @[fetch.scala 150:27]
  reg  valid_bits_113; // @[fetch.scala 150:27]
  reg  valid_bits_114; // @[fetch.scala 150:27]
  reg  valid_bits_115; // @[fetch.scala 150:27]
  reg  valid_bits_116; // @[fetch.scala 150:27]
  reg  valid_bits_117; // @[fetch.scala 150:27]
  reg  valid_bits_118; // @[fetch.scala 150:27]
  reg  valid_bits_119; // @[fetch.scala 150:27]
  reg  valid_bits_120; // @[fetch.scala 150:27]
  reg  valid_bits_121; // @[fetch.scala 150:27]
  reg  valid_bits_122; // @[fetch.scala 150:27]
  reg  valid_bits_123; // @[fetch.scala 150:27]
  reg  valid_bits_124; // @[fetch.scala 150:27]
  reg  valid_bits_125; // @[fetch.scala 150:27]
  reg  valid_bits_126; // @[fetch.scala 150:27]
  reg  valid_bits_127; // @[fetch.scala 150:27]
  reg  valid_bits_128; // @[fetch.scala 150:27]
  reg  valid_bits_129; // @[fetch.scala 150:27]
  reg  valid_bits_130; // @[fetch.scala 150:27]
  reg  valid_bits_131; // @[fetch.scala 150:27]
  reg  valid_bits_132; // @[fetch.scala 150:27]
  reg  valid_bits_133; // @[fetch.scala 150:27]
  reg  valid_bits_134; // @[fetch.scala 150:27]
  reg  valid_bits_135; // @[fetch.scala 150:27]
  reg  valid_bits_136; // @[fetch.scala 150:27]
  reg  valid_bits_137; // @[fetch.scala 150:27]
  reg  valid_bits_138; // @[fetch.scala 150:27]
  reg  valid_bits_139; // @[fetch.scala 150:27]
  reg  valid_bits_140; // @[fetch.scala 150:27]
  reg  valid_bits_141; // @[fetch.scala 150:27]
  reg  valid_bits_142; // @[fetch.scala 150:27]
  reg  valid_bits_143; // @[fetch.scala 150:27]
  reg  valid_bits_144; // @[fetch.scala 150:27]
  reg  valid_bits_145; // @[fetch.scala 150:27]
  reg  valid_bits_146; // @[fetch.scala 150:27]
  reg  valid_bits_147; // @[fetch.scala 150:27]
  reg  valid_bits_148; // @[fetch.scala 150:27]
  reg  valid_bits_149; // @[fetch.scala 150:27]
  reg  valid_bits_150; // @[fetch.scala 150:27]
  reg  valid_bits_151; // @[fetch.scala 150:27]
  reg  valid_bits_152; // @[fetch.scala 150:27]
  reg  valid_bits_153; // @[fetch.scala 150:27]
  reg  valid_bits_154; // @[fetch.scala 150:27]
  reg  valid_bits_155; // @[fetch.scala 150:27]
  reg  valid_bits_156; // @[fetch.scala 150:27]
  reg  valid_bits_157; // @[fetch.scala 150:27]
  reg  valid_bits_158; // @[fetch.scala 150:27]
  reg  valid_bits_159; // @[fetch.scala 150:27]
  reg  valid_bits_160; // @[fetch.scala 150:27]
  reg  valid_bits_161; // @[fetch.scala 150:27]
  reg  valid_bits_162; // @[fetch.scala 150:27]
  reg  valid_bits_163; // @[fetch.scala 150:27]
  reg  valid_bits_164; // @[fetch.scala 150:27]
  reg  valid_bits_165; // @[fetch.scala 150:27]
  reg  valid_bits_166; // @[fetch.scala 150:27]
  reg  valid_bits_167; // @[fetch.scala 150:27]
  reg  valid_bits_168; // @[fetch.scala 150:27]
  reg  valid_bits_169; // @[fetch.scala 150:27]
  reg  valid_bits_170; // @[fetch.scala 150:27]
  reg  valid_bits_171; // @[fetch.scala 150:27]
  reg  valid_bits_172; // @[fetch.scala 150:27]
  reg  valid_bits_173; // @[fetch.scala 150:27]
  reg  valid_bits_174; // @[fetch.scala 150:27]
  reg  valid_bits_175; // @[fetch.scala 150:27]
  reg  valid_bits_176; // @[fetch.scala 150:27]
  reg  valid_bits_177; // @[fetch.scala 150:27]
  reg  valid_bits_178; // @[fetch.scala 150:27]
  reg  valid_bits_179; // @[fetch.scala 150:27]
  reg  valid_bits_180; // @[fetch.scala 150:27]
  reg  valid_bits_181; // @[fetch.scala 150:27]
  reg  valid_bits_182; // @[fetch.scala 150:27]
  reg  valid_bits_183; // @[fetch.scala 150:27]
  reg  valid_bits_184; // @[fetch.scala 150:27]
  reg  valid_bits_185; // @[fetch.scala 150:27]
  reg  valid_bits_186; // @[fetch.scala 150:27]
  reg  valid_bits_187; // @[fetch.scala 150:27]
  reg  valid_bits_188; // @[fetch.scala 150:27]
  reg  valid_bits_189; // @[fetch.scala 150:27]
  reg  valid_bits_190; // @[fetch.scala 150:27]
  reg  valid_bits_191; // @[fetch.scala 150:27]
  reg  valid_bits_192; // @[fetch.scala 150:27]
  reg  valid_bits_193; // @[fetch.scala 150:27]
  reg  valid_bits_194; // @[fetch.scala 150:27]
  reg  valid_bits_195; // @[fetch.scala 150:27]
  reg  valid_bits_196; // @[fetch.scala 150:27]
  reg  valid_bits_197; // @[fetch.scala 150:27]
  reg  valid_bits_198; // @[fetch.scala 150:27]
  reg  valid_bits_199; // @[fetch.scala 150:27]
  reg  valid_bits_200; // @[fetch.scala 150:27]
  reg  valid_bits_201; // @[fetch.scala 150:27]
  reg  valid_bits_202; // @[fetch.scala 150:27]
  reg  valid_bits_203; // @[fetch.scala 150:27]
  reg  valid_bits_204; // @[fetch.scala 150:27]
  reg  valid_bits_205; // @[fetch.scala 150:27]
  reg  valid_bits_206; // @[fetch.scala 150:27]
  reg  valid_bits_207; // @[fetch.scala 150:27]
  reg  valid_bits_208; // @[fetch.scala 150:27]
  reg  valid_bits_209; // @[fetch.scala 150:27]
  reg  valid_bits_210; // @[fetch.scala 150:27]
  reg  valid_bits_211; // @[fetch.scala 150:27]
  reg  valid_bits_212; // @[fetch.scala 150:27]
  reg  valid_bits_213; // @[fetch.scala 150:27]
  reg  valid_bits_214; // @[fetch.scala 150:27]
  reg  valid_bits_215; // @[fetch.scala 150:27]
  reg  valid_bits_216; // @[fetch.scala 150:27]
  reg  valid_bits_217; // @[fetch.scala 150:27]
  reg  valid_bits_218; // @[fetch.scala 150:27]
  reg  valid_bits_219; // @[fetch.scala 150:27]
  reg  valid_bits_220; // @[fetch.scala 150:27]
  reg  valid_bits_221; // @[fetch.scala 150:27]
  reg  valid_bits_222; // @[fetch.scala 150:27]
  reg  valid_bits_223; // @[fetch.scala 150:27]
  reg  valid_bits_224; // @[fetch.scala 150:27]
  reg  valid_bits_225; // @[fetch.scala 150:27]
  reg  valid_bits_226; // @[fetch.scala 150:27]
  reg  valid_bits_227; // @[fetch.scala 150:27]
  reg  valid_bits_228; // @[fetch.scala 150:27]
  reg  valid_bits_229; // @[fetch.scala 150:27]
  reg  valid_bits_230; // @[fetch.scala 150:27]
  reg  valid_bits_231; // @[fetch.scala 150:27]
  reg  valid_bits_232; // @[fetch.scala 150:27]
  reg  valid_bits_233; // @[fetch.scala 150:27]
  reg  valid_bits_234; // @[fetch.scala 150:27]
  reg  valid_bits_235; // @[fetch.scala 150:27]
  reg  valid_bits_236; // @[fetch.scala 150:27]
  reg  valid_bits_237; // @[fetch.scala 150:27]
  reg  valid_bits_238; // @[fetch.scala 150:27]
  reg  valid_bits_239; // @[fetch.scala 150:27]
  reg  valid_bits_240; // @[fetch.scala 150:27]
  reg  valid_bits_241; // @[fetch.scala 150:27]
  reg  valid_bits_242; // @[fetch.scala 150:27]
  reg  valid_bits_243; // @[fetch.scala 150:27]
  reg  valid_bits_244; // @[fetch.scala 150:27]
  reg  valid_bits_245; // @[fetch.scala 150:27]
  reg  valid_bits_246; // @[fetch.scala 150:27]
  reg  valid_bits_247; // @[fetch.scala 150:27]
  reg  valid_bits_248; // @[fetch.scala 150:27]
  reg  valid_bits_249; // @[fetch.scala 150:27]
  reg  valid_bits_250; // @[fetch.scala 150:27]
  reg  valid_bits_251; // @[fetch.scala 150:27]
  reg  valid_bits_252; // @[fetch.scala 150:27]
  reg  valid_bits_253; // @[fetch.scala 150:27]
  reg  valid_bits_254; // @[fetch.scala 150:27]
  reg  valid_bits_255; // @[fetch.scala 150:27]
  wire  _GEN_0 = 8'h0 == result_addr | valid_bits_0; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_1 = 8'h1 == result_addr | valid_bits_1; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_2 = 8'h2 == result_addr | valid_bits_2; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_3 = 8'h3 == result_addr | valid_bits_3; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_4 = 8'h4 == result_addr | valid_bits_4; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_5 = 8'h5 == result_addr | valid_bits_5; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_6 = 8'h6 == result_addr | valid_bits_6; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_7 = 8'h7 == result_addr | valid_bits_7; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_8 = 8'h8 == result_addr | valid_bits_8; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_9 = 8'h9 == result_addr | valid_bits_9; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_10 = 8'ha == result_addr | valid_bits_10; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_11 = 8'hb == result_addr | valid_bits_11; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_12 = 8'hc == result_addr | valid_bits_12; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_13 = 8'hd == result_addr | valid_bits_13; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_14 = 8'he == result_addr | valid_bits_14; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_15 = 8'hf == result_addr | valid_bits_15; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_16 = 8'h10 == result_addr | valid_bits_16; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_17 = 8'h11 == result_addr | valid_bits_17; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_18 = 8'h12 == result_addr | valid_bits_18; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_19 = 8'h13 == result_addr | valid_bits_19; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_20 = 8'h14 == result_addr | valid_bits_20; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_21 = 8'h15 == result_addr | valid_bits_21; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_22 = 8'h16 == result_addr | valid_bits_22; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_23 = 8'h17 == result_addr | valid_bits_23; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_24 = 8'h18 == result_addr | valid_bits_24; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_25 = 8'h19 == result_addr | valid_bits_25; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_26 = 8'h1a == result_addr | valid_bits_26; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_27 = 8'h1b == result_addr | valid_bits_27; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_28 = 8'h1c == result_addr | valid_bits_28; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_29 = 8'h1d == result_addr | valid_bits_29; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_30 = 8'h1e == result_addr | valid_bits_30; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_31 = 8'h1f == result_addr | valid_bits_31; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_32 = 8'h20 == result_addr | valid_bits_32; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_33 = 8'h21 == result_addr | valid_bits_33; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_34 = 8'h22 == result_addr | valid_bits_34; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_35 = 8'h23 == result_addr | valid_bits_35; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_36 = 8'h24 == result_addr | valid_bits_36; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_37 = 8'h25 == result_addr | valid_bits_37; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_38 = 8'h26 == result_addr | valid_bits_38; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_39 = 8'h27 == result_addr | valid_bits_39; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_40 = 8'h28 == result_addr | valid_bits_40; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_41 = 8'h29 == result_addr | valid_bits_41; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_42 = 8'h2a == result_addr | valid_bits_42; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_43 = 8'h2b == result_addr | valid_bits_43; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_44 = 8'h2c == result_addr | valid_bits_44; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_45 = 8'h2d == result_addr | valid_bits_45; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_46 = 8'h2e == result_addr | valid_bits_46; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_47 = 8'h2f == result_addr | valid_bits_47; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_48 = 8'h30 == result_addr | valid_bits_48; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_49 = 8'h31 == result_addr | valid_bits_49; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_50 = 8'h32 == result_addr | valid_bits_50; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_51 = 8'h33 == result_addr | valid_bits_51; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_52 = 8'h34 == result_addr | valid_bits_52; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_53 = 8'h35 == result_addr | valid_bits_53; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_54 = 8'h36 == result_addr | valid_bits_54; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_55 = 8'h37 == result_addr | valid_bits_55; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_56 = 8'h38 == result_addr | valid_bits_56; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_57 = 8'h39 == result_addr | valid_bits_57; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_58 = 8'h3a == result_addr | valid_bits_58; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_59 = 8'h3b == result_addr | valid_bits_59; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_60 = 8'h3c == result_addr | valid_bits_60; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_61 = 8'h3d == result_addr | valid_bits_61; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_62 = 8'h3e == result_addr | valid_bits_62; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_63 = 8'h3f == result_addr | valid_bits_63; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_64 = 8'h40 == result_addr | valid_bits_64; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_65 = 8'h41 == result_addr | valid_bits_65; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_66 = 8'h42 == result_addr | valid_bits_66; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_67 = 8'h43 == result_addr | valid_bits_67; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_68 = 8'h44 == result_addr | valid_bits_68; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_69 = 8'h45 == result_addr | valid_bits_69; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_70 = 8'h46 == result_addr | valid_bits_70; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_71 = 8'h47 == result_addr | valid_bits_71; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_72 = 8'h48 == result_addr | valid_bits_72; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_73 = 8'h49 == result_addr | valid_bits_73; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_74 = 8'h4a == result_addr | valid_bits_74; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_75 = 8'h4b == result_addr | valid_bits_75; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_76 = 8'h4c == result_addr | valid_bits_76; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_77 = 8'h4d == result_addr | valid_bits_77; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_78 = 8'h4e == result_addr | valid_bits_78; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_79 = 8'h4f == result_addr | valid_bits_79; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_80 = 8'h50 == result_addr | valid_bits_80; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_81 = 8'h51 == result_addr | valid_bits_81; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_82 = 8'h52 == result_addr | valid_bits_82; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_83 = 8'h53 == result_addr | valid_bits_83; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_84 = 8'h54 == result_addr | valid_bits_84; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_85 = 8'h55 == result_addr | valid_bits_85; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_86 = 8'h56 == result_addr | valid_bits_86; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_87 = 8'h57 == result_addr | valid_bits_87; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_88 = 8'h58 == result_addr | valid_bits_88; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_89 = 8'h59 == result_addr | valid_bits_89; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_90 = 8'h5a == result_addr | valid_bits_90; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_91 = 8'h5b == result_addr | valid_bits_91; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_92 = 8'h5c == result_addr | valid_bits_92; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_93 = 8'h5d == result_addr | valid_bits_93; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_94 = 8'h5e == result_addr | valid_bits_94; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_95 = 8'h5f == result_addr | valid_bits_95; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_96 = 8'h60 == result_addr | valid_bits_96; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_97 = 8'h61 == result_addr | valid_bits_97; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_98 = 8'h62 == result_addr | valid_bits_98; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_99 = 8'h63 == result_addr | valid_bits_99; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_100 = 8'h64 == result_addr | valid_bits_100; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_101 = 8'h65 == result_addr | valid_bits_101; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_102 = 8'h66 == result_addr | valid_bits_102; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_103 = 8'h67 == result_addr | valid_bits_103; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_104 = 8'h68 == result_addr | valid_bits_104; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_105 = 8'h69 == result_addr | valid_bits_105; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_106 = 8'h6a == result_addr | valid_bits_106; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_107 = 8'h6b == result_addr | valid_bits_107; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_108 = 8'h6c == result_addr | valid_bits_108; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_109 = 8'h6d == result_addr | valid_bits_109; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_110 = 8'h6e == result_addr | valid_bits_110; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_111 = 8'h6f == result_addr | valid_bits_111; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_112 = 8'h70 == result_addr | valid_bits_112; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_113 = 8'h71 == result_addr | valid_bits_113; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_114 = 8'h72 == result_addr | valid_bits_114; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_115 = 8'h73 == result_addr | valid_bits_115; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_116 = 8'h74 == result_addr | valid_bits_116; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_117 = 8'h75 == result_addr | valid_bits_117; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_118 = 8'h76 == result_addr | valid_bits_118; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_119 = 8'h77 == result_addr | valid_bits_119; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_120 = 8'h78 == result_addr | valid_bits_120; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_121 = 8'h79 == result_addr | valid_bits_121; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_122 = 8'h7a == result_addr | valid_bits_122; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_123 = 8'h7b == result_addr | valid_bits_123; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_124 = 8'h7c == result_addr | valid_bits_124; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_125 = 8'h7d == result_addr | valid_bits_125; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_126 = 8'h7e == result_addr | valid_bits_126; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_127 = 8'h7f == result_addr | valid_bits_127; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_128 = 8'h80 == result_addr | valid_bits_128; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_129 = 8'h81 == result_addr | valid_bits_129; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_130 = 8'h82 == result_addr | valid_bits_130; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_131 = 8'h83 == result_addr | valid_bits_131; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_132 = 8'h84 == result_addr | valid_bits_132; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_133 = 8'h85 == result_addr | valid_bits_133; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_134 = 8'h86 == result_addr | valid_bits_134; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_135 = 8'h87 == result_addr | valid_bits_135; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_136 = 8'h88 == result_addr | valid_bits_136; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_137 = 8'h89 == result_addr | valid_bits_137; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_138 = 8'h8a == result_addr | valid_bits_138; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_139 = 8'h8b == result_addr | valid_bits_139; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_140 = 8'h8c == result_addr | valid_bits_140; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_141 = 8'h8d == result_addr | valid_bits_141; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_142 = 8'h8e == result_addr | valid_bits_142; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_143 = 8'h8f == result_addr | valid_bits_143; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_144 = 8'h90 == result_addr | valid_bits_144; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_145 = 8'h91 == result_addr | valid_bits_145; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_146 = 8'h92 == result_addr | valid_bits_146; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_147 = 8'h93 == result_addr | valid_bits_147; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_148 = 8'h94 == result_addr | valid_bits_148; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_149 = 8'h95 == result_addr | valid_bits_149; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_150 = 8'h96 == result_addr | valid_bits_150; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_151 = 8'h97 == result_addr | valid_bits_151; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_152 = 8'h98 == result_addr | valid_bits_152; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_153 = 8'h99 == result_addr | valid_bits_153; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_154 = 8'h9a == result_addr | valid_bits_154; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_155 = 8'h9b == result_addr | valid_bits_155; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_156 = 8'h9c == result_addr | valid_bits_156; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_157 = 8'h9d == result_addr | valid_bits_157; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_158 = 8'h9e == result_addr | valid_bits_158; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_159 = 8'h9f == result_addr | valid_bits_159; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_160 = 8'ha0 == result_addr | valid_bits_160; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_161 = 8'ha1 == result_addr | valid_bits_161; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_162 = 8'ha2 == result_addr | valid_bits_162; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_163 = 8'ha3 == result_addr | valid_bits_163; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_164 = 8'ha4 == result_addr | valid_bits_164; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_165 = 8'ha5 == result_addr | valid_bits_165; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_166 = 8'ha6 == result_addr | valid_bits_166; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_167 = 8'ha7 == result_addr | valid_bits_167; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_168 = 8'ha8 == result_addr | valid_bits_168; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_169 = 8'ha9 == result_addr | valid_bits_169; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_170 = 8'haa == result_addr | valid_bits_170; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_171 = 8'hab == result_addr | valid_bits_171; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_172 = 8'hac == result_addr | valid_bits_172; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_173 = 8'had == result_addr | valid_bits_173; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_174 = 8'hae == result_addr | valid_bits_174; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_175 = 8'haf == result_addr | valid_bits_175; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_176 = 8'hb0 == result_addr | valid_bits_176; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_177 = 8'hb1 == result_addr | valid_bits_177; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_178 = 8'hb2 == result_addr | valid_bits_178; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_179 = 8'hb3 == result_addr | valid_bits_179; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_180 = 8'hb4 == result_addr | valid_bits_180; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_181 = 8'hb5 == result_addr | valid_bits_181; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_182 = 8'hb6 == result_addr | valid_bits_182; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_183 = 8'hb7 == result_addr | valid_bits_183; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_184 = 8'hb8 == result_addr | valid_bits_184; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_185 = 8'hb9 == result_addr | valid_bits_185; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_186 = 8'hba == result_addr | valid_bits_186; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_187 = 8'hbb == result_addr | valid_bits_187; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_188 = 8'hbc == result_addr | valid_bits_188; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_189 = 8'hbd == result_addr | valid_bits_189; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_190 = 8'hbe == result_addr | valid_bits_190; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_191 = 8'hbf == result_addr | valid_bits_191; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_192 = 8'hc0 == result_addr | valid_bits_192; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_193 = 8'hc1 == result_addr | valid_bits_193; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_194 = 8'hc2 == result_addr | valid_bits_194; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_195 = 8'hc3 == result_addr | valid_bits_195; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_196 = 8'hc4 == result_addr | valid_bits_196; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_197 = 8'hc5 == result_addr | valid_bits_197; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_198 = 8'hc6 == result_addr | valid_bits_198; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_199 = 8'hc7 == result_addr | valid_bits_199; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_200 = 8'hc8 == result_addr | valid_bits_200; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_201 = 8'hc9 == result_addr | valid_bits_201; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_202 = 8'hca == result_addr | valid_bits_202; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_203 = 8'hcb == result_addr | valid_bits_203; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_204 = 8'hcc == result_addr | valid_bits_204; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_205 = 8'hcd == result_addr | valid_bits_205; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_206 = 8'hce == result_addr | valid_bits_206; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_207 = 8'hcf == result_addr | valid_bits_207; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_208 = 8'hd0 == result_addr | valid_bits_208; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_209 = 8'hd1 == result_addr | valid_bits_209; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_210 = 8'hd2 == result_addr | valid_bits_210; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_211 = 8'hd3 == result_addr | valid_bits_211; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_212 = 8'hd4 == result_addr | valid_bits_212; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_213 = 8'hd5 == result_addr | valid_bits_213; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_214 = 8'hd6 == result_addr | valid_bits_214; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_215 = 8'hd7 == result_addr | valid_bits_215; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_216 = 8'hd8 == result_addr | valid_bits_216; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_217 = 8'hd9 == result_addr | valid_bits_217; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_218 = 8'hda == result_addr | valid_bits_218; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_219 = 8'hdb == result_addr | valid_bits_219; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_220 = 8'hdc == result_addr | valid_bits_220; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_221 = 8'hdd == result_addr | valid_bits_221; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_222 = 8'hde == result_addr | valid_bits_222; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_223 = 8'hdf == result_addr | valid_bits_223; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_224 = 8'he0 == result_addr | valid_bits_224; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_225 = 8'he1 == result_addr | valid_bits_225; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_226 = 8'he2 == result_addr | valid_bits_226; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_227 = 8'he3 == result_addr | valid_bits_227; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_228 = 8'he4 == result_addr | valid_bits_228; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_229 = 8'he5 == result_addr | valid_bits_229; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_230 = 8'he6 == result_addr | valid_bits_230; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_231 = 8'he7 == result_addr | valid_bits_231; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_232 = 8'he8 == result_addr | valid_bits_232; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_233 = 8'he9 == result_addr | valid_bits_233; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_234 = 8'hea == result_addr | valid_bits_234; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_235 = 8'heb == result_addr | valid_bits_235; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_236 = 8'hec == result_addr | valid_bits_236; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_237 = 8'hed == result_addr | valid_bits_237; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_238 = 8'hee == result_addr | valid_bits_238; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_239 = 8'hef == result_addr | valid_bits_239; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_240 = 8'hf0 == result_addr | valid_bits_240; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_241 = 8'hf1 == result_addr | valid_bits_241; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_242 = 8'hf2 == result_addr | valid_bits_242; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_243 = 8'hf3 == result_addr | valid_bits_243; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_244 = 8'hf4 == result_addr | valid_bits_244; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_245 = 8'hf5 == result_addr | valid_bits_245; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_246 = 8'hf6 == result_addr | valid_bits_246; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_247 = 8'hf7 == result_addr | valid_bits_247; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_248 = 8'hf8 == result_addr | valid_bits_248; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_249 = 8'hf9 == result_addr | valid_bits_249; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_250 = 8'hfa == result_addr | valid_bits_250; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_251 = 8'hfb == result_addr | valid_bits_251; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_252 = 8'hfc == result_addr | valid_bits_252; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_253 = 8'hfd == result_addr | valid_bits_253; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_254 = 8'hfe == result_addr | valid_bits_254; // @[fetch.scala 150:27 156:{31,31}]
  wire  _GEN_255 = 8'hff == result_addr | valid_bits_255; // @[fetch.scala 150:27 156:{31,31}]
  wire  _T_1 = ~(counters_MPORT_2_data == 2'h3); // @[fetch.scala 161:14]
  wire  _T_5 = ~(counters_MPORT_5_data == 2'h0); // @[fetch.scala 165:14]
  wire  _GEN_271 = io_branchres_branchTaken & _T_1; // @[fetch.scala 149:21 160:37]
  wire  _GEN_276 = io_branchres_branchTaken ? 1'h0 : 1'h1; // @[fetch.scala 149:21 160:37 165:24]
  wire  _GEN_279 = io_branchres_branchTaken ? 1'h0 : _T_5; // @[fetch.scala 149:21 160:37]
  wire  _GEN_1351 = 8'h1 == btb_addr ? valid_bits_1 : valid_bits_0; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1352 = 8'h2 == btb_addr ? valid_bits_2 : _GEN_1351; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1353 = 8'h3 == btb_addr ? valid_bits_3 : _GEN_1352; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1354 = 8'h4 == btb_addr ? valid_bits_4 : _GEN_1353; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1355 = 8'h5 == btb_addr ? valid_bits_5 : _GEN_1354; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1356 = 8'h6 == btb_addr ? valid_bits_6 : _GEN_1355; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1357 = 8'h7 == btb_addr ? valid_bits_7 : _GEN_1356; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1358 = 8'h8 == btb_addr ? valid_bits_8 : _GEN_1357; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1359 = 8'h9 == btb_addr ? valid_bits_9 : _GEN_1358; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1360 = 8'ha == btb_addr ? valid_bits_10 : _GEN_1359; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1361 = 8'hb == btb_addr ? valid_bits_11 : _GEN_1360; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1362 = 8'hc == btb_addr ? valid_bits_12 : _GEN_1361; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1363 = 8'hd == btb_addr ? valid_bits_13 : _GEN_1362; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1364 = 8'he == btb_addr ? valid_bits_14 : _GEN_1363; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1365 = 8'hf == btb_addr ? valid_bits_15 : _GEN_1364; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1366 = 8'h10 == btb_addr ? valid_bits_16 : _GEN_1365; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1367 = 8'h11 == btb_addr ? valid_bits_17 : _GEN_1366; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1368 = 8'h12 == btb_addr ? valid_bits_18 : _GEN_1367; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1369 = 8'h13 == btb_addr ? valid_bits_19 : _GEN_1368; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1370 = 8'h14 == btb_addr ? valid_bits_20 : _GEN_1369; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1371 = 8'h15 == btb_addr ? valid_bits_21 : _GEN_1370; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1372 = 8'h16 == btb_addr ? valid_bits_22 : _GEN_1371; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1373 = 8'h17 == btb_addr ? valid_bits_23 : _GEN_1372; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1374 = 8'h18 == btb_addr ? valid_bits_24 : _GEN_1373; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1375 = 8'h19 == btb_addr ? valid_bits_25 : _GEN_1374; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1376 = 8'h1a == btb_addr ? valid_bits_26 : _GEN_1375; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1377 = 8'h1b == btb_addr ? valid_bits_27 : _GEN_1376; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1378 = 8'h1c == btb_addr ? valid_bits_28 : _GEN_1377; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1379 = 8'h1d == btb_addr ? valid_bits_29 : _GEN_1378; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1380 = 8'h1e == btb_addr ? valid_bits_30 : _GEN_1379; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1381 = 8'h1f == btb_addr ? valid_bits_31 : _GEN_1380; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1382 = 8'h20 == btb_addr ? valid_bits_32 : _GEN_1381; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1383 = 8'h21 == btb_addr ? valid_bits_33 : _GEN_1382; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1384 = 8'h22 == btb_addr ? valid_bits_34 : _GEN_1383; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1385 = 8'h23 == btb_addr ? valid_bits_35 : _GEN_1384; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1386 = 8'h24 == btb_addr ? valid_bits_36 : _GEN_1385; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1387 = 8'h25 == btb_addr ? valid_bits_37 : _GEN_1386; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1388 = 8'h26 == btb_addr ? valid_bits_38 : _GEN_1387; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1389 = 8'h27 == btb_addr ? valid_bits_39 : _GEN_1388; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1390 = 8'h28 == btb_addr ? valid_bits_40 : _GEN_1389; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1391 = 8'h29 == btb_addr ? valid_bits_41 : _GEN_1390; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1392 = 8'h2a == btb_addr ? valid_bits_42 : _GEN_1391; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1393 = 8'h2b == btb_addr ? valid_bits_43 : _GEN_1392; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1394 = 8'h2c == btb_addr ? valid_bits_44 : _GEN_1393; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1395 = 8'h2d == btb_addr ? valid_bits_45 : _GEN_1394; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1396 = 8'h2e == btb_addr ? valid_bits_46 : _GEN_1395; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1397 = 8'h2f == btb_addr ? valid_bits_47 : _GEN_1396; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1398 = 8'h30 == btb_addr ? valid_bits_48 : _GEN_1397; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1399 = 8'h31 == btb_addr ? valid_bits_49 : _GEN_1398; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1400 = 8'h32 == btb_addr ? valid_bits_50 : _GEN_1399; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1401 = 8'h33 == btb_addr ? valid_bits_51 : _GEN_1400; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1402 = 8'h34 == btb_addr ? valid_bits_52 : _GEN_1401; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1403 = 8'h35 == btb_addr ? valid_bits_53 : _GEN_1402; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1404 = 8'h36 == btb_addr ? valid_bits_54 : _GEN_1403; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1405 = 8'h37 == btb_addr ? valid_bits_55 : _GEN_1404; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1406 = 8'h38 == btb_addr ? valid_bits_56 : _GEN_1405; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1407 = 8'h39 == btb_addr ? valid_bits_57 : _GEN_1406; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1408 = 8'h3a == btb_addr ? valid_bits_58 : _GEN_1407; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1409 = 8'h3b == btb_addr ? valid_bits_59 : _GEN_1408; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1410 = 8'h3c == btb_addr ? valid_bits_60 : _GEN_1409; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1411 = 8'h3d == btb_addr ? valid_bits_61 : _GEN_1410; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1412 = 8'h3e == btb_addr ? valid_bits_62 : _GEN_1411; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1413 = 8'h3f == btb_addr ? valid_bits_63 : _GEN_1412; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1414 = 8'h40 == btb_addr ? valid_bits_64 : _GEN_1413; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1415 = 8'h41 == btb_addr ? valid_bits_65 : _GEN_1414; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1416 = 8'h42 == btb_addr ? valid_bits_66 : _GEN_1415; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1417 = 8'h43 == btb_addr ? valid_bits_67 : _GEN_1416; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1418 = 8'h44 == btb_addr ? valid_bits_68 : _GEN_1417; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1419 = 8'h45 == btb_addr ? valid_bits_69 : _GEN_1418; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1420 = 8'h46 == btb_addr ? valid_bits_70 : _GEN_1419; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1421 = 8'h47 == btb_addr ? valid_bits_71 : _GEN_1420; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1422 = 8'h48 == btb_addr ? valid_bits_72 : _GEN_1421; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1423 = 8'h49 == btb_addr ? valid_bits_73 : _GEN_1422; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1424 = 8'h4a == btb_addr ? valid_bits_74 : _GEN_1423; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1425 = 8'h4b == btb_addr ? valid_bits_75 : _GEN_1424; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1426 = 8'h4c == btb_addr ? valid_bits_76 : _GEN_1425; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1427 = 8'h4d == btb_addr ? valid_bits_77 : _GEN_1426; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1428 = 8'h4e == btb_addr ? valid_bits_78 : _GEN_1427; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1429 = 8'h4f == btb_addr ? valid_bits_79 : _GEN_1428; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1430 = 8'h50 == btb_addr ? valid_bits_80 : _GEN_1429; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1431 = 8'h51 == btb_addr ? valid_bits_81 : _GEN_1430; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1432 = 8'h52 == btb_addr ? valid_bits_82 : _GEN_1431; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1433 = 8'h53 == btb_addr ? valid_bits_83 : _GEN_1432; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1434 = 8'h54 == btb_addr ? valid_bits_84 : _GEN_1433; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1435 = 8'h55 == btb_addr ? valid_bits_85 : _GEN_1434; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1436 = 8'h56 == btb_addr ? valid_bits_86 : _GEN_1435; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1437 = 8'h57 == btb_addr ? valid_bits_87 : _GEN_1436; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1438 = 8'h58 == btb_addr ? valid_bits_88 : _GEN_1437; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1439 = 8'h59 == btb_addr ? valid_bits_89 : _GEN_1438; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1440 = 8'h5a == btb_addr ? valid_bits_90 : _GEN_1439; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1441 = 8'h5b == btb_addr ? valid_bits_91 : _GEN_1440; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1442 = 8'h5c == btb_addr ? valid_bits_92 : _GEN_1441; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1443 = 8'h5d == btb_addr ? valid_bits_93 : _GEN_1442; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1444 = 8'h5e == btb_addr ? valid_bits_94 : _GEN_1443; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1445 = 8'h5f == btb_addr ? valid_bits_95 : _GEN_1444; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1446 = 8'h60 == btb_addr ? valid_bits_96 : _GEN_1445; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1447 = 8'h61 == btb_addr ? valid_bits_97 : _GEN_1446; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1448 = 8'h62 == btb_addr ? valid_bits_98 : _GEN_1447; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1449 = 8'h63 == btb_addr ? valid_bits_99 : _GEN_1448; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1450 = 8'h64 == btb_addr ? valid_bits_100 : _GEN_1449; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1451 = 8'h65 == btb_addr ? valid_bits_101 : _GEN_1450; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1452 = 8'h66 == btb_addr ? valid_bits_102 : _GEN_1451; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1453 = 8'h67 == btb_addr ? valid_bits_103 : _GEN_1452; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1454 = 8'h68 == btb_addr ? valid_bits_104 : _GEN_1453; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1455 = 8'h69 == btb_addr ? valid_bits_105 : _GEN_1454; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1456 = 8'h6a == btb_addr ? valid_bits_106 : _GEN_1455; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1457 = 8'h6b == btb_addr ? valid_bits_107 : _GEN_1456; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1458 = 8'h6c == btb_addr ? valid_bits_108 : _GEN_1457; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1459 = 8'h6d == btb_addr ? valid_bits_109 : _GEN_1458; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1460 = 8'h6e == btb_addr ? valid_bits_110 : _GEN_1459; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1461 = 8'h6f == btb_addr ? valid_bits_111 : _GEN_1460; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1462 = 8'h70 == btb_addr ? valid_bits_112 : _GEN_1461; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1463 = 8'h71 == btb_addr ? valid_bits_113 : _GEN_1462; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1464 = 8'h72 == btb_addr ? valid_bits_114 : _GEN_1463; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1465 = 8'h73 == btb_addr ? valid_bits_115 : _GEN_1464; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1466 = 8'h74 == btb_addr ? valid_bits_116 : _GEN_1465; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1467 = 8'h75 == btb_addr ? valid_bits_117 : _GEN_1466; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1468 = 8'h76 == btb_addr ? valid_bits_118 : _GEN_1467; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1469 = 8'h77 == btb_addr ? valid_bits_119 : _GEN_1468; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1470 = 8'h78 == btb_addr ? valid_bits_120 : _GEN_1469; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1471 = 8'h79 == btb_addr ? valid_bits_121 : _GEN_1470; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1472 = 8'h7a == btb_addr ? valid_bits_122 : _GEN_1471; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1473 = 8'h7b == btb_addr ? valid_bits_123 : _GEN_1472; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1474 = 8'h7c == btb_addr ? valid_bits_124 : _GEN_1473; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1475 = 8'h7d == btb_addr ? valid_bits_125 : _GEN_1474; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1476 = 8'h7e == btb_addr ? valid_bits_126 : _GEN_1475; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1477 = 8'h7f == btb_addr ? valid_bits_127 : _GEN_1476; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1478 = 8'h80 == btb_addr ? valid_bits_128 : _GEN_1477; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1479 = 8'h81 == btb_addr ? valid_bits_129 : _GEN_1478; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1480 = 8'h82 == btb_addr ? valid_bits_130 : _GEN_1479; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1481 = 8'h83 == btb_addr ? valid_bits_131 : _GEN_1480; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1482 = 8'h84 == btb_addr ? valid_bits_132 : _GEN_1481; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1483 = 8'h85 == btb_addr ? valid_bits_133 : _GEN_1482; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1484 = 8'h86 == btb_addr ? valid_bits_134 : _GEN_1483; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1485 = 8'h87 == btb_addr ? valid_bits_135 : _GEN_1484; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1486 = 8'h88 == btb_addr ? valid_bits_136 : _GEN_1485; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1487 = 8'h89 == btb_addr ? valid_bits_137 : _GEN_1486; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1488 = 8'h8a == btb_addr ? valid_bits_138 : _GEN_1487; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1489 = 8'h8b == btb_addr ? valid_bits_139 : _GEN_1488; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1490 = 8'h8c == btb_addr ? valid_bits_140 : _GEN_1489; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1491 = 8'h8d == btb_addr ? valid_bits_141 : _GEN_1490; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1492 = 8'h8e == btb_addr ? valid_bits_142 : _GEN_1491; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1493 = 8'h8f == btb_addr ? valid_bits_143 : _GEN_1492; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1494 = 8'h90 == btb_addr ? valid_bits_144 : _GEN_1493; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1495 = 8'h91 == btb_addr ? valid_bits_145 : _GEN_1494; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1496 = 8'h92 == btb_addr ? valid_bits_146 : _GEN_1495; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1497 = 8'h93 == btb_addr ? valid_bits_147 : _GEN_1496; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1498 = 8'h94 == btb_addr ? valid_bits_148 : _GEN_1497; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1499 = 8'h95 == btb_addr ? valid_bits_149 : _GEN_1498; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1500 = 8'h96 == btb_addr ? valid_bits_150 : _GEN_1499; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1501 = 8'h97 == btb_addr ? valid_bits_151 : _GEN_1500; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1502 = 8'h98 == btb_addr ? valid_bits_152 : _GEN_1501; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1503 = 8'h99 == btb_addr ? valid_bits_153 : _GEN_1502; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1504 = 8'h9a == btb_addr ? valid_bits_154 : _GEN_1503; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1505 = 8'h9b == btb_addr ? valid_bits_155 : _GEN_1504; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1506 = 8'h9c == btb_addr ? valid_bits_156 : _GEN_1505; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1507 = 8'h9d == btb_addr ? valid_bits_157 : _GEN_1506; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1508 = 8'h9e == btb_addr ? valid_bits_158 : _GEN_1507; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1509 = 8'h9f == btb_addr ? valid_bits_159 : _GEN_1508; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1510 = 8'ha0 == btb_addr ? valid_bits_160 : _GEN_1509; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1511 = 8'ha1 == btb_addr ? valid_bits_161 : _GEN_1510; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1512 = 8'ha2 == btb_addr ? valid_bits_162 : _GEN_1511; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1513 = 8'ha3 == btb_addr ? valid_bits_163 : _GEN_1512; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1514 = 8'ha4 == btb_addr ? valid_bits_164 : _GEN_1513; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1515 = 8'ha5 == btb_addr ? valid_bits_165 : _GEN_1514; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1516 = 8'ha6 == btb_addr ? valid_bits_166 : _GEN_1515; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1517 = 8'ha7 == btb_addr ? valid_bits_167 : _GEN_1516; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1518 = 8'ha8 == btb_addr ? valid_bits_168 : _GEN_1517; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1519 = 8'ha9 == btb_addr ? valid_bits_169 : _GEN_1518; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1520 = 8'haa == btb_addr ? valid_bits_170 : _GEN_1519; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1521 = 8'hab == btb_addr ? valid_bits_171 : _GEN_1520; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1522 = 8'hac == btb_addr ? valid_bits_172 : _GEN_1521; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1523 = 8'had == btb_addr ? valid_bits_173 : _GEN_1522; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1524 = 8'hae == btb_addr ? valid_bits_174 : _GEN_1523; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1525 = 8'haf == btb_addr ? valid_bits_175 : _GEN_1524; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1526 = 8'hb0 == btb_addr ? valid_bits_176 : _GEN_1525; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1527 = 8'hb1 == btb_addr ? valid_bits_177 : _GEN_1526; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1528 = 8'hb2 == btb_addr ? valid_bits_178 : _GEN_1527; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1529 = 8'hb3 == btb_addr ? valid_bits_179 : _GEN_1528; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1530 = 8'hb4 == btb_addr ? valid_bits_180 : _GEN_1529; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1531 = 8'hb5 == btb_addr ? valid_bits_181 : _GEN_1530; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1532 = 8'hb6 == btb_addr ? valid_bits_182 : _GEN_1531; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1533 = 8'hb7 == btb_addr ? valid_bits_183 : _GEN_1532; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1534 = 8'hb8 == btb_addr ? valid_bits_184 : _GEN_1533; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1535 = 8'hb9 == btb_addr ? valid_bits_185 : _GEN_1534; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1536 = 8'hba == btb_addr ? valid_bits_186 : _GEN_1535; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1537 = 8'hbb == btb_addr ? valid_bits_187 : _GEN_1536; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1538 = 8'hbc == btb_addr ? valid_bits_188 : _GEN_1537; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1539 = 8'hbd == btb_addr ? valid_bits_189 : _GEN_1538; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1540 = 8'hbe == btb_addr ? valid_bits_190 : _GEN_1539; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1541 = 8'hbf == btb_addr ? valid_bits_191 : _GEN_1540; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1542 = 8'hc0 == btb_addr ? valid_bits_192 : _GEN_1541; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1543 = 8'hc1 == btb_addr ? valid_bits_193 : _GEN_1542; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1544 = 8'hc2 == btb_addr ? valid_bits_194 : _GEN_1543; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1545 = 8'hc3 == btb_addr ? valid_bits_195 : _GEN_1544; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1546 = 8'hc4 == btb_addr ? valid_bits_196 : _GEN_1545; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1547 = 8'hc5 == btb_addr ? valid_bits_197 : _GEN_1546; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1548 = 8'hc6 == btb_addr ? valid_bits_198 : _GEN_1547; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1549 = 8'hc7 == btb_addr ? valid_bits_199 : _GEN_1548; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1550 = 8'hc8 == btb_addr ? valid_bits_200 : _GEN_1549; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1551 = 8'hc9 == btb_addr ? valid_bits_201 : _GEN_1550; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1552 = 8'hca == btb_addr ? valid_bits_202 : _GEN_1551; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1553 = 8'hcb == btb_addr ? valid_bits_203 : _GEN_1552; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1554 = 8'hcc == btb_addr ? valid_bits_204 : _GEN_1553; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1555 = 8'hcd == btb_addr ? valid_bits_205 : _GEN_1554; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1556 = 8'hce == btb_addr ? valid_bits_206 : _GEN_1555; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1557 = 8'hcf == btb_addr ? valid_bits_207 : _GEN_1556; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1558 = 8'hd0 == btb_addr ? valid_bits_208 : _GEN_1557; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1559 = 8'hd1 == btb_addr ? valid_bits_209 : _GEN_1558; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1560 = 8'hd2 == btb_addr ? valid_bits_210 : _GEN_1559; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1561 = 8'hd3 == btb_addr ? valid_bits_211 : _GEN_1560; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1562 = 8'hd4 == btb_addr ? valid_bits_212 : _GEN_1561; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1563 = 8'hd5 == btb_addr ? valid_bits_213 : _GEN_1562; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1564 = 8'hd6 == btb_addr ? valid_bits_214 : _GEN_1563; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1565 = 8'hd7 == btb_addr ? valid_bits_215 : _GEN_1564; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1566 = 8'hd8 == btb_addr ? valid_bits_216 : _GEN_1565; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1567 = 8'hd9 == btb_addr ? valid_bits_217 : _GEN_1566; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1568 = 8'hda == btb_addr ? valid_bits_218 : _GEN_1567; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1569 = 8'hdb == btb_addr ? valid_bits_219 : _GEN_1568; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1570 = 8'hdc == btb_addr ? valid_bits_220 : _GEN_1569; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1571 = 8'hdd == btb_addr ? valid_bits_221 : _GEN_1570; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1572 = 8'hde == btb_addr ? valid_bits_222 : _GEN_1571; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1573 = 8'hdf == btb_addr ? valid_bits_223 : _GEN_1572; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1574 = 8'he0 == btb_addr ? valid_bits_224 : _GEN_1573; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1575 = 8'he1 == btb_addr ? valid_bits_225 : _GEN_1574; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1576 = 8'he2 == btb_addr ? valid_bits_226 : _GEN_1575; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1577 = 8'he3 == btb_addr ? valid_bits_227 : _GEN_1576; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1578 = 8'he4 == btb_addr ? valid_bits_228 : _GEN_1577; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1579 = 8'he5 == btb_addr ? valid_bits_229 : _GEN_1578; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1580 = 8'he6 == btb_addr ? valid_bits_230 : _GEN_1579; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1581 = 8'he7 == btb_addr ? valid_bits_231 : _GEN_1580; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1582 = 8'he8 == btb_addr ? valid_bits_232 : _GEN_1581; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1583 = 8'he9 == btb_addr ? valid_bits_233 : _GEN_1582; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1584 = 8'hea == btb_addr ? valid_bits_234 : _GEN_1583; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1585 = 8'heb == btb_addr ? valid_bits_235 : _GEN_1584; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1586 = 8'hec == btb_addr ? valid_bits_236 : _GEN_1585; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1587 = 8'hed == btb_addr ? valid_bits_237 : _GEN_1586; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1588 = 8'hee == btb_addr ? valid_bits_238 : _GEN_1587; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1589 = 8'hef == btb_addr ? valid_bits_239 : _GEN_1588; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1590 = 8'hf0 == btb_addr ? valid_bits_240 : _GEN_1589; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1591 = 8'hf1 == btb_addr ? valid_bits_241 : _GEN_1590; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1592 = 8'hf2 == btb_addr ? valid_bits_242 : _GEN_1591; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1593 = 8'hf3 == btb_addr ? valid_bits_243 : _GEN_1592; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1594 = 8'hf4 == btb_addr ? valid_bits_244 : _GEN_1593; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1595 = 8'hf5 == btb_addr ? valid_bits_245 : _GEN_1594; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1596 = 8'hf6 == btb_addr ? valid_bits_246 : _GEN_1595; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1597 = 8'hf7 == btb_addr ? valid_bits_247 : _GEN_1596; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1598 = 8'hf8 == btb_addr ? valid_bits_248 : _GEN_1597; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1599 = 8'hf9 == btb_addr ? valid_bits_249 : _GEN_1598; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1600 = 8'hfa == btb_addr ? valid_bits_250 : _GEN_1599; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1601 = 8'hfb == btb_addr ? valid_bits_251 : _GEN_1600; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1602 = 8'hfc == btb_addr ? valid_bits_252 : _GEN_1601; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1603 = 8'hfd == btb_addr ? valid_bits_253 : _GEN_1602; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1604 = 8'hfe == btb_addr ? valid_bits_254 : _GEN_1603; // @[fetch.scala 176:{37,37}]
  wire  _GEN_1605 = 8'hff == btb_addr ? valid_bits_255 : _GEN_1604; // @[fetch.scala 176:{37,37}]
  wire  btb_hit = _GEN_1605 & tag_store_btb_hit_MPORT_data == tag; // @[fetch.scala 176:44]
  wire  prediction = counters_prediction_MPORT_data[1]; // @[fetch.scala 177:47]
  wire [63:0] _io_next_pc_T_2 = io_curr_pc + 64'h4; // @[fetch.scala 182:70]
  wire  _GEN_1606 = correct_history_en ? io_branchres_branchTaken : correct_history_output_0; // @[fetch.scala 187:29 188:39 194:41]
  wire  _GEN_1607 = correct_history_output_1; // @[fetch.scala 187:29 190:41 194:41]
  wire  _GEN_1608 = correct_history_output_2; // @[fetch.scala 187:29 190:41 194:41]
  wire  _GEN_1609 = correct_history_output_3; // @[fetch.scala 187:29 190:41 194:41]
  wire  _GEN_1610 = correct_history_output_4; // @[fetch.scala 187:29 190:41 194:41]
  shiftReg correct_history ( // @[fetch.scala 123:31]
    .clock(correct_history_clock),
    .reset(correct_history_reset),
    .in(correct_history_in),
    .en(correct_history_en),
    .output_0(correct_history_output_0),
    .output_1(correct_history_output_1),
    .output_2(correct_history_output_2),
    .output_3(correct_history_output_3),
    .output_4(correct_history_output_4)
  );
  updateShiftReg predicted_history ( // @[fetch.scala 124:33]
    .clock(predicted_history_clock),
    .reset(predicted_history_reset),
    .in(predicted_history_in),
    .en(predicted_history_en),
    .output_0(predicted_history_output_0),
    .output_1(predicted_history_output_1),
    .output_2(predicted_history_output_2),
    .output_3(predicted_history_output_3),
    .output_4(predicted_history_output_4),
    .updateVals_0(predicted_history_updateVals_0),
    .updateVals_1(predicted_history_updateVals_1),
    .updateVals_2(predicted_history_updateVals_2),
    .updateVals_3(predicted_history_updateVals_3),
    .updateVals_4(predicted_history_updateVals_4),
    .update(predicted_history_update)
  );
  assign btb_io_next_pc_MPORT_en = 1'h1;
  assign btb_io_next_pc_MPORT_addr = io_curr_pc[9:2];
  assign btb_io_next_pc_MPORT_data = btb[btb_io_next_pc_MPORT_addr]; // @[fetch.scala 148:16]
  assign btb_MPORT_1_data = io_branchres_pcAfterBrnach;
  assign btb_MPORT_1_addr = io_branchres_pc[9:2];
  assign btb_MPORT_1_mask = 1'h1;
  assign btb_MPORT_1_en = io_branchres_fired;
  assign counters_MPORT_2_en = io_branchres_fired & io_branchres_branchTaken;
  assign counters_MPORT_2_addr = {io_branchres_pc[7:2],_counterIndex_train_T_15};
  assign counters_MPORT_2_data = counters[counters_MPORT_2_addr]; // @[fetch.scala 149:21]
  assign counters_MPORT_4_en = io_branchres_fired & _GEN_271;
  assign counters_MPORT_4_addr = {io_branchres_pc[7:2],_counterIndex_train_T_15};
  assign counters_MPORT_4_data = counters[counters_MPORT_4_addr]; // @[fetch.scala 149:21]
  assign counters_MPORT_5_en = io_branchres_fired & _GEN_276;
  assign counters_MPORT_5_addr = {io_branchres_pc[7:2],_counterIndex_train_T_15};
  assign counters_MPORT_5_data = counters[counters_MPORT_5_addr]; // @[fetch.scala 149:21]
  assign counters_MPORT_7_en = io_branchres_fired & _GEN_279;
  assign counters_MPORT_7_addr = {io_branchres_pc[7:2],_counterIndex_train_T_15};
  assign counters_MPORT_7_data = counters[counters_MPORT_7_addr]; // @[fetch.scala 149:21]
  assign counters_prediction_MPORT_en = 1'h1;
  assign counters_prediction_MPORT_addr = {io_curr_pc[7:2],_counterIndex_pred_T_15};
  assign counters_prediction_MPORT_data = counters[counters_prediction_MPORT_addr]; // @[fetch.scala 149:21]
  assign counters_MPORT_3_data = counters_MPORT_4_data + 2'h1;
  assign counters_MPORT_3_addr = {io_branchres_pc[7:2],_counterIndex_train_T_15};
  assign counters_MPORT_3_mask = 1'h1;
  assign counters_MPORT_3_en = io_branchres_fired & _GEN_271;
  assign counters_MPORT_6_data = counters_MPORT_7_data - 2'h1;
  assign counters_MPORT_6_addr = {io_branchres_pc[7:2],_counterIndex_train_T_15};
  assign counters_MPORT_6_mask = 1'h1;
  assign counters_MPORT_6_en = io_branchres_fired & _GEN_279;
  assign tag_store_btb_hit_MPORT_en = 1'h1;
  assign tag_store_btb_hit_MPORT_addr = io_curr_pc[9:2];
  assign tag_store_btb_hit_MPORT_data = tag_store[tag_store_btb_hit_MPORT_addr]; // @[fetch.scala 151:22]
  assign tag_store_MPORT_data = io_branchres_pc[63:10];
  assign tag_store_MPORT_addr = io_branchres_pc[9:2];
  assign tag_store_MPORT_mask = 1'h1;
  assign tag_store_MPORT_en = io_branchres_fired;
  assign io_next_pc = btb_hit & prediction ? btb_io_next_pc_MPORT_data : _io_next_pc_T_2; // @[fetch.scala 182:20]
  assign correct_history_clock = clock;
  assign correct_history_reset = reset;
  assign correct_history_in = io_branchres_branchTaken; // @[fetch.scala 126:22]
  assign correct_history_en = io_branchres_fired; // @[fetch.scala 125:44]
  assign predicted_history_clock = clock;
  assign predicted_history_reset = reset;
  assign predicted_history_in = counters_prediction_MPORT_data[1]; // @[fetch.scala 177:47]
  assign predicted_history_en = ~mispredicted & btb_hit & requestSent; // @[fetch.scala 179:52]
  assign predicted_history_updateVals_0 = mispredicted ? _GEN_1606 : correct_history_output_0; // @[fetch.scala 185:22 129:37]
  assign predicted_history_updateVals_1 = mispredicted ? _GEN_1607 : correct_history_output_1; // @[fetch.scala 185:22 129:37]
  assign predicted_history_updateVals_2 = mispredicted ? _GEN_1608 : correct_history_output_2; // @[fetch.scala 185:22 129:37]
  assign predicted_history_updateVals_3 = mispredicted ? _GEN_1609 : correct_history_output_3; // @[fetch.scala 185:22 129:37]
  assign predicted_history_updateVals_4 = mispredicted ? _GEN_1610 : correct_history_output_4; // @[fetch.scala 185:22 129:37]
  assign predicted_history_update = mispredicted; // @[fetch.scala 185:22 186:30 198:30]
  always @(posedge clock) begin
    if (btb_MPORT_1_en & btb_MPORT_1_mask) begin
      btb[btb_MPORT_1_addr] <= btb_MPORT_1_data; // @[fetch.scala 148:16]
    end
    if (counters_MPORT_3_en & counters_MPORT_3_mask) begin
      counters[counters_MPORT_3_addr] <= counters_MPORT_3_data; // @[fetch.scala 149:21]
    end
    if (counters_MPORT_6_en & counters_MPORT_6_mask) begin
      counters[counters_MPORT_6_addr] <= counters_MPORT_6_data; // @[fetch.scala 149:21]
    end
    if (tag_store_MPORT_en & tag_store_MPORT_mask) begin
      tag_store[tag_store_MPORT_addr] <= tag_store_MPORT_data; // @[fetch.scala 151:22]
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_0 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_0 <= _GEN_0;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_1 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_1 <= _GEN_1;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_2 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_2 <= _GEN_2;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_3 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_3 <= _GEN_3;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_4 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_4 <= _GEN_4;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_5 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_5 <= _GEN_5;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_6 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_6 <= _GEN_6;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_7 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_7 <= _GEN_7;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_8 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_8 <= _GEN_8;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_9 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_9 <= _GEN_9;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_10 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_10 <= _GEN_10;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_11 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_11 <= _GEN_11;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_12 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_12 <= _GEN_12;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_13 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_13 <= _GEN_13;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_14 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_14 <= _GEN_14;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_15 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_15 <= _GEN_15;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_16 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_16 <= _GEN_16;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_17 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_17 <= _GEN_17;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_18 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_18 <= _GEN_18;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_19 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_19 <= _GEN_19;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_20 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_20 <= _GEN_20;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_21 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_21 <= _GEN_21;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_22 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_22 <= _GEN_22;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_23 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_23 <= _GEN_23;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_24 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_24 <= _GEN_24;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_25 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_25 <= _GEN_25;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_26 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_26 <= _GEN_26;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_27 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_27 <= _GEN_27;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_28 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_28 <= _GEN_28;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_29 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_29 <= _GEN_29;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_30 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_30 <= _GEN_30;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_31 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_31 <= _GEN_31;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_32 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_32 <= _GEN_32;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_33 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_33 <= _GEN_33;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_34 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_34 <= _GEN_34;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_35 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_35 <= _GEN_35;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_36 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_36 <= _GEN_36;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_37 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_37 <= _GEN_37;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_38 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_38 <= _GEN_38;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_39 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_39 <= _GEN_39;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_40 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_40 <= _GEN_40;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_41 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_41 <= _GEN_41;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_42 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_42 <= _GEN_42;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_43 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_43 <= _GEN_43;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_44 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_44 <= _GEN_44;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_45 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_45 <= _GEN_45;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_46 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_46 <= _GEN_46;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_47 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_47 <= _GEN_47;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_48 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_48 <= _GEN_48;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_49 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_49 <= _GEN_49;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_50 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_50 <= _GEN_50;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_51 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_51 <= _GEN_51;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_52 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_52 <= _GEN_52;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_53 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_53 <= _GEN_53;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_54 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_54 <= _GEN_54;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_55 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_55 <= _GEN_55;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_56 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_56 <= _GEN_56;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_57 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_57 <= _GEN_57;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_58 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_58 <= _GEN_58;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_59 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_59 <= _GEN_59;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_60 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_60 <= _GEN_60;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_61 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_61 <= _GEN_61;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_62 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_62 <= _GEN_62;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_63 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_63 <= _GEN_63;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_64 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_64 <= _GEN_64;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_65 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_65 <= _GEN_65;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_66 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_66 <= _GEN_66;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_67 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_67 <= _GEN_67;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_68 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_68 <= _GEN_68;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_69 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_69 <= _GEN_69;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_70 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_70 <= _GEN_70;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_71 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_71 <= _GEN_71;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_72 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_72 <= _GEN_72;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_73 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_73 <= _GEN_73;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_74 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_74 <= _GEN_74;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_75 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_75 <= _GEN_75;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_76 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_76 <= _GEN_76;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_77 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_77 <= _GEN_77;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_78 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_78 <= _GEN_78;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_79 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_79 <= _GEN_79;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_80 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_80 <= _GEN_80;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_81 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_81 <= _GEN_81;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_82 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_82 <= _GEN_82;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_83 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_83 <= _GEN_83;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_84 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_84 <= _GEN_84;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_85 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_85 <= _GEN_85;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_86 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_86 <= _GEN_86;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_87 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_87 <= _GEN_87;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_88 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_88 <= _GEN_88;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_89 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_89 <= _GEN_89;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_90 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_90 <= _GEN_90;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_91 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_91 <= _GEN_91;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_92 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_92 <= _GEN_92;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_93 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_93 <= _GEN_93;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_94 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_94 <= _GEN_94;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_95 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_95 <= _GEN_95;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_96 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_96 <= _GEN_96;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_97 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_97 <= _GEN_97;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_98 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_98 <= _GEN_98;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_99 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_99 <= _GEN_99;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_100 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_100 <= _GEN_100;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_101 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_101 <= _GEN_101;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_102 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_102 <= _GEN_102;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_103 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_103 <= _GEN_103;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_104 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_104 <= _GEN_104;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_105 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_105 <= _GEN_105;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_106 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_106 <= _GEN_106;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_107 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_107 <= _GEN_107;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_108 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_108 <= _GEN_108;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_109 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_109 <= _GEN_109;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_110 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_110 <= _GEN_110;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_111 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_111 <= _GEN_111;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_112 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_112 <= _GEN_112;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_113 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_113 <= _GEN_113;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_114 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_114 <= _GEN_114;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_115 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_115 <= _GEN_115;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_116 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_116 <= _GEN_116;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_117 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_117 <= _GEN_117;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_118 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_118 <= _GEN_118;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_119 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_119 <= _GEN_119;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_120 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_120 <= _GEN_120;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_121 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_121 <= _GEN_121;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_122 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_122 <= _GEN_122;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_123 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_123 <= _GEN_123;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_124 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_124 <= _GEN_124;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_125 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_125 <= _GEN_125;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_126 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_126 <= _GEN_126;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_127 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_127 <= _GEN_127;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_128 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_128 <= _GEN_128;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_129 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_129 <= _GEN_129;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_130 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_130 <= _GEN_130;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_131 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_131 <= _GEN_131;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_132 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_132 <= _GEN_132;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_133 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_133 <= _GEN_133;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_134 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_134 <= _GEN_134;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_135 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_135 <= _GEN_135;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_136 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_136 <= _GEN_136;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_137 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_137 <= _GEN_137;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_138 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_138 <= _GEN_138;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_139 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_139 <= _GEN_139;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_140 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_140 <= _GEN_140;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_141 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_141 <= _GEN_141;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_142 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_142 <= _GEN_142;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_143 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_143 <= _GEN_143;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_144 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_144 <= _GEN_144;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_145 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_145 <= _GEN_145;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_146 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_146 <= _GEN_146;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_147 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_147 <= _GEN_147;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_148 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_148 <= _GEN_148;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_149 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_149 <= _GEN_149;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_150 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_150 <= _GEN_150;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_151 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_151 <= _GEN_151;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_152 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_152 <= _GEN_152;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_153 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_153 <= _GEN_153;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_154 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_154 <= _GEN_154;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_155 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_155 <= _GEN_155;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_156 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_156 <= _GEN_156;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_157 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_157 <= _GEN_157;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_158 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_158 <= _GEN_158;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_159 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_159 <= _GEN_159;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_160 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_160 <= _GEN_160;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_161 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_161 <= _GEN_161;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_162 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_162 <= _GEN_162;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_163 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_163 <= _GEN_163;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_164 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_164 <= _GEN_164;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_165 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_165 <= _GEN_165;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_166 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_166 <= _GEN_166;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_167 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_167 <= _GEN_167;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_168 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_168 <= _GEN_168;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_169 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_169 <= _GEN_169;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_170 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_170 <= _GEN_170;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_171 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_171 <= _GEN_171;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_172 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_172 <= _GEN_172;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_173 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_173 <= _GEN_173;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_174 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_174 <= _GEN_174;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_175 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_175 <= _GEN_175;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_176 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_176 <= _GEN_176;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_177 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_177 <= _GEN_177;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_178 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_178 <= _GEN_178;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_179 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_179 <= _GEN_179;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_180 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_180 <= _GEN_180;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_181 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_181 <= _GEN_181;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_182 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_182 <= _GEN_182;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_183 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_183 <= _GEN_183;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_184 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_184 <= _GEN_184;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_185 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_185 <= _GEN_185;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_186 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_186 <= _GEN_186;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_187 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_187 <= _GEN_187;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_188 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_188 <= _GEN_188;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_189 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_189 <= _GEN_189;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_190 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_190 <= _GEN_190;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_191 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_191 <= _GEN_191;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_192 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_192 <= _GEN_192;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_193 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_193 <= _GEN_193;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_194 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_194 <= _GEN_194;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_195 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_195 <= _GEN_195;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_196 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_196 <= _GEN_196;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_197 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_197 <= _GEN_197;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_198 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_198 <= _GEN_198;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_199 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_199 <= _GEN_199;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_200 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_200 <= _GEN_200;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_201 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_201 <= _GEN_201;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_202 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_202 <= _GEN_202;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_203 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_203 <= _GEN_203;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_204 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_204 <= _GEN_204;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_205 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_205 <= _GEN_205;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_206 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_206 <= _GEN_206;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_207 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_207 <= _GEN_207;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_208 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_208 <= _GEN_208;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_209 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_209 <= _GEN_209;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_210 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_210 <= _GEN_210;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_211 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_211 <= _GEN_211;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_212 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_212 <= _GEN_212;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_213 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_213 <= _GEN_213;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_214 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_214 <= _GEN_214;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_215 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_215 <= _GEN_215;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_216 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_216 <= _GEN_216;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_217 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_217 <= _GEN_217;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_218 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_218 <= _GEN_218;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_219 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_219 <= _GEN_219;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_220 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_220 <= _GEN_220;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_221 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_221 <= _GEN_221;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_222 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_222 <= _GEN_222;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_223 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_223 <= _GEN_223;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_224 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_224 <= _GEN_224;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_225 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_225 <= _GEN_225;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_226 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_226 <= _GEN_226;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_227 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_227 <= _GEN_227;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_228 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_228 <= _GEN_228;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_229 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_229 <= _GEN_229;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_230 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_230 <= _GEN_230;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_231 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_231 <= _GEN_231;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_232 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_232 <= _GEN_232;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_233 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_233 <= _GEN_233;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_234 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_234 <= _GEN_234;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_235 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_235 <= _GEN_235;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_236 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_236 <= _GEN_236;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_237 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_237 <= _GEN_237;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_238 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_238 <= _GEN_238;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_239 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_239 <= _GEN_239;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_240 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_240 <= _GEN_240;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_241 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_241 <= _GEN_241;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_242 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_242 <= _GEN_242;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_243 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_243 <= _GEN_243;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_244 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_244 <= _GEN_244;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_245 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_245 <= _GEN_245;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_246 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_246 <= _GEN_246;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_247 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_247 <= _GEN_247;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_248 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_248 <= _GEN_248;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_249 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_249 <= _GEN_249;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_250 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_250 <= _GEN_250;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_251 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_251 <= _GEN_251;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_252 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_252 <= _GEN_252;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_253 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_253 <= _GEN_253;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_254 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_254 <= _GEN_254;
    end
    if (reset) begin // @[fetch.scala 150:27]
      valid_bits_255 <= 1'h0; // @[fetch.scala 150:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 154:27]
      valid_bits_255 <= _GEN_255;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    btb[initvar] = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    counters[initvar] = _RAND_1[1:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    tag_store[initvar] = _RAND_2[53:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  valid_bits_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  valid_bits_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  valid_bits_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  valid_bits_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  valid_bits_4 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  valid_bits_5 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  valid_bits_6 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  valid_bits_7 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  valid_bits_8 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  valid_bits_9 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  valid_bits_10 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  valid_bits_11 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  valid_bits_12 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  valid_bits_13 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  valid_bits_14 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  valid_bits_15 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  valid_bits_16 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  valid_bits_17 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  valid_bits_18 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  valid_bits_19 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  valid_bits_20 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  valid_bits_21 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  valid_bits_22 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid_bits_23 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  valid_bits_24 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  valid_bits_25 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  valid_bits_26 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  valid_bits_27 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  valid_bits_28 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  valid_bits_29 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  valid_bits_30 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  valid_bits_31 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  valid_bits_32 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  valid_bits_33 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  valid_bits_34 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  valid_bits_35 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  valid_bits_36 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  valid_bits_37 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  valid_bits_38 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  valid_bits_39 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  valid_bits_40 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  valid_bits_41 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  valid_bits_42 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  valid_bits_43 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  valid_bits_44 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  valid_bits_45 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  valid_bits_46 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  valid_bits_47 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  valid_bits_48 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  valid_bits_49 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  valid_bits_50 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  valid_bits_51 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  valid_bits_52 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  valid_bits_53 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  valid_bits_54 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  valid_bits_55 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  valid_bits_56 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  valid_bits_57 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  valid_bits_58 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  valid_bits_59 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  valid_bits_60 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  valid_bits_61 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  valid_bits_62 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  valid_bits_63 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  valid_bits_64 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  valid_bits_65 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  valid_bits_66 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  valid_bits_67 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  valid_bits_68 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  valid_bits_69 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  valid_bits_70 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  valid_bits_71 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  valid_bits_72 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  valid_bits_73 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  valid_bits_74 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  valid_bits_75 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  valid_bits_76 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  valid_bits_77 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_bits_78 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_bits_79 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_bits_80 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_bits_81 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_bits_82 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_bits_83 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_bits_84 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_bits_85 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_bits_86 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_bits_87 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_bits_88 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_bits_89 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_bits_90 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_bits_91 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_bits_92 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  valid_bits_93 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  valid_bits_94 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  valid_bits_95 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  valid_bits_96 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  valid_bits_97 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  valid_bits_98 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  valid_bits_99 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  valid_bits_100 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  valid_bits_101 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  valid_bits_102 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  valid_bits_103 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  valid_bits_104 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  valid_bits_105 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  valid_bits_106 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  valid_bits_107 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  valid_bits_108 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  valid_bits_109 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  valid_bits_110 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  valid_bits_111 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  valid_bits_112 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  valid_bits_113 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  valid_bits_114 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  valid_bits_115 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  valid_bits_116 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  valid_bits_117 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  valid_bits_118 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  valid_bits_119 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  valid_bits_120 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  valid_bits_121 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  valid_bits_122 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  valid_bits_123 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  valid_bits_124 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  valid_bits_125 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_bits_126 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_bits_127 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_bits_128 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_bits_129 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_bits_130 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_bits_131 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  valid_bits_132 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  valid_bits_133 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  valid_bits_134 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  valid_bits_135 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  valid_bits_136 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  valid_bits_137 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  valid_bits_138 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  valid_bits_139 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  valid_bits_140 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  valid_bits_141 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  valid_bits_142 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  valid_bits_143 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  valid_bits_144 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  valid_bits_145 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  valid_bits_146 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  valid_bits_147 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  valid_bits_148 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  valid_bits_149 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  valid_bits_150 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  valid_bits_151 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  valid_bits_152 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  valid_bits_153 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  valid_bits_154 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  valid_bits_155 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  valid_bits_156 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  valid_bits_157 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_bits_158 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_bits_159 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_bits_160 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  valid_bits_161 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  valid_bits_162 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  valid_bits_163 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  valid_bits_164 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  valid_bits_165 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  valid_bits_166 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  valid_bits_167 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  valid_bits_168 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  valid_bits_169 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  valid_bits_170 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  valid_bits_171 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  valid_bits_172 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  valid_bits_173 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  valid_bits_174 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  valid_bits_175 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  valid_bits_176 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  valid_bits_177 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  valid_bits_178 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  valid_bits_179 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  valid_bits_180 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  valid_bits_181 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  valid_bits_182 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  valid_bits_183 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  valid_bits_184 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  valid_bits_185 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  valid_bits_186 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  valid_bits_187 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  valid_bits_188 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  valid_bits_189 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  valid_bits_190 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  valid_bits_191 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  valid_bits_192 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  valid_bits_193 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  valid_bits_194 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  valid_bits_195 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  valid_bits_196 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  valid_bits_197 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  valid_bits_198 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  valid_bits_199 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  valid_bits_200 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  valid_bits_201 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  valid_bits_202 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  valid_bits_203 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  valid_bits_204 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  valid_bits_205 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  valid_bits_206 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  valid_bits_207 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  valid_bits_208 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  valid_bits_209 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  valid_bits_210 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  valid_bits_211 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  valid_bits_212 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  valid_bits_213 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  valid_bits_214 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  valid_bits_215 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  valid_bits_216 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  valid_bits_217 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  valid_bits_218 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  valid_bits_219 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  valid_bits_220 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  valid_bits_221 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  valid_bits_222 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  valid_bits_223 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  valid_bits_224 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  valid_bits_225 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  valid_bits_226 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  valid_bits_227 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  valid_bits_228 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  valid_bits_229 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  valid_bits_230 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  valid_bits_231 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  valid_bits_232 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  valid_bits_233 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  valid_bits_234 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  valid_bits_235 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  valid_bits_236 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  valid_bits_237 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  valid_bits_238 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  valid_bits_239 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  valid_bits_240 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  valid_bits_241 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  valid_bits_242 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  valid_bits_243 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  valid_bits_244 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  valid_bits_245 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  valid_bits_246 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  valid_bits_247 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  valid_bits_248 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  valid_bits_249 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  valid_bits_250 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  valid_bits_251 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  valid_bits_252 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  valid_bits_253 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  valid_bits_254 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  valid_bits_255 = _RAND_258[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module regFifo(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [127:0] io_enq_bits,
  input          io_deq_ready,
  output         io_deq_valid,
  output [127:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] memReg [0:3]; // @[Fifo.scala 21:19]
  wire  memReg_io_deq_bits_MPORT_en; // @[Fifo.scala 21:19]
  wire [1:0] memReg_io_deq_bits_MPORT_addr; // @[Fifo.scala 21:19]
  wire [127:0] memReg_io_deq_bits_MPORT_data; // @[Fifo.scala 21:19]
  wire [127:0] memReg_MPORT_data; // @[Fifo.scala 21:19]
  wire [1:0] memReg_MPORT_addr; // @[Fifo.scala 21:19]
  wire  memReg_MPORT_mask; // @[Fifo.scala 21:19]
  wire  memReg_MPORT_en; // @[Fifo.scala 21:19]
  wire [127:0] memReg_MPORT_1_data; // @[Fifo.scala 21:19]
  wire [1:0] memReg_MPORT_1_addr; // @[Fifo.scala 21:19]
  wire  memReg_MPORT_1_mask; // @[Fifo.scala 21:19]
  wire  memReg_MPORT_1_en; // @[Fifo.scala 21:19]
  reg [1:0] readPtr; // @[Fifo.scala 12:26]
  wire [1:0] _nextVal_T_2 = readPtr + 2'h1; // @[Fifo.scala 13:60]
  wire [1:0] nextRead = readPtr == 2'h3 ? 2'h0 : _nextVal_T_2; // @[Fifo.scala 13:22]
  wire  _T = io_deq_ready & io_deq_valid; // @[Fifo.scala 30:21]
  wire  _T_1 = io_deq_ready & io_deq_valid & io_enq_valid; // @[Fifo.scala 30:37]
  wire  _T_2 = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready; // @[Fifo.scala 30:53]
  wire  _T_3 = io_enq_valid & io_enq_ready; // @[Fifo.scala 34:27]
  wire  _GEN_12 = io_enq_valid & io_enq_ready ? 1'h0 : _T; // @[Fifo.scala 34:44]
  wire  incrRead = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready | _GEN_12; // @[Fifo.scala 30:70 33:14]
  reg [1:0] writePtr; // @[Fifo.scala 12:26]
  wire [1:0] _nextVal_T_5 = writePtr + 2'h1; // @[Fifo.scala 13:60]
  wire [1:0] nextWrite = writePtr == 2'h3 ? 2'h0 : _nextVal_T_5; // @[Fifo.scala 13:22]
  wire  incrWrite = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready | _T_3; // @[Fifo.scala 30:70 32:15]
  reg  emptyReg; // @[Fifo.scala 26:25]
  reg  fullReg; // @[Fifo.scala 27:24]
  wire  _GEN_3 = _T ? nextRead == writePtr : emptyReg; // @[Fifo.scala 39:44 41:14 26:25]
  wire  _GEN_10 = io_enq_valid & io_enq_ready ? 1'h0 : _GEN_3; // @[Fifo.scala 34:44 36:14]
  wire  _GEN_25 = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready ? emptyReg : _GEN_10; // @[Fifo.scala 26:25 30:70]
  assign memReg_io_deq_bits_MPORT_en = 1'h1;
  assign memReg_io_deq_bits_MPORT_addr = readPtr;
  assign memReg_io_deq_bits_MPORT_data = memReg[memReg_io_deq_bits_MPORT_addr]; // @[Fifo.scala 21:19]
  assign memReg_MPORT_data = io_enq_bits;
  assign memReg_MPORT_addr = writePtr;
  assign memReg_MPORT_mask = 1'h1;
  assign memReg_MPORT_en = _T_1 & io_enq_ready;
  assign memReg_MPORT_1_data = io_enq_bits;
  assign memReg_MPORT_1_addr = writePtr;
  assign memReg_MPORT_1_mask = 1'h1;
  assign memReg_MPORT_1_en = _T_2 ? 1'h0 : _T_3;
  assign io_enq_ready = ~fullReg | io_deq_valid & io_deq_ready; // @[Fifo.scala 46:28]
  assign io_deq_valid = ~emptyReg; // @[Fifo.scala 47:19]
  assign io_deq_bits = memReg_io_deq_bits_MPORT_data; // @[Fifo.scala 45:15]
  always @(posedge clock) begin
    if (memReg_MPORT_en & memReg_MPORT_mask) begin
      memReg[memReg_MPORT_addr] <= memReg_MPORT_data; // @[Fifo.scala 21:19]
    end
    if (memReg_MPORT_1_en & memReg_MPORT_1_mask) begin
      memReg[memReg_MPORT_1_addr] <= memReg_MPORT_1_data; // @[Fifo.scala 21:19]
    end
    if (reset) begin // @[Fifo.scala 12:26]
      readPtr <= 2'h0; // @[Fifo.scala 12:26]
    end else if (incrRead) begin // @[Fifo.scala 14:17]
      if (readPtr == 2'h3) begin // @[Fifo.scala 13:22]
        readPtr <= 2'h0;
      end else begin
        readPtr <= _nextVal_T_2;
      end
    end
    if (reset) begin // @[Fifo.scala 12:26]
      writePtr <= 2'h0; // @[Fifo.scala 12:26]
    end else if (incrWrite) begin // @[Fifo.scala 14:17]
      if (writePtr == 2'h3) begin // @[Fifo.scala 13:22]
        writePtr <= 2'h0;
      end else begin
        writePtr <= _nextVal_T_5;
      end
    end
    emptyReg <= reset | _GEN_25; // @[Fifo.scala 26:{25,25}]
    if (reset) begin // @[Fifo.scala 27:24]
      fullReg <= 1'h0; // @[Fifo.scala 27:24]
    end else if (!(io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready)) begin // @[Fifo.scala 30:70]
      if (io_enq_valid & io_enq_ready) begin // @[Fifo.scala 34:44]
        fullReg <= nextWrite == readPtr; // @[Fifo.scala 37:13]
      end else if (_T) begin // @[Fifo.scala 39:44]
        fullReg <= 1'h0; // @[Fifo.scala 40:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    memReg[initvar] = _RAND_0[127:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  readPtr = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  writePtr = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  emptyReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  fullReg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module fetch(
  input         clock,
  input         reset,
  input         cache_req_ready,
  output        cache_req_valid,
  output [63:0] cache_req_bits,
  output        cache_resp_ready,
  input         cache_resp_valid,
  input  [31:0] cache_resp_bits,
  output        toDecode_ready,
  input         toDecode_fired,
  output [63:0] toDecode_pc,
  output [31:0] toDecode_instruction,
  input         toDecode_expected_valid,
  input  [63:0] toDecode_expected_pc,
  input         toDecode_expected_coherency,
  input         branchRes_fired,
  input         branchRes_branchTaken,
  input  [63:0] branchRes_pc,
  input  [63:0] branchRes_pcAfterBrnach,
  output        carryOutFence_ready,
  input         carryOutFence_fired,
  output        updateAllCachelines_ready,
  input         updateAllCachelines_fired,
  output        cachelinesUpdatesResp_ready,
  input         cachelinesUpdatesResp_fired,
  output        fdbg_probe_redirect_bit,
  output        fdbg_probe_fifo_enq_ready,
  output        fdbg_probe_is_fence,
  output        fdbg_probe_handle_fence
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  predictor_clock; // @[fetch.scala 259:25]
  wire  predictor_reset; // @[fetch.scala 259:25]
  wire  predictor_io_branchres_fired; // @[fetch.scala 259:25]
  wire  predictor_io_branchres_branchTaken; // @[fetch.scala 259:25]
  wire [63:0] predictor_io_branchres_pc; // @[fetch.scala 259:25]
  wire [63:0] predictor_io_branchres_pcAfterBrnach; // @[fetch.scala 259:25]
  wire [63:0] predictor_io_curr_pc; // @[fetch.scala 259:25]
  wire [63:0] predictor_io_next_pc; // @[fetch.scala 259:25]
  wire  predictor_requestSent; // @[fetch.scala 259:25]
  wire  predictor_mispredicted; // @[fetch.scala 259:25]
  wire  PC_fifo_clock; // @[fetch.scala 262:23]
  wire  PC_fifo_reset; // @[fetch.scala 262:23]
  wire  PC_fifo_io_enq_ready; // @[fetch.scala 262:23]
  wire  PC_fifo_io_enq_valid; // @[fetch.scala 262:23]
  wire [127:0] PC_fifo_io_enq_bits; // @[fetch.scala 262:23]
  wire  PC_fifo_io_deq_ready; // @[fetch.scala 262:23]
  wire  PC_fifo_io_deq_valid; // @[fetch.scala 262:23]
  wire [127:0] PC_fifo_io_deq_bits; // @[fetch.scala 262:23]
  reg [63:0] PC; // @[fetch.scala 250:19]
  reg  redirect_bit; // @[fetch.scala 251:28]
  reg  handle_fenceI; // @[fetch.scala 252:29]
  reg  clear_cache_req; // @[fetch.scala 253:31]
  reg  cache_cleared; // @[fetch.scala 254:29]
  reg  fence_pending; // @[fetch.scala 255:29]
  wire  _PC_fifo_io_enq_valid_T = cache_req_valid & cache_req_ready; // @[fetch.scala 266:43]
  wire  is_fenceI = toDecode_instruction[6:2] == 5'h3 & toDecode_instruction[14:13] == 2'h0 & toDecode_fired; // @[fetch.scala 271:102]
  wire  _T_1 = ~handle_fenceI; // @[fetch.scala 275:23]
  wire  _T_2 = ~clear_cache_req; // @[fetch.scala 278:26]
  wire  _T_3 = ~cache_cleared; // @[fetch.scala 278:49]
  wire  _T_5 = ~fence_pending; // @[fetch.scala 278:72]
  wire  redirect = ~(toDecode_expected_pc == toDecode_pc) & toDecode_expected_valid; // @[fetch.scala 307:55]
  wire  _T_19 = ~redirect_bit; // @[fetch.scala 311:20]
  wire  _T_20 = ~redirect_bit & PC_fifo_io_deq_valid; // @[fetch.scala 311:27]
  wire  _T_21 = ~PC_fifo_io_deq_valid; // @[fetch.scala 313:36]
  wire [127:0] _PC_T_1 = PC_fifo_io_deq_bits + 128'h4; // @[fetch.scala 322:31]
  wire [63:0] _GEN_11 = _PC_fifo_io_enq_valid_T ? predictor_io_next_pc : PC; // @[fetch.scala 250:19 323:49 324:8]
  wire [127:0] _GEN_12 = is_fenceI ? _PC_T_1 : {{64'd0}, _GEN_11}; // @[fetch.scala 321:25 322:8]
  wire [127:0] _GEN_13 = redirect_bit ? {{64'd0}, toDecode_expected_pc} : _GEN_12; // @[fetch.scala 319:28 320:8]
  reg  misPredicted; // @[fetch.scala 353:29]
  wire  _GEN_15 = _T_20 & (redirect & ~toDecode_expected_coherency); // @[fetch.scala 354:51 355:18 357:18]
  wire [127:0] _GEN_17 = reset ? 128'h10000000 : _GEN_13; // @[fetch.scala 250:{19,19}]
  gshare_predictor predictor ( // @[fetch.scala 259:25]
    .clock(predictor_clock),
    .reset(predictor_reset),
    .io_branchres_fired(predictor_io_branchres_fired),
    .io_branchres_branchTaken(predictor_io_branchres_branchTaken),
    .io_branchres_pc(predictor_io_branchres_pc),
    .io_branchres_pcAfterBrnach(predictor_io_branchres_pcAfterBrnach),
    .io_curr_pc(predictor_io_curr_pc),
    .io_next_pc(predictor_io_next_pc),
    .requestSent(predictor_requestSent),
    .mispredicted(predictor_mispredicted)
  );
  regFifo PC_fifo ( // @[fetch.scala 262:23]
    .clock(PC_fifo_clock),
    .reset(PC_fifo_reset),
    .io_enq_ready(PC_fifo_io_enq_ready),
    .io_enq_valid(PC_fifo_io_enq_valid),
    .io_enq_bits(PC_fifo_io_enq_bits),
    .io_deq_ready(PC_fifo_io_deq_ready),
    .io_deq_valid(PC_fifo_io_deq_valid),
    .io_deq_bits(PC_fifo_io_deq_bits)
  );
  assign cache_req_valid = _T_19 & PC_fifo_io_enq_ready & ~is_fenceI & _T_1; // @[fetch.scala 329:79]
  assign cache_req_bits = PC; // @[fetch.scala 326:18]
  assign cache_resp_ready = handle_fenceI | (redirect_bit | toDecode_fired) & _T_1; // @[fetch.scala 330:20 361:{30,49}]
  assign toDecode_ready = redirect | redirect_bit | ~cache_resp_valid | _T_21 | handle_fenceI ? 1'h0 : 1'h1; // @[fetch.scala 342:109 343:20 345:20]
  assign toDecode_pc = PC_fifo_io_deq_bits[63:0]; // @[fetch.scala 268:15]
  assign toDecode_instruction = cache_resp_bits; // @[fetch.scala 348:24]
  assign carryOutFence_ready = fence_pending; // @[fetch.scala 295:23]
  assign updateAllCachelines_ready = clear_cache_req; // @[fetch.scala 331:29]
  assign cachelinesUpdatesResp_ready = cache_cleared; // @[fetch.scala 332:31]
  assign fdbg_probe_redirect_bit = redirect_bit; // @[fetch.scala 336:27]
  assign fdbg_probe_fifo_enq_ready = PC_fifo_io_enq_ready; // @[fetch.scala 337:29]
  assign fdbg_probe_is_fence = toDecode_instruction[6:2] == 5'h3 & toDecode_instruction[14:13] == 2'h0 & toDecode_fired; // @[fetch.scala 271:102]
  assign fdbg_probe_handle_fence = handle_fenceI; // @[fetch.scala 339:27]
  assign predictor_clock = clock;
  assign predictor_reset = reset;
  assign predictor_io_branchres_fired = branchRes_fired; // @[fetch.scala 260:26]
  assign predictor_io_branchres_branchTaken = branchRes_branchTaken; // @[fetch.scala 260:26]
  assign predictor_io_branchres_pc = branchRes_pc; // @[fetch.scala 260:26]
  assign predictor_io_branchres_pcAfterBrnach = branchRes_pcAfterBrnach; // @[fetch.scala 260:26]
  assign predictor_io_curr_pc = PC; // @[fetch.scala 261:24]
  assign predictor_requestSent = cache_req_valid & cache_req_ready; // @[fetch.scala 350:44]
  assign predictor_mispredicted = misPredicted; // @[fetch.scala 360:26]
  assign PC_fifo_clock = clock;
  assign PC_fifo_reset = handle_fenceI | reset; // @[fetch.scala 272:29 273:18]
  assign PC_fifo_io_enq_valid = cache_req_valid & cache_req_ready; // @[fetch.scala 266:43]
  assign PC_fifo_io_enq_bits = {{64'd0}, PC}; // @[fetch.scala 265:23]
  assign PC_fifo_io_deq_ready = cache_resp_valid & cache_resp_ready; // @[fetch.scala 267:44]
  always @(posedge clock) begin
    PC <= _GEN_17[63:0]; // @[fetch.scala 250:{19,19}]
    if (reset) begin // @[fetch.scala 251:28]
      redirect_bit <= 1'h0; // @[fetch.scala 251:28]
    end else if (~redirect_bit & PC_fifo_io_deq_valid) begin // @[fetch.scala 311:50]
      redirect_bit <= redirect; // @[fetch.scala 312:18]
    end else if (~PC_fifo_io_deq_valid) begin // @[fetch.scala 313:44]
      redirect_bit <= 1'h0; // @[fetch.scala 314:18]
    end
    if (reset) begin // @[fetch.scala 252:29]
      handle_fenceI <= 1'h0; // @[fetch.scala 252:29]
    end else if (~handle_fenceI) begin // @[fetch.scala 275:31]
      handle_fenceI <= is_fenceI; // @[fetch.scala 276:19]
    end else if (~clear_cache_req & ~cache_cleared & ~fence_pending) begin // @[fetch.scala 278:79]
      handle_fenceI <= 1'h0; // @[fetch.scala 279:21]
    end
    if (reset) begin // @[fetch.scala 253:31]
      clear_cache_req <= 1'h0; // @[fetch.scala 253:31]
    end else if (_T_2 & _T_1) begin // @[fetch.scala 283:54]
      clear_cache_req <= is_fenceI; // @[fetch.scala 284:21]
    end else if (updateAllCachelines_fired) begin // @[fetch.scala 285:40]
      clear_cache_req <= 1'h0; // @[fetch.scala 286:21]
    end
    if (reset) begin // @[fetch.scala 254:29]
      cache_cleared <= 1'h0; // @[fetch.scala 254:29]
    end else if (_T_3 & _T_1) begin // @[fetch.scala 289:54]
      cache_cleared <= is_fenceI; // @[fetch.scala 290:19]
    end else if (cachelinesUpdatesResp_fired) begin // @[fetch.scala 291:43]
      cache_cleared <= 1'h0; // @[fetch.scala 292:19]
    end
    if (reset) begin // @[fetch.scala 255:29]
      fence_pending <= 1'h0; // @[fetch.scala 255:29]
    end else if (_T_5 & _T_1) begin // @[fetch.scala 297:52]
      fence_pending <= is_fenceI; // @[fetch.scala 298:18]
    end else if (carryOutFence_fired) begin // @[fetch.scala 299:34]
      fence_pending <= 1'h0; // @[fetch.scala 300:18]
    end
    if (reset) begin // @[fetch.scala 353:29]
      misPredicted <= 1'h0; // @[fetch.scala 353:29]
    end else begin
      misPredicted <= _GEN_15;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  PC = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  redirect_bit = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  handle_fenceI = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  clear_cache_req = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  cache_cleared = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  fence_pending = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  misPredicted = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module core_Anon(
  input         clock,
  input         reset,
  output        fromFetch_ready,
  input         fromFetch_fired,
  input  [63:0] fromFetch_pc,
  input  [31:0] fromFetch_instruction,
  output        fromFetch_expected_valid,
  output [63:0] fromFetch_expected_pc,
  output        fromFetch_expected_coherency,
  output        toExec_ready,
  input         toExec_fired,
  output [31:0] toExec_instruction,
  output [63:0] toExec_pc,
  output [5:0]  toExec_PRFDest,
  output [5:0]  toExec_rs1Addr,
  output        toExec_rs1Ready,
  output [5:0]  toExec_rs2Addr,
  output        toExec_rs2Ready,
  output [4:0]  toExec_branchMask,
  input         writeBackResult_fired,
  input  [31:0] writeBackResult_instruction,
  input  [4:0]  writeBackResult_rdAddr,
  input  [5:0]  writeBackResult_PRFDest,
  input  [63:0] writeBackResult_data,
  input  [5:0]  writeAddrPRF_exec1Addr,
  input  [5:0]  writeAddrPRF_exec2Addr,
  input  [5:0]  writeAddrPRF_exec3Addr,
  input         writeAddrPRF_exec1Valid,
  input         writeAddrPRF_exec2Valid,
  input         writeAddrPRF_exec3Valid,
  output        jumpAddrWrite_ready,
  input         jumpAddrWrite_fired,
  output [5:0]  jumpAddrWrite_PRFDest,
  output [63:0] jumpAddrWrite_linkAddr,
  output        branchPCs_branchPCReady,
  output [63:0] branchPCs_branchPC,
  output        branchPCs_predictedPCReady,
  output [63:0] branchPCs_predictedPC,
  output [4:0]  branchPCs_branchMask,
  input         branchEvalIn_fired,
  input         branchEvalIn_passFail,
  input  [4:0]  branchEvalIn_branchMask,
  input  [63:0] branchEvalIn_targetPC,
  input  [63:0] interruptedPC,
  output        canTakeInterrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [63:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [63:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [63:0] _RAND_856;
  reg [63:0] _RAND_857;
  reg [63:0] _RAND_858;
  reg [63:0] _RAND_859;
  reg [63:0] _RAND_860;
  reg [63:0] _RAND_861;
  reg [63:0] _RAND_862;
  reg [63:0] _RAND_863;
  reg [63:0] _RAND_864;
  reg [63:0] _RAND_865;
  reg [63:0] _RAND_866;
  reg [63:0] _RAND_867;
  reg [63:0] _RAND_868;
  reg [63:0] _RAND_869;
  reg [63:0] _RAND_870;
  reg [63:0] _RAND_871;
  reg [63:0] _RAND_872;
  reg [63:0] _RAND_873;
  reg [63:0] _RAND_874;
  reg [63:0] _RAND_875;
  reg [63:0] _RAND_876;
  reg [63:0] _RAND_877;
  reg [63:0] _RAND_878;
  reg [63:0] _RAND_879;
  reg [63:0] _RAND_880;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] inputBuffer_pc; // @[decode.scala 111:28]
  reg [31:0] inputBuffer_instruction; // @[decode.scala 111:28]
  reg [31:0] outputBuffer_instruction; // @[decode.scala 120:29]
  reg [63:0] outputBuffer_pc; // @[decode.scala 120:29]
  reg [5:0] outputBuffer_PRFDest; // @[decode.scala 120:29]
  reg [5:0] outputBuffer_rs1Addr; // @[decode.scala 120:29]
  reg [5:0] outputBuffer_rs2Addr; // @[decode.scala 120:29]
  reg [63:0] outputBuffer_immediate; // @[decode.scala 120:29]
  reg  branchBuffer_branchPCReady; // @[decode.scala 142:29]
  reg  branchBuffer_predictedPCReady; // @[decode.scala 142:29]
  reg [63:0] branchBuffer_branchPC; // @[decode.scala 142:29]
  reg [63:0] branchBuffer_predictedPC; // @[decode.scala 142:29]
  reg  branchBuffer_branchMask_0; // @[decode.scala 142:29]
  reg  branchBuffer_branchMask_1; // @[decode.scala 142:29]
  reg  branchBuffer_branchMask_2; // @[decode.scala 142:29]
  reg  branchBuffer_branchMask_3; // @[decode.scala 142:29]
  reg  branchBuffer_branchMask_4; // @[decode.scala 142:29]
  reg [2:0] branchTracker; // @[decode.scala 178:30]
  reg [63:0] expectedPC; // @[decode.scala 188:27]
  reg  coherency; // @[decode.scala 189:26]
  reg  stateRegInputBuf; // @[decode.scala 193:34]
  reg  stateRegOutputBuf; // @[decode.scala 194:34]
  reg  stallReg; // @[decode.scala 196:25]
  reg [63:0] ecallPC; // @[decode.scala 197:20]
  reg  PRFValidList_0; // @[decode.scala 199:29]
  reg  PRFValidList_1; // @[decode.scala 199:29]
  reg  PRFValidList_2; // @[decode.scala 199:29]
  reg  PRFValidList_3; // @[decode.scala 199:29]
  reg  PRFValidList_4; // @[decode.scala 199:29]
  reg  PRFValidList_5; // @[decode.scala 199:29]
  reg  PRFValidList_6; // @[decode.scala 199:29]
  reg  PRFValidList_7; // @[decode.scala 199:29]
  reg  PRFValidList_8; // @[decode.scala 199:29]
  reg  PRFValidList_9; // @[decode.scala 199:29]
  reg  PRFValidList_10; // @[decode.scala 199:29]
  reg  PRFValidList_11; // @[decode.scala 199:29]
  reg  PRFValidList_12; // @[decode.scala 199:29]
  reg  PRFValidList_13; // @[decode.scala 199:29]
  reg  PRFValidList_14; // @[decode.scala 199:29]
  reg  PRFValidList_15; // @[decode.scala 199:29]
  reg  PRFValidList_16; // @[decode.scala 199:29]
  reg  PRFValidList_17; // @[decode.scala 199:29]
  reg  PRFValidList_18; // @[decode.scala 199:29]
  reg  PRFValidList_19; // @[decode.scala 199:29]
  reg  PRFValidList_20; // @[decode.scala 199:29]
  reg  PRFValidList_21; // @[decode.scala 199:29]
  reg  PRFValidList_22; // @[decode.scala 199:29]
  reg  PRFValidList_23; // @[decode.scala 199:29]
  reg  PRFValidList_24; // @[decode.scala 199:29]
  reg  PRFValidList_25; // @[decode.scala 199:29]
  reg  PRFValidList_26; // @[decode.scala 199:29]
  reg  PRFValidList_27; // @[decode.scala 199:29]
  reg  PRFValidList_28; // @[decode.scala 199:29]
  reg  PRFValidList_29; // @[decode.scala 199:29]
  reg  PRFValidList_30; // @[decode.scala 199:29]
  reg  PRFValidList_31; // @[decode.scala 199:29]
  reg  PRFValidList_32; // @[decode.scala 199:29]
  reg  PRFValidList_33; // @[decode.scala 199:29]
  reg  PRFValidList_34; // @[decode.scala 199:29]
  reg  PRFValidList_35; // @[decode.scala 199:29]
  reg  PRFValidList_36; // @[decode.scala 199:29]
  reg  PRFValidList_37; // @[decode.scala 199:29]
  reg  PRFValidList_38; // @[decode.scala 199:29]
  reg  PRFValidList_39; // @[decode.scala 199:29]
  reg  PRFValidList_40; // @[decode.scala 199:29]
  reg  PRFValidList_41; // @[decode.scala 199:29]
  reg  PRFValidList_42; // @[decode.scala 199:29]
  reg  PRFValidList_43; // @[decode.scala 199:29]
  reg  PRFValidList_44; // @[decode.scala 199:29]
  reg  PRFValidList_45; // @[decode.scala 199:29]
  reg  PRFValidList_46; // @[decode.scala 199:29]
  reg  PRFValidList_47; // @[decode.scala 199:29]
  reg  PRFValidList_48; // @[decode.scala 199:29]
  reg  PRFValidList_49; // @[decode.scala 199:29]
  reg  PRFValidList_50; // @[decode.scala 199:29]
  reg  PRFValidList_51; // @[decode.scala 199:29]
  reg  PRFValidList_52; // @[decode.scala 199:29]
  reg  PRFValidList_53; // @[decode.scala 199:29]
  reg  PRFValidList_54; // @[decode.scala 199:29]
  reg  PRFValidList_55; // @[decode.scala 199:29]
  reg  PRFValidList_56; // @[decode.scala 199:29]
  reg  PRFValidList_57; // @[decode.scala 199:29]
  reg  PRFValidList_58; // @[decode.scala 199:29]
  reg  PRFValidList_59; // @[decode.scala 199:29]
  reg  PRFValidList_60; // @[decode.scala 199:29]
  reg  PRFValidList_61; // @[decode.scala 199:29]
  reg  PRFValidList_62; // @[decode.scala 199:29]
  reg  PRFValidList_63; // @[decode.scala 199:29]
  wire  _T_434 = ~branchEvalIn_passFail; // @[decode.scala 794:34]
  wire  _T_435 = branchEvalIn_fired & ~branchEvalIn_passFail; // @[decode.scala 794:31]
  wire  _GEN_13361 = branchEvalIn_fired & ~branchEvalIn_passFail ? 1'h0 : 1'h1; // @[decode.scala 794:58 797:26 801:23]
  wire  _GEN_13363 = stallReg ? 1'h0 : _GEN_13361; // @[decode.scala 812:22 813:23]
  wire [4:0] rs1 = inputBuffer_instruction[19:15]; // @[decode.scala 297:16]
  reg [5:0] frontEndRegMap_31; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_30; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_29; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_28; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_27; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_26; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_25; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_24; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_23; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_22; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_21; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_20; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_19; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_18; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_17; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_16; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_15; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_14; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_13; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_12; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_11; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_10; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_9; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_8; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_7; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_6; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_5; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_4; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_3; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_2; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_1; // @[decode.scala 308:36]
  reg [5:0] frontEndRegMap_0; // @[decode.scala 308:36]
  wire [5:0] _GEN_209 = 5'h1 == rs1 ? frontEndRegMap_1 : frontEndRegMap_0; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_210 = 5'h2 == rs1 ? frontEndRegMap_2 : _GEN_209; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_211 = 5'h3 == rs1 ? frontEndRegMap_3 : _GEN_210; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_212 = 5'h4 == rs1 ? frontEndRegMap_4 : _GEN_211; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_213 = 5'h5 == rs1 ? frontEndRegMap_5 : _GEN_212; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_214 = 5'h6 == rs1 ? frontEndRegMap_6 : _GEN_213; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_215 = 5'h7 == rs1 ? frontEndRegMap_7 : _GEN_214; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_216 = 5'h8 == rs1 ? frontEndRegMap_8 : _GEN_215; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_217 = 5'h9 == rs1 ? frontEndRegMap_9 : _GEN_216; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_218 = 5'ha == rs1 ? frontEndRegMap_10 : _GEN_217; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_219 = 5'hb == rs1 ? frontEndRegMap_11 : _GEN_218; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_220 = 5'hc == rs1 ? frontEndRegMap_12 : _GEN_219; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_221 = 5'hd == rs1 ? frontEndRegMap_13 : _GEN_220; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_222 = 5'he == rs1 ? frontEndRegMap_14 : _GEN_221; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_223 = 5'hf == rs1 ? frontEndRegMap_15 : _GEN_222; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_224 = 5'h10 == rs1 ? frontEndRegMap_16 : _GEN_223; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_225 = 5'h11 == rs1 ? frontEndRegMap_17 : _GEN_224; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_226 = 5'h12 == rs1 ? frontEndRegMap_18 : _GEN_225; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_227 = 5'h13 == rs1 ? frontEndRegMap_19 : _GEN_226; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_228 = 5'h14 == rs1 ? frontEndRegMap_20 : _GEN_227; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_229 = 5'h15 == rs1 ? frontEndRegMap_21 : _GEN_228; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_230 = 5'h16 == rs1 ? frontEndRegMap_22 : _GEN_229; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_231 = 5'h17 == rs1 ? frontEndRegMap_23 : _GEN_230; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_232 = 5'h18 == rs1 ? frontEndRegMap_24 : _GEN_231; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_233 = 5'h19 == rs1 ? frontEndRegMap_25 : _GEN_232; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_234 = 5'h1a == rs1 ? frontEndRegMap_26 : _GEN_233; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_235 = 5'h1b == rs1 ? frontEndRegMap_27 : _GEN_234; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_236 = 5'h1c == rs1 ? frontEndRegMap_28 : _GEN_235; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_237 = 5'h1d == rs1 ? frontEndRegMap_29 : _GEN_236; // @[decode.scala 332:{12,12}]
  wire [5:0] _GEN_238 = 5'h1e == rs1 ? frontEndRegMap_30 : _GEN_237; // @[decode.scala 332:{12,12}]
  wire [5:0] rs1Addr = 5'h1f == rs1 ? frontEndRegMap_31 : _GEN_238; // @[decode.scala 332:{12,12}]
  reg  PRFFreeList_0; // @[decode.scala 310:36]
  reg  PRFFreeList_1; // @[decode.scala 310:36]
  reg  PRFFreeList_2; // @[decode.scala 310:36]
  reg  PRFFreeList_3; // @[decode.scala 310:36]
  reg  PRFFreeList_4; // @[decode.scala 310:36]
  reg  PRFFreeList_5; // @[decode.scala 310:36]
  reg  PRFFreeList_6; // @[decode.scala 310:36]
  reg  PRFFreeList_7; // @[decode.scala 310:36]
  reg  PRFFreeList_8; // @[decode.scala 310:36]
  reg  PRFFreeList_9; // @[decode.scala 310:36]
  reg  PRFFreeList_10; // @[decode.scala 310:36]
  reg  PRFFreeList_11; // @[decode.scala 310:36]
  reg  PRFFreeList_12; // @[decode.scala 310:36]
  reg  PRFFreeList_13; // @[decode.scala 310:36]
  reg  PRFFreeList_14; // @[decode.scala 310:36]
  reg  PRFFreeList_15; // @[decode.scala 310:36]
  reg  PRFFreeList_16; // @[decode.scala 310:36]
  reg  PRFFreeList_17; // @[decode.scala 310:36]
  reg  PRFFreeList_18; // @[decode.scala 310:36]
  reg  PRFFreeList_19; // @[decode.scala 310:36]
  reg  PRFFreeList_20; // @[decode.scala 310:36]
  reg  PRFFreeList_21; // @[decode.scala 310:36]
  reg  PRFFreeList_22; // @[decode.scala 310:36]
  reg  PRFFreeList_23; // @[decode.scala 310:36]
  reg  PRFFreeList_24; // @[decode.scala 310:36]
  reg  PRFFreeList_25; // @[decode.scala 310:36]
  reg  PRFFreeList_26; // @[decode.scala 310:36]
  reg  PRFFreeList_27; // @[decode.scala 310:36]
  reg  PRFFreeList_28; // @[decode.scala 310:36]
  reg  PRFFreeList_29; // @[decode.scala 310:36]
  reg  PRFFreeList_30; // @[decode.scala 310:36]
  reg  PRFFreeList_31; // @[decode.scala 310:36]
  reg  PRFFreeList_32; // @[decode.scala 310:36]
  reg  PRFFreeList_33; // @[decode.scala 310:36]
  reg  PRFFreeList_34; // @[decode.scala 310:36]
  reg  PRFFreeList_35; // @[decode.scala 310:36]
  reg  PRFFreeList_36; // @[decode.scala 310:36]
  reg  PRFFreeList_37; // @[decode.scala 310:36]
  reg  PRFFreeList_38; // @[decode.scala 310:36]
  reg  PRFFreeList_39; // @[decode.scala 310:36]
  reg  PRFFreeList_40; // @[decode.scala 310:36]
  reg  PRFFreeList_41; // @[decode.scala 310:36]
  reg  PRFFreeList_42; // @[decode.scala 310:36]
  reg  PRFFreeList_43; // @[decode.scala 310:36]
  reg  PRFFreeList_44; // @[decode.scala 310:36]
  reg  PRFFreeList_45; // @[decode.scala 310:36]
  reg  PRFFreeList_46; // @[decode.scala 310:36]
  reg  PRFFreeList_47; // @[decode.scala 310:36]
  reg  PRFFreeList_48; // @[decode.scala 310:36]
  reg  PRFFreeList_49; // @[decode.scala 310:36]
  reg  PRFFreeList_50; // @[decode.scala 310:36]
  reg  PRFFreeList_51; // @[decode.scala 310:36]
  reg  PRFFreeList_52; // @[decode.scala 310:36]
  reg  PRFFreeList_53; // @[decode.scala 310:36]
  reg  PRFFreeList_54; // @[decode.scala 310:36]
  reg  PRFFreeList_55; // @[decode.scala 310:36]
  reg  PRFFreeList_56; // @[decode.scala 310:36]
  reg  PRFFreeList_57; // @[decode.scala 310:36]
  reg  PRFFreeList_58; // @[decode.scala 310:36]
  reg  PRFFreeList_59; // @[decode.scala 310:36]
  reg  PRFFreeList_60; // @[decode.scala 310:36]
  reg  PRFFreeList_61; // @[decode.scala 310:36]
  reg  PRFFreeList_62; // @[decode.scala 310:36]
  wire [5:0] _freeRegAddr_T = PRFFreeList_62 ? 6'h3e : 6'h3f; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_1 = PRFFreeList_61 ? 6'h3d : _freeRegAddr_T; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_2 = PRFFreeList_60 ? 6'h3c : _freeRegAddr_T_1; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_3 = PRFFreeList_59 ? 6'h3b : _freeRegAddr_T_2; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_4 = PRFFreeList_58 ? 6'h3a : _freeRegAddr_T_3; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_5 = PRFFreeList_57 ? 6'h39 : _freeRegAddr_T_4; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_6 = PRFFreeList_56 ? 6'h38 : _freeRegAddr_T_5; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_7 = PRFFreeList_55 ? 6'h37 : _freeRegAddr_T_6; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_8 = PRFFreeList_54 ? 6'h36 : _freeRegAddr_T_7; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_9 = PRFFreeList_53 ? 6'h35 : _freeRegAddr_T_8; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_10 = PRFFreeList_52 ? 6'h34 : _freeRegAddr_T_9; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_11 = PRFFreeList_51 ? 6'h33 : _freeRegAddr_T_10; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_12 = PRFFreeList_50 ? 6'h32 : _freeRegAddr_T_11; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_13 = PRFFreeList_49 ? 6'h31 : _freeRegAddr_T_12; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_14 = PRFFreeList_48 ? 6'h30 : _freeRegAddr_T_13; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_15 = PRFFreeList_47 ? 6'h2f : _freeRegAddr_T_14; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_16 = PRFFreeList_46 ? 6'h2e : _freeRegAddr_T_15; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_17 = PRFFreeList_45 ? 6'h2d : _freeRegAddr_T_16; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_18 = PRFFreeList_44 ? 6'h2c : _freeRegAddr_T_17; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_19 = PRFFreeList_43 ? 6'h2b : _freeRegAddr_T_18; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_20 = PRFFreeList_42 ? 6'h2a : _freeRegAddr_T_19; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_21 = PRFFreeList_41 ? 6'h29 : _freeRegAddr_T_20; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_22 = PRFFreeList_40 ? 6'h28 : _freeRegAddr_T_21; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_23 = PRFFreeList_39 ? 6'h27 : _freeRegAddr_T_22; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_24 = PRFFreeList_38 ? 6'h26 : _freeRegAddr_T_23; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_25 = PRFFreeList_37 ? 6'h25 : _freeRegAddr_T_24; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_26 = PRFFreeList_36 ? 6'h24 : _freeRegAddr_T_25; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_27 = PRFFreeList_35 ? 6'h23 : _freeRegAddr_T_26; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_28 = PRFFreeList_34 ? 6'h22 : _freeRegAddr_T_27; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_29 = PRFFreeList_33 ? 6'h21 : _freeRegAddr_T_28; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_30 = PRFFreeList_32 ? 6'h20 : _freeRegAddr_T_29; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_31 = PRFFreeList_31 ? 6'h1f : _freeRegAddr_T_30; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_32 = PRFFreeList_30 ? 6'h1e : _freeRegAddr_T_31; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_33 = PRFFreeList_29 ? 6'h1d : _freeRegAddr_T_32; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_34 = PRFFreeList_28 ? 6'h1c : _freeRegAddr_T_33; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_35 = PRFFreeList_27 ? 6'h1b : _freeRegAddr_T_34; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_36 = PRFFreeList_26 ? 6'h1a : _freeRegAddr_T_35; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_37 = PRFFreeList_25 ? 6'h19 : _freeRegAddr_T_36; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_38 = PRFFreeList_24 ? 6'h18 : _freeRegAddr_T_37; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_39 = PRFFreeList_23 ? 6'h17 : _freeRegAddr_T_38; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_40 = PRFFreeList_22 ? 6'h16 : _freeRegAddr_T_39; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_41 = PRFFreeList_21 ? 6'h15 : _freeRegAddr_T_40; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_42 = PRFFreeList_20 ? 6'h14 : _freeRegAddr_T_41; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_43 = PRFFreeList_19 ? 6'h13 : _freeRegAddr_T_42; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_44 = PRFFreeList_18 ? 6'h12 : _freeRegAddr_T_43; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_45 = PRFFreeList_17 ? 6'h11 : _freeRegAddr_T_44; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_46 = PRFFreeList_16 ? 6'h10 : _freeRegAddr_T_45; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_47 = PRFFreeList_15 ? 6'hf : _freeRegAddr_T_46; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_48 = PRFFreeList_14 ? 6'he : _freeRegAddr_T_47; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_49 = PRFFreeList_13 ? 6'hd : _freeRegAddr_T_48; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_50 = PRFFreeList_12 ? 6'hc : _freeRegAddr_T_49; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_51 = PRFFreeList_11 ? 6'hb : _freeRegAddr_T_50; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_52 = PRFFreeList_10 ? 6'ha : _freeRegAddr_T_51; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_53 = PRFFreeList_9 ? 6'h9 : _freeRegAddr_T_52; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_54 = PRFFreeList_8 ? 6'h8 : _freeRegAddr_T_53; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_55 = PRFFreeList_7 ? 6'h7 : _freeRegAddr_T_54; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_56 = PRFFreeList_6 ? 6'h6 : _freeRegAddr_T_55; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_57 = PRFFreeList_5 ? 6'h5 : _freeRegAddr_T_56; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_58 = PRFFreeList_4 ? 6'h4 : _freeRegAddr_T_57; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_59 = PRFFreeList_3 ? 6'h3 : _freeRegAddr_T_58; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_60 = PRFFreeList_2 ? 6'h2 : _freeRegAddr_T_59; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_61 = PRFFreeList_1 ? 6'h1 : _freeRegAddr_T_60; // @[Mux.scala 47:70]
  wire [5:0] freeRegAddr = PRFFreeList_0 ? 6'h0 : _freeRegAddr_T_61; // @[Mux.scala 47:70]
  wire  _T_21 = rs1Addr == freeRegAddr; // @[decode.scala 342:16]
  wire [4:0] rs2 = inputBuffer_instruction[24:20]; // @[decode.scala 298:16]
  wire [5:0] _GEN_241 = 5'h1 == rs2 ? frontEndRegMap_1 : frontEndRegMap_0; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_242 = 5'h2 == rs2 ? frontEndRegMap_2 : _GEN_241; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_243 = 5'h3 == rs2 ? frontEndRegMap_3 : _GEN_242; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_244 = 5'h4 == rs2 ? frontEndRegMap_4 : _GEN_243; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_245 = 5'h5 == rs2 ? frontEndRegMap_5 : _GEN_244; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_246 = 5'h6 == rs2 ? frontEndRegMap_6 : _GEN_245; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_247 = 5'h7 == rs2 ? frontEndRegMap_7 : _GEN_246; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_248 = 5'h8 == rs2 ? frontEndRegMap_8 : _GEN_247; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_249 = 5'h9 == rs2 ? frontEndRegMap_9 : _GEN_248; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_250 = 5'ha == rs2 ? frontEndRegMap_10 : _GEN_249; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_251 = 5'hb == rs2 ? frontEndRegMap_11 : _GEN_250; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_252 = 5'hc == rs2 ? frontEndRegMap_12 : _GEN_251; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_253 = 5'hd == rs2 ? frontEndRegMap_13 : _GEN_252; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_254 = 5'he == rs2 ? frontEndRegMap_14 : _GEN_253; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_255 = 5'hf == rs2 ? frontEndRegMap_15 : _GEN_254; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_256 = 5'h10 == rs2 ? frontEndRegMap_16 : _GEN_255; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_257 = 5'h11 == rs2 ? frontEndRegMap_17 : _GEN_256; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_258 = 5'h12 == rs2 ? frontEndRegMap_18 : _GEN_257; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_259 = 5'h13 == rs2 ? frontEndRegMap_19 : _GEN_258; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_260 = 5'h14 == rs2 ? frontEndRegMap_20 : _GEN_259; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_261 = 5'h15 == rs2 ? frontEndRegMap_21 : _GEN_260; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_262 = 5'h16 == rs2 ? frontEndRegMap_22 : _GEN_261; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_263 = 5'h17 == rs2 ? frontEndRegMap_23 : _GEN_262; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_264 = 5'h18 == rs2 ? frontEndRegMap_24 : _GEN_263; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_265 = 5'h19 == rs2 ? frontEndRegMap_25 : _GEN_264; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_266 = 5'h1a == rs2 ? frontEndRegMap_26 : _GEN_265; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_267 = 5'h1b == rs2 ? frontEndRegMap_27 : _GEN_266; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_268 = 5'h1c == rs2 ? frontEndRegMap_28 : _GEN_267; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_269 = 5'h1d == rs2 ? frontEndRegMap_29 : _GEN_268; // @[decode.scala 333:{12,12}]
  wire [5:0] _GEN_270 = 5'h1e == rs2 ? frontEndRegMap_30 : _GEN_269; // @[decode.scala 333:{12,12}]
  wire [5:0] rs2Addr = 5'h1f == rs2 ? frontEndRegMap_31 : _GEN_270; // @[decode.scala 333:{12,12}]
  wire  _T_22 = rs2Addr == freeRegAddr; // @[decode.scala 342:43]
  wire [6:0] opcode = inputBuffer_instruction[6:0]; // @[decode.scala 296:16]
  wire  _T_5 = 7'h6f == opcode; // @[decode.scala 338:69]
  wire  _T_6 = 7'h67 == opcode; // @[decode.scala 338:69]
  wire  _T_7 = 7'h63 == opcode; // @[decode.scala 338:69]
  wire  _T_20 = freeRegAddr == 6'h3f | (7'h6f == opcode | 7'h67 == opcode | 7'h63 == opcode) & (
    branchBuffer_branchMask_0 & branchBuffer_branchMask_1 & branchBuffer_branchMask_2 & branchBuffer_branchMask_3 &
    branchBuffer_branchMask_4); // @[decode.scala 338:29]
  wire  stall = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr | _T_20; // @[decode.scala 342:60 343:11]
  wire  _T_441 = opcode == 7'h63; // @[decode.scala 823:56]
  wire  _T_442 = opcode == 7'h6f; // @[decode.scala 823:78]
  wire  _T_444 = opcode == 7'h67; // @[decode.scala 823:99]
  wire  _T_445 = opcode == 7'h63 | opcode == 7'h6f | opcode == 7'h67; // @[decode.scala 823:89]
  wire  _T_448 = ~stall & ~(branchEvalIn_fired & (opcode == 7'h63 | opcode == 7'h6f | opcode == 7'h67)); // @[decode.scala 823:21]
  wire  _GEN_13392 = _T_435 ? 1'h0 : toExec_fired; // @[decode.scala 861:58 864:27]
  wire  readyOutputBuf = ~stateRegOutputBuf ? _GEN_13361 : stateRegOutputBuf & _GEN_13392; // @[decode.scala 846:29]
  wire  _GEN_13368 = ~stall & ~(branchEvalIn_fired & (opcode == 7'h63 | opcode == 7'h6f | opcode == 7'h67)) &
    readyOutputBuf; // @[decode.scala 823:114]
  wire  _GEN_13372 = _T_435 ? 1'h0 : _GEN_13368; // @[decode.scala 817:58 820:26]
  wire  _GEN_13374 = stallReg ? 1'h0 : _GEN_13372; // @[decode.scala 837:22 838:23]
  wire  readyInputBuf = ~stateRegInputBuf ? _GEN_13363 : stateRegInputBuf & _GEN_13374; // @[decode.scala 792:28]
  wire  _GEN_0 = fromFetch_instruction[6:0] == 7'h73 | stallReg; // @[decode.scala 205:97 206:16 196:25]
  wire  _GEN_4 = fromFetch_fired & readyInputBuf ? _GEN_0 : stallReg; // @[decode.scala 196:25 202:42]
  wire  _GEN_13371 = _T_435 ? 1'h0 : _T_448; // @[decode.scala 817:58 819:26]
  wire  validInputBuf = ~stateRegInputBuf ? 1'h0 : stateRegInputBuf & _GEN_13371; // @[decode.scala 792:28]
  wire  _T_3 = validInputBuf & readyOutputBuf; // @[decode.scala 212:22]
  wire [2:0] _GEN_188 = 7'hf == opcode ? 3'h6 : 3'h0; // @[utils.scala 10:20 48:17]
  wire [2:0] _GEN_189 = 7'h73 == opcode ? 3'h1 : _GEN_188; // @[utils.scala 10:20 45:17]
  wire [2:0] _GEN_190 = 7'h3b == opcode ? 3'h0 : _GEN_189; // @[utils.scala 10:20 42:17]
  wire [2:0] _GEN_191 = 7'h33 == opcode ? 3'h0 : _GEN_190; // @[utils.scala 10:20 39:17]
  wire [2:0] _GEN_192 = 7'h1b == opcode ? 3'h1 : _GEN_191; // @[utils.scala 10:20 36:17]
  wire [2:0] _GEN_193 = 7'h13 == opcode ? 3'h1 : _GEN_192; // @[utils.scala 10:20 33:17]
  wire [2:0] _GEN_194 = 7'h23 == opcode ? 3'h2 : _GEN_193; // @[utils.scala 10:20 30:17]
  wire [2:0] _GEN_195 = 7'h3 == opcode ? 3'h1 : _GEN_194; // @[utils.scala 10:20 27:17]
  wire [2:0] _GEN_196 = _T_7 ? 3'h3 : _GEN_195; // @[utils.scala 10:20 24:17]
  wire [2:0] _GEN_197 = _T_6 ? 3'h1 : _GEN_196; // @[utils.scala 10:20 21:17]
  wire [2:0] _GEN_198 = _T_5 ? 3'h5 : _GEN_197; // @[utils.scala 10:20 18:17]
  wire [2:0] _GEN_199 = 7'h17 == opcode ? 3'h4 : _GEN_198; // @[utils.scala 10:20 15:17]
  wire [2:0] insType_insType = 7'h37 == opcode ? 3'h4 : _GEN_199; // @[utils.scala 10:20 12:17]
  wire [52:0] _immediate_immediate_T_2 = inputBuffer_instruction[31] ? 53'h1fffffffffffff : 53'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _immediate_immediate_T_4 = {_immediate_immediate_T_2,inputBuffer_instruction[30:20]}; // @[Cat.scala 33:92]
  wire [63:0] _immediate_immediate_T_10 = {_immediate_immediate_T_2,inputBuffer_instruction[30:25],
    inputBuffer_instruction[11:7]}; // @[Cat.scala 33:92]
  wire [64:0] _immediate_immediate_T_17 = {_immediate_immediate_T_2,inputBuffer_instruction[7],inputBuffer_instruction[
    30:25],inputBuffer_instruction[11:8],1'h0}; // @[Cat.scala 33:92]
  wire [31:0] _immediate_immediate_T_20 = inputBuffer_instruction[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _immediate_immediate_T_22 = {_immediate_immediate_T_20,inputBuffer_instruction[31:12],12'h0}; // @[Cat.scala 33:92]
  wire [43:0] _immediate_immediate_T_25 = inputBuffer_instruction[31] ? 44'hfffffffffff : 44'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _immediate_immediate_T_30 = {_immediate_immediate_T_25,inputBuffer_instruction[19:12],
    inputBuffer_instruction[20],inputBuffer_instruction[30:25],inputBuffer_instruction[24:21],1'h0}; // @[Cat.scala 33:92]
  wire [63:0] _GEN_203 = 3'h5 == insType_insType ? _immediate_immediate_T_30 : 64'h0; // @[utils.scala 59:29 73:19]
  wire [63:0] _GEN_204 = 3'h4 == insType_insType ? _immediate_immediate_T_22 : _GEN_203; // @[utils.scala 59:29 70:19]
  wire [64:0] _GEN_205 = 3'h3 == insType_insType ? _immediate_immediate_T_17 : {{1'd0}, _GEN_204}; // @[utils.scala 59:29 67:19]
  wire [64:0] _GEN_206 = 3'h2 == insType_insType ? {{1'd0}, _immediate_immediate_T_10} : _GEN_205; // @[utils.scala 59:29 64:19]
  wire [64:0] _GEN_207 = 3'h1 == insType_insType ? {{1'd0}, _immediate_immediate_T_4} : _GEN_206; // @[utils.scala 59:29 61:19]
  wire [63:0] immediate_immediate = _GEN_207[63:0];
  reg [4:0] branchPCMask; // @[decode.scala 225:29]
  reg  branchReg; // @[decode.scala 226:29]
  reg [63:0] csrReadDataReg; // @[decode.scala 240:31]
  reg [11:0] csrAddrReg; // @[decode.scala 242:27]
  reg [63:0] csrImmReg; // @[decode.scala 243:26]
  wire  _GEN_13 = 6'h1 == outputBuffer_rs1Addr ? PRFValidList_1 : PRFValidList_0; // @[decode.scala 254:{22,22}]
  wire  _GEN_14 = 6'h2 == outputBuffer_rs1Addr ? PRFValidList_2 : _GEN_13; // @[decode.scala 254:{22,22}]
  wire  _GEN_15 = 6'h3 == outputBuffer_rs1Addr ? PRFValidList_3 : _GEN_14; // @[decode.scala 254:{22,22}]
  wire  _GEN_16 = 6'h4 == outputBuffer_rs1Addr ? PRFValidList_4 : _GEN_15; // @[decode.scala 254:{22,22}]
  wire  _GEN_17 = 6'h5 == outputBuffer_rs1Addr ? PRFValidList_5 : _GEN_16; // @[decode.scala 254:{22,22}]
  wire  _GEN_18 = 6'h6 == outputBuffer_rs1Addr ? PRFValidList_6 : _GEN_17; // @[decode.scala 254:{22,22}]
  wire  _GEN_19 = 6'h7 == outputBuffer_rs1Addr ? PRFValidList_7 : _GEN_18; // @[decode.scala 254:{22,22}]
  wire  _GEN_20 = 6'h8 == outputBuffer_rs1Addr ? PRFValidList_8 : _GEN_19; // @[decode.scala 254:{22,22}]
  wire  _GEN_21 = 6'h9 == outputBuffer_rs1Addr ? PRFValidList_9 : _GEN_20; // @[decode.scala 254:{22,22}]
  wire  _GEN_22 = 6'ha == outputBuffer_rs1Addr ? PRFValidList_10 : _GEN_21; // @[decode.scala 254:{22,22}]
  wire  _GEN_23 = 6'hb == outputBuffer_rs1Addr ? PRFValidList_11 : _GEN_22; // @[decode.scala 254:{22,22}]
  wire  _GEN_24 = 6'hc == outputBuffer_rs1Addr ? PRFValidList_12 : _GEN_23; // @[decode.scala 254:{22,22}]
  wire  _GEN_25 = 6'hd == outputBuffer_rs1Addr ? PRFValidList_13 : _GEN_24; // @[decode.scala 254:{22,22}]
  wire  _GEN_26 = 6'he == outputBuffer_rs1Addr ? PRFValidList_14 : _GEN_25; // @[decode.scala 254:{22,22}]
  wire  _GEN_27 = 6'hf == outputBuffer_rs1Addr ? PRFValidList_15 : _GEN_26; // @[decode.scala 254:{22,22}]
  wire  _GEN_28 = 6'h10 == outputBuffer_rs1Addr ? PRFValidList_16 : _GEN_27; // @[decode.scala 254:{22,22}]
  wire  _GEN_29 = 6'h11 == outputBuffer_rs1Addr ? PRFValidList_17 : _GEN_28; // @[decode.scala 254:{22,22}]
  wire  _GEN_30 = 6'h12 == outputBuffer_rs1Addr ? PRFValidList_18 : _GEN_29; // @[decode.scala 254:{22,22}]
  wire  _GEN_31 = 6'h13 == outputBuffer_rs1Addr ? PRFValidList_19 : _GEN_30; // @[decode.scala 254:{22,22}]
  wire  _GEN_32 = 6'h14 == outputBuffer_rs1Addr ? PRFValidList_20 : _GEN_31; // @[decode.scala 254:{22,22}]
  wire  _GEN_33 = 6'h15 == outputBuffer_rs1Addr ? PRFValidList_21 : _GEN_32; // @[decode.scala 254:{22,22}]
  wire  _GEN_34 = 6'h16 == outputBuffer_rs1Addr ? PRFValidList_22 : _GEN_33; // @[decode.scala 254:{22,22}]
  wire  _GEN_35 = 6'h17 == outputBuffer_rs1Addr ? PRFValidList_23 : _GEN_34; // @[decode.scala 254:{22,22}]
  wire  _GEN_36 = 6'h18 == outputBuffer_rs1Addr ? PRFValidList_24 : _GEN_35; // @[decode.scala 254:{22,22}]
  wire  _GEN_37 = 6'h19 == outputBuffer_rs1Addr ? PRFValidList_25 : _GEN_36; // @[decode.scala 254:{22,22}]
  wire  _GEN_38 = 6'h1a == outputBuffer_rs1Addr ? PRFValidList_26 : _GEN_37; // @[decode.scala 254:{22,22}]
  wire  _GEN_39 = 6'h1b == outputBuffer_rs1Addr ? PRFValidList_27 : _GEN_38; // @[decode.scala 254:{22,22}]
  wire  _GEN_40 = 6'h1c == outputBuffer_rs1Addr ? PRFValidList_28 : _GEN_39; // @[decode.scala 254:{22,22}]
  wire  _GEN_41 = 6'h1d == outputBuffer_rs1Addr ? PRFValidList_29 : _GEN_40; // @[decode.scala 254:{22,22}]
  wire  _GEN_42 = 6'h1e == outputBuffer_rs1Addr ? PRFValidList_30 : _GEN_41; // @[decode.scala 254:{22,22}]
  wire  _GEN_43 = 6'h1f == outputBuffer_rs1Addr ? PRFValidList_31 : _GEN_42; // @[decode.scala 254:{22,22}]
  wire  _GEN_44 = 6'h20 == outputBuffer_rs1Addr ? PRFValidList_32 : _GEN_43; // @[decode.scala 254:{22,22}]
  wire  _GEN_45 = 6'h21 == outputBuffer_rs1Addr ? PRFValidList_33 : _GEN_44; // @[decode.scala 254:{22,22}]
  wire  _GEN_46 = 6'h22 == outputBuffer_rs1Addr ? PRFValidList_34 : _GEN_45; // @[decode.scala 254:{22,22}]
  wire  _GEN_47 = 6'h23 == outputBuffer_rs1Addr ? PRFValidList_35 : _GEN_46; // @[decode.scala 254:{22,22}]
  wire  _GEN_48 = 6'h24 == outputBuffer_rs1Addr ? PRFValidList_36 : _GEN_47; // @[decode.scala 254:{22,22}]
  wire  _GEN_49 = 6'h25 == outputBuffer_rs1Addr ? PRFValidList_37 : _GEN_48; // @[decode.scala 254:{22,22}]
  wire  _GEN_50 = 6'h26 == outputBuffer_rs1Addr ? PRFValidList_38 : _GEN_49; // @[decode.scala 254:{22,22}]
  wire  _GEN_51 = 6'h27 == outputBuffer_rs1Addr ? PRFValidList_39 : _GEN_50; // @[decode.scala 254:{22,22}]
  wire  _GEN_52 = 6'h28 == outputBuffer_rs1Addr ? PRFValidList_40 : _GEN_51; // @[decode.scala 254:{22,22}]
  wire  _GEN_53 = 6'h29 == outputBuffer_rs1Addr ? PRFValidList_41 : _GEN_52; // @[decode.scala 254:{22,22}]
  wire  _GEN_54 = 6'h2a == outputBuffer_rs1Addr ? PRFValidList_42 : _GEN_53; // @[decode.scala 254:{22,22}]
  wire  _GEN_55 = 6'h2b == outputBuffer_rs1Addr ? PRFValidList_43 : _GEN_54; // @[decode.scala 254:{22,22}]
  wire  _GEN_56 = 6'h2c == outputBuffer_rs1Addr ? PRFValidList_44 : _GEN_55; // @[decode.scala 254:{22,22}]
  wire  _GEN_57 = 6'h2d == outputBuffer_rs1Addr ? PRFValidList_45 : _GEN_56; // @[decode.scala 254:{22,22}]
  wire  _GEN_58 = 6'h2e == outputBuffer_rs1Addr ? PRFValidList_46 : _GEN_57; // @[decode.scala 254:{22,22}]
  wire  _GEN_59 = 6'h2f == outputBuffer_rs1Addr ? PRFValidList_47 : _GEN_58; // @[decode.scala 254:{22,22}]
  wire  _GEN_60 = 6'h30 == outputBuffer_rs1Addr ? PRFValidList_48 : _GEN_59; // @[decode.scala 254:{22,22}]
  wire  _GEN_61 = 6'h31 == outputBuffer_rs1Addr ? PRFValidList_49 : _GEN_60; // @[decode.scala 254:{22,22}]
  wire  _GEN_62 = 6'h32 == outputBuffer_rs1Addr ? PRFValidList_50 : _GEN_61; // @[decode.scala 254:{22,22}]
  wire  _GEN_63 = 6'h33 == outputBuffer_rs1Addr ? PRFValidList_51 : _GEN_62; // @[decode.scala 254:{22,22}]
  wire  _GEN_64 = 6'h34 == outputBuffer_rs1Addr ? PRFValidList_52 : _GEN_63; // @[decode.scala 254:{22,22}]
  wire  _GEN_65 = 6'h35 == outputBuffer_rs1Addr ? PRFValidList_53 : _GEN_64; // @[decode.scala 254:{22,22}]
  wire  _GEN_66 = 6'h36 == outputBuffer_rs1Addr ? PRFValidList_54 : _GEN_65; // @[decode.scala 254:{22,22}]
  wire  _GEN_67 = 6'h37 == outputBuffer_rs1Addr ? PRFValidList_55 : _GEN_66; // @[decode.scala 254:{22,22}]
  wire  _GEN_68 = 6'h38 == outputBuffer_rs1Addr ? PRFValidList_56 : _GEN_67; // @[decode.scala 254:{22,22}]
  wire  _GEN_69 = 6'h39 == outputBuffer_rs1Addr ? PRFValidList_57 : _GEN_68; // @[decode.scala 254:{22,22}]
  wire  _GEN_70 = 6'h3a == outputBuffer_rs1Addr ? PRFValidList_58 : _GEN_69; // @[decode.scala 254:{22,22}]
  wire  _GEN_71 = 6'h3b == outputBuffer_rs1Addr ? PRFValidList_59 : _GEN_70; // @[decode.scala 254:{22,22}]
  wire  _GEN_72 = 6'h3c == outputBuffer_rs1Addr ? PRFValidList_60 : _GEN_71; // @[decode.scala 254:{22,22}]
  wire  _GEN_73 = 6'h3d == outputBuffer_rs1Addr ? PRFValidList_61 : _GEN_72; // @[decode.scala 254:{22,22}]
  wire  _GEN_74 = 6'h3e == outputBuffer_rs1Addr ? PRFValidList_62 : _GEN_73; // @[decode.scala 254:{22,22}]
  wire [2:0] _GEN_77 = 7'hf == outputBuffer_instruction[6:0] ? 3'h6 : 3'h0; // @[utils.scala 10:20 48:17]
  wire [2:0] _GEN_78 = 7'h73 == outputBuffer_instruction[6:0] ? 3'h1 : _GEN_77; // @[utils.scala 10:20 45:17]
  wire [2:0] _GEN_79 = 7'h3b == outputBuffer_instruction[6:0] ? 3'h0 : _GEN_78; // @[utils.scala 10:20 42:17]
  wire [2:0] _GEN_80 = 7'h33 == outputBuffer_instruction[6:0] ? 3'h0 : _GEN_79; // @[utils.scala 10:20 39:17]
  wire [2:0] _GEN_81 = 7'h1b == outputBuffer_instruction[6:0] ? 3'h1 : _GEN_80; // @[utils.scala 10:20 36:17]
  wire [2:0] _GEN_82 = 7'h13 == outputBuffer_instruction[6:0] ? 3'h1 : _GEN_81; // @[utils.scala 10:20 33:17]
  wire [2:0] _GEN_83 = 7'h23 == outputBuffer_instruction[6:0] ? 3'h2 : _GEN_82; // @[utils.scala 10:20 30:17]
  wire [2:0] _GEN_84 = 7'h3 == outputBuffer_instruction[6:0] ? 3'h1 : _GEN_83; // @[utils.scala 10:20 27:17]
  wire [2:0] _GEN_85 = 7'h63 == outputBuffer_instruction[6:0] ? 3'h3 : _GEN_84; // @[utils.scala 10:20 24:17]
  wire [2:0] _GEN_86 = 7'h67 == outputBuffer_instruction[6:0] ? 3'h1 : _GEN_85; // @[utils.scala 10:20 21:17]
  wire [2:0] _GEN_87 = 7'h6f == outputBuffer_instruction[6:0] ? 3'h5 : _GEN_86; // @[utils.scala 10:20 18:17]
  wire [2:0] _GEN_88 = 7'h17 == outputBuffer_instruction[6:0] ? 3'h4 : _GEN_87; // @[utils.scala 10:20 15:17]
  wire [2:0] toExec_rs2Ready_insType = 7'h37 == outputBuffer_instruction[6:0] ? 3'h4 : _GEN_88; // @[utils.scala 10:20 12:17]
  wire  _GEN_119 = 6'h1 == outputBuffer_rs2Addr ? PRFValidList_1 : PRFValidList_0; // @[decode.scala 256:{60,60}]
  wire  _GEN_120 = 6'h2 == outputBuffer_rs2Addr ? PRFValidList_2 : _GEN_119; // @[decode.scala 256:{60,60}]
  wire  _GEN_121 = 6'h3 == outputBuffer_rs2Addr ? PRFValidList_3 : _GEN_120; // @[decode.scala 256:{60,60}]
  wire  _GEN_122 = 6'h4 == outputBuffer_rs2Addr ? PRFValidList_4 : _GEN_121; // @[decode.scala 256:{60,60}]
  wire  _GEN_123 = 6'h5 == outputBuffer_rs2Addr ? PRFValidList_5 : _GEN_122; // @[decode.scala 256:{60,60}]
  wire  _GEN_124 = 6'h6 == outputBuffer_rs2Addr ? PRFValidList_6 : _GEN_123; // @[decode.scala 256:{60,60}]
  wire  _GEN_125 = 6'h7 == outputBuffer_rs2Addr ? PRFValidList_7 : _GEN_124; // @[decode.scala 256:{60,60}]
  wire  _GEN_126 = 6'h8 == outputBuffer_rs2Addr ? PRFValidList_8 : _GEN_125; // @[decode.scala 256:{60,60}]
  wire  _GEN_127 = 6'h9 == outputBuffer_rs2Addr ? PRFValidList_9 : _GEN_126; // @[decode.scala 256:{60,60}]
  wire  _GEN_128 = 6'ha == outputBuffer_rs2Addr ? PRFValidList_10 : _GEN_127; // @[decode.scala 256:{60,60}]
  wire  _GEN_129 = 6'hb == outputBuffer_rs2Addr ? PRFValidList_11 : _GEN_128; // @[decode.scala 256:{60,60}]
  wire  _GEN_130 = 6'hc == outputBuffer_rs2Addr ? PRFValidList_12 : _GEN_129; // @[decode.scala 256:{60,60}]
  wire  _GEN_131 = 6'hd == outputBuffer_rs2Addr ? PRFValidList_13 : _GEN_130; // @[decode.scala 256:{60,60}]
  wire  _GEN_132 = 6'he == outputBuffer_rs2Addr ? PRFValidList_14 : _GEN_131; // @[decode.scala 256:{60,60}]
  wire  _GEN_133 = 6'hf == outputBuffer_rs2Addr ? PRFValidList_15 : _GEN_132; // @[decode.scala 256:{60,60}]
  wire  _GEN_134 = 6'h10 == outputBuffer_rs2Addr ? PRFValidList_16 : _GEN_133; // @[decode.scala 256:{60,60}]
  wire  _GEN_135 = 6'h11 == outputBuffer_rs2Addr ? PRFValidList_17 : _GEN_134; // @[decode.scala 256:{60,60}]
  wire  _GEN_136 = 6'h12 == outputBuffer_rs2Addr ? PRFValidList_18 : _GEN_135; // @[decode.scala 256:{60,60}]
  wire  _GEN_137 = 6'h13 == outputBuffer_rs2Addr ? PRFValidList_19 : _GEN_136; // @[decode.scala 256:{60,60}]
  wire  _GEN_138 = 6'h14 == outputBuffer_rs2Addr ? PRFValidList_20 : _GEN_137; // @[decode.scala 256:{60,60}]
  wire  _GEN_139 = 6'h15 == outputBuffer_rs2Addr ? PRFValidList_21 : _GEN_138; // @[decode.scala 256:{60,60}]
  wire  _GEN_140 = 6'h16 == outputBuffer_rs2Addr ? PRFValidList_22 : _GEN_139; // @[decode.scala 256:{60,60}]
  wire  _GEN_141 = 6'h17 == outputBuffer_rs2Addr ? PRFValidList_23 : _GEN_140; // @[decode.scala 256:{60,60}]
  wire  _GEN_142 = 6'h18 == outputBuffer_rs2Addr ? PRFValidList_24 : _GEN_141; // @[decode.scala 256:{60,60}]
  wire  _GEN_143 = 6'h19 == outputBuffer_rs2Addr ? PRFValidList_25 : _GEN_142; // @[decode.scala 256:{60,60}]
  wire  _GEN_144 = 6'h1a == outputBuffer_rs2Addr ? PRFValidList_26 : _GEN_143; // @[decode.scala 256:{60,60}]
  wire  _GEN_145 = 6'h1b == outputBuffer_rs2Addr ? PRFValidList_27 : _GEN_144; // @[decode.scala 256:{60,60}]
  wire  _GEN_146 = 6'h1c == outputBuffer_rs2Addr ? PRFValidList_28 : _GEN_145; // @[decode.scala 256:{60,60}]
  wire  _GEN_147 = 6'h1d == outputBuffer_rs2Addr ? PRFValidList_29 : _GEN_146; // @[decode.scala 256:{60,60}]
  wire  _GEN_148 = 6'h1e == outputBuffer_rs2Addr ? PRFValidList_30 : _GEN_147; // @[decode.scala 256:{60,60}]
  wire  _GEN_149 = 6'h1f == outputBuffer_rs2Addr ? PRFValidList_31 : _GEN_148; // @[decode.scala 256:{60,60}]
  wire  _GEN_150 = 6'h20 == outputBuffer_rs2Addr ? PRFValidList_32 : _GEN_149; // @[decode.scala 256:{60,60}]
  wire  _GEN_151 = 6'h21 == outputBuffer_rs2Addr ? PRFValidList_33 : _GEN_150; // @[decode.scala 256:{60,60}]
  wire  _GEN_152 = 6'h22 == outputBuffer_rs2Addr ? PRFValidList_34 : _GEN_151; // @[decode.scala 256:{60,60}]
  wire  _GEN_153 = 6'h23 == outputBuffer_rs2Addr ? PRFValidList_35 : _GEN_152; // @[decode.scala 256:{60,60}]
  wire  _GEN_154 = 6'h24 == outputBuffer_rs2Addr ? PRFValidList_36 : _GEN_153; // @[decode.scala 256:{60,60}]
  wire  _GEN_155 = 6'h25 == outputBuffer_rs2Addr ? PRFValidList_37 : _GEN_154; // @[decode.scala 256:{60,60}]
  wire  _GEN_156 = 6'h26 == outputBuffer_rs2Addr ? PRFValidList_38 : _GEN_155; // @[decode.scala 256:{60,60}]
  wire  _GEN_157 = 6'h27 == outputBuffer_rs2Addr ? PRFValidList_39 : _GEN_156; // @[decode.scala 256:{60,60}]
  wire  _GEN_158 = 6'h28 == outputBuffer_rs2Addr ? PRFValidList_40 : _GEN_157; // @[decode.scala 256:{60,60}]
  wire  _GEN_159 = 6'h29 == outputBuffer_rs2Addr ? PRFValidList_41 : _GEN_158; // @[decode.scala 256:{60,60}]
  wire  _GEN_160 = 6'h2a == outputBuffer_rs2Addr ? PRFValidList_42 : _GEN_159; // @[decode.scala 256:{60,60}]
  wire  _GEN_161 = 6'h2b == outputBuffer_rs2Addr ? PRFValidList_43 : _GEN_160; // @[decode.scala 256:{60,60}]
  wire  _GEN_162 = 6'h2c == outputBuffer_rs2Addr ? PRFValidList_44 : _GEN_161; // @[decode.scala 256:{60,60}]
  wire  _GEN_163 = 6'h2d == outputBuffer_rs2Addr ? PRFValidList_45 : _GEN_162; // @[decode.scala 256:{60,60}]
  wire  _GEN_164 = 6'h2e == outputBuffer_rs2Addr ? PRFValidList_46 : _GEN_163; // @[decode.scala 256:{60,60}]
  wire  _GEN_165 = 6'h2f == outputBuffer_rs2Addr ? PRFValidList_47 : _GEN_164; // @[decode.scala 256:{60,60}]
  wire  _GEN_166 = 6'h30 == outputBuffer_rs2Addr ? PRFValidList_48 : _GEN_165; // @[decode.scala 256:{60,60}]
  wire  _GEN_167 = 6'h31 == outputBuffer_rs2Addr ? PRFValidList_49 : _GEN_166; // @[decode.scala 256:{60,60}]
  wire  _GEN_168 = 6'h32 == outputBuffer_rs2Addr ? PRFValidList_50 : _GEN_167; // @[decode.scala 256:{60,60}]
  wire  _GEN_169 = 6'h33 == outputBuffer_rs2Addr ? PRFValidList_51 : _GEN_168; // @[decode.scala 256:{60,60}]
  wire  _GEN_170 = 6'h34 == outputBuffer_rs2Addr ? PRFValidList_52 : _GEN_169; // @[decode.scala 256:{60,60}]
  wire  _GEN_171 = 6'h35 == outputBuffer_rs2Addr ? PRFValidList_53 : _GEN_170; // @[decode.scala 256:{60,60}]
  wire  _GEN_172 = 6'h36 == outputBuffer_rs2Addr ? PRFValidList_54 : _GEN_171; // @[decode.scala 256:{60,60}]
  wire  _GEN_173 = 6'h37 == outputBuffer_rs2Addr ? PRFValidList_55 : _GEN_172; // @[decode.scala 256:{60,60}]
  wire  _GEN_174 = 6'h38 == outputBuffer_rs2Addr ? PRFValidList_56 : _GEN_173; // @[decode.scala 256:{60,60}]
  wire  _GEN_175 = 6'h39 == outputBuffer_rs2Addr ? PRFValidList_57 : _GEN_174; // @[decode.scala 256:{60,60}]
  wire  _GEN_176 = 6'h3a == outputBuffer_rs2Addr ? PRFValidList_58 : _GEN_175; // @[decode.scala 256:{60,60}]
  wire  _GEN_177 = 6'h3b == outputBuffer_rs2Addr ? PRFValidList_59 : _GEN_176; // @[decode.scala 256:{60,60}]
  wire  _GEN_178 = 6'h3c == outputBuffer_rs2Addr ? PRFValidList_60 : _GEN_177; // @[decode.scala 256:{60,60}]
  wire  _GEN_179 = 6'h3d == outputBuffer_rs2Addr ? PRFValidList_61 : _GEN_178; // @[decode.scala 256:{60,60}]
  wire  _GEN_180 = 6'h3e == outputBuffer_rs2Addr ? PRFValidList_62 : _GEN_179; // @[decode.scala 256:{60,60}]
  wire  _GEN_181 = 6'h3f == outputBuffer_rs2Addr ? PRFValidList_63 : _GEN_180; // @[decode.scala 256:{60,60}]
  wire [1:0] toExec_branchMask_lo = {branchBuffer_branchMask_1,branchBuffer_branchMask_0}; // @[decode.scala 258:49]
  wire [2:0] toExec_branchMask_hi = {branchBuffer_branchMask_4,branchBuffer_branchMask_3,branchBuffer_branchMask_2}; // @[decode.scala 258:49]
  wire [4:0] _toExec_branchMask_T = {branchBuffer_branchMask_4,branchBuffer_branchMask_3,branchBuffer_branchMask_2,
    branchBuffer_branchMask_1,branchBuffer_branchMask_0}; // @[decode.scala 258:49]
  wire  _fromFetch_expected_valid_T = expectedPC != 64'h0; // @[decode.scala 261:42]
  wire  unconditionalJumps = outputBuffer_instruction[6:0] == 7'h6f | outputBuffer_instruction[6:0] == 7'h67 |
    outputBuffer_instruction[6:0] == 7'h37 | outputBuffer_instruction[6:0] == 7'h17; // @[decode.scala 305:154]
  wire  csrIns = outputBuffer_instruction[6:0] == 7'h73 & outputBuffer_instruction[14:12] != 3'h0; // @[decode.scala 306:56]
  wire  validOutputBuf = ~stateRegOutputBuf ? 1'h0 : stateRegOutputBuf & _GEN_13361; // @[decode.scala 846:29]
  wire [31:0] _jumpAddrWrite_linkAddr_T_2 = outputBuffer_instruction[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _jumpAddrWrite_linkAddr_T_4 = {_jumpAddrWrite_linkAddr_T_2,outputBuffer_instruction[31:12],12'h0}; // @[Cat.scala 33:92]
  wire [63:0] _jumpAddrWrite_linkAddr_T_6 = outputBuffer_pc + _jumpAddrWrite_linkAddr_T_4; // @[decode.scala 269:24]
  wire [63:0] _jumpAddrWrite_linkAddr_T_13 = outputBuffer_pc + 64'h4; // @[decode.scala 272:23]
  wire [63:0] _GEN_183 = 2'h1 == outputBuffer_instruction[6:5] ? _jumpAddrWrite_linkAddr_T_4 :
    _jumpAddrWrite_linkAddr_T_6; // @[decode.scala 268:{28,28}]
  wire [63:0] _GEN_184 = 2'h2 == outputBuffer_instruction[6:5] ? 64'h0 : _GEN_183; // @[decode.scala 268:{28,28}]
  wire [63:0] _GEN_185 = 2'h3 == outputBuffer_instruction[6:5] ? _jumpAddrWrite_linkAddr_T_13 : _GEN_184; // @[decode.scala 268:{28,28}]
  wire [2:0] fun3 = inputBuffer_instruction[14:12]; // @[decode.scala 300:16]
  reg [5:0] architecturalRegMap_0; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_1; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_2; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_3; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_4; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_5; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_6; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_7; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_8; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_9; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_10; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_11; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_12; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_13; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_14; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_15; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_16; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_17; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_18; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_19; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_20; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_21; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_22; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_23; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_24; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_25; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_26; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_27; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_28; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_29; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_30; // @[decode.scala 309:36]
  reg [5:0] architecturalRegMap_31; // @[decode.scala 309:36]
  reg [5:0] reservedRegMap1_0; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_1; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_2; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_3; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_4; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_5; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_6; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_7; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_8; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_9; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_10; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_11; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_12; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_13; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_14; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_15; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_16; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_17; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_18; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_19; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_20; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_21; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_22; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_23; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_24; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_25; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_26; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_27; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_28; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_29; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_30; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap1_31; // @[decode.scala 317:28]
  reg [5:0] reservedRegMap2_0; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_1; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_2; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_3; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_4; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_5; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_6; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_7; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_8; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_9; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_10; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_11; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_12; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_13; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_14; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_15; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_16; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_17; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_18; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_19; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_20; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_21; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_22; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_23; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_24; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_25; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_26; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_27; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_28; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_29; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_30; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap2_31; // @[decode.scala 318:28]
  reg [5:0] reservedRegMap3_0; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_1; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_2; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_3; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_4; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_5; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_6; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_7; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_8; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_9; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_10; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_11; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_12; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_13; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_14; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_15; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_16; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_17; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_18; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_19; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_20; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_21; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_22; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_23; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_24; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_25; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_26; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_27; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_28; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_29; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_30; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap3_31; // @[decode.scala 319:28]
  reg [5:0] reservedRegMap4_0; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_1; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_2; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_3; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_4; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_5; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_6; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_7; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_8; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_9; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_10; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_11; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_12; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_13; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_14; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_15; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_16; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_17; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_18; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_19; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_20; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_21; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_22; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_23; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_24; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_25; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_26; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_27; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_28; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_29; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_30; // @[decode.scala 320:28]
  reg [5:0] reservedRegMap4_31; // @[decode.scala 320:28]
  reg  reservedFreeList1_0; // @[decode.scala 322:30]
  reg  reservedFreeList1_1; // @[decode.scala 322:30]
  reg  reservedFreeList1_2; // @[decode.scala 322:30]
  reg  reservedFreeList1_3; // @[decode.scala 322:30]
  reg  reservedFreeList1_4; // @[decode.scala 322:30]
  reg  reservedFreeList1_5; // @[decode.scala 322:30]
  reg  reservedFreeList1_6; // @[decode.scala 322:30]
  reg  reservedFreeList1_7; // @[decode.scala 322:30]
  reg  reservedFreeList1_8; // @[decode.scala 322:30]
  reg  reservedFreeList1_9; // @[decode.scala 322:30]
  reg  reservedFreeList1_10; // @[decode.scala 322:30]
  reg  reservedFreeList1_11; // @[decode.scala 322:30]
  reg  reservedFreeList1_12; // @[decode.scala 322:30]
  reg  reservedFreeList1_13; // @[decode.scala 322:30]
  reg  reservedFreeList1_14; // @[decode.scala 322:30]
  reg  reservedFreeList1_15; // @[decode.scala 322:30]
  reg  reservedFreeList1_16; // @[decode.scala 322:30]
  reg  reservedFreeList1_17; // @[decode.scala 322:30]
  reg  reservedFreeList1_18; // @[decode.scala 322:30]
  reg  reservedFreeList1_19; // @[decode.scala 322:30]
  reg  reservedFreeList1_20; // @[decode.scala 322:30]
  reg  reservedFreeList1_21; // @[decode.scala 322:30]
  reg  reservedFreeList1_22; // @[decode.scala 322:30]
  reg  reservedFreeList1_23; // @[decode.scala 322:30]
  reg  reservedFreeList1_24; // @[decode.scala 322:30]
  reg  reservedFreeList1_25; // @[decode.scala 322:30]
  reg  reservedFreeList1_26; // @[decode.scala 322:30]
  reg  reservedFreeList1_27; // @[decode.scala 322:30]
  reg  reservedFreeList1_28; // @[decode.scala 322:30]
  reg  reservedFreeList1_29; // @[decode.scala 322:30]
  reg  reservedFreeList1_30; // @[decode.scala 322:30]
  reg  reservedFreeList1_31; // @[decode.scala 322:30]
  reg  reservedFreeList1_32; // @[decode.scala 322:30]
  reg  reservedFreeList1_33; // @[decode.scala 322:30]
  reg  reservedFreeList1_34; // @[decode.scala 322:30]
  reg  reservedFreeList1_35; // @[decode.scala 322:30]
  reg  reservedFreeList1_36; // @[decode.scala 322:30]
  reg  reservedFreeList1_37; // @[decode.scala 322:30]
  reg  reservedFreeList1_38; // @[decode.scala 322:30]
  reg  reservedFreeList1_39; // @[decode.scala 322:30]
  reg  reservedFreeList1_40; // @[decode.scala 322:30]
  reg  reservedFreeList1_41; // @[decode.scala 322:30]
  reg  reservedFreeList1_42; // @[decode.scala 322:30]
  reg  reservedFreeList1_43; // @[decode.scala 322:30]
  reg  reservedFreeList1_44; // @[decode.scala 322:30]
  reg  reservedFreeList1_45; // @[decode.scala 322:30]
  reg  reservedFreeList1_46; // @[decode.scala 322:30]
  reg  reservedFreeList1_47; // @[decode.scala 322:30]
  reg  reservedFreeList1_48; // @[decode.scala 322:30]
  reg  reservedFreeList1_49; // @[decode.scala 322:30]
  reg  reservedFreeList1_50; // @[decode.scala 322:30]
  reg  reservedFreeList1_51; // @[decode.scala 322:30]
  reg  reservedFreeList1_52; // @[decode.scala 322:30]
  reg  reservedFreeList1_53; // @[decode.scala 322:30]
  reg  reservedFreeList1_54; // @[decode.scala 322:30]
  reg  reservedFreeList1_55; // @[decode.scala 322:30]
  reg  reservedFreeList1_56; // @[decode.scala 322:30]
  reg  reservedFreeList1_57; // @[decode.scala 322:30]
  reg  reservedFreeList1_58; // @[decode.scala 322:30]
  reg  reservedFreeList1_59; // @[decode.scala 322:30]
  reg  reservedFreeList1_60; // @[decode.scala 322:30]
  reg  reservedFreeList1_61; // @[decode.scala 322:30]
  reg  reservedFreeList1_62; // @[decode.scala 322:30]
  reg  reservedFreeList2_0; // @[decode.scala 323:30]
  reg  reservedFreeList2_1; // @[decode.scala 323:30]
  reg  reservedFreeList2_2; // @[decode.scala 323:30]
  reg  reservedFreeList2_3; // @[decode.scala 323:30]
  reg  reservedFreeList2_4; // @[decode.scala 323:30]
  reg  reservedFreeList2_5; // @[decode.scala 323:30]
  reg  reservedFreeList2_6; // @[decode.scala 323:30]
  reg  reservedFreeList2_7; // @[decode.scala 323:30]
  reg  reservedFreeList2_8; // @[decode.scala 323:30]
  reg  reservedFreeList2_9; // @[decode.scala 323:30]
  reg  reservedFreeList2_10; // @[decode.scala 323:30]
  reg  reservedFreeList2_11; // @[decode.scala 323:30]
  reg  reservedFreeList2_12; // @[decode.scala 323:30]
  reg  reservedFreeList2_13; // @[decode.scala 323:30]
  reg  reservedFreeList2_14; // @[decode.scala 323:30]
  reg  reservedFreeList2_15; // @[decode.scala 323:30]
  reg  reservedFreeList2_16; // @[decode.scala 323:30]
  reg  reservedFreeList2_17; // @[decode.scala 323:30]
  reg  reservedFreeList2_18; // @[decode.scala 323:30]
  reg  reservedFreeList2_19; // @[decode.scala 323:30]
  reg  reservedFreeList2_20; // @[decode.scala 323:30]
  reg  reservedFreeList2_21; // @[decode.scala 323:30]
  reg  reservedFreeList2_22; // @[decode.scala 323:30]
  reg  reservedFreeList2_23; // @[decode.scala 323:30]
  reg  reservedFreeList2_24; // @[decode.scala 323:30]
  reg  reservedFreeList2_25; // @[decode.scala 323:30]
  reg  reservedFreeList2_26; // @[decode.scala 323:30]
  reg  reservedFreeList2_27; // @[decode.scala 323:30]
  reg  reservedFreeList2_28; // @[decode.scala 323:30]
  reg  reservedFreeList2_29; // @[decode.scala 323:30]
  reg  reservedFreeList2_30; // @[decode.scala 323:30]
  reg  reservedFreeList2_31; // @[decode.scala 323:30]
  reg  reservedFreeList2_32; // @[decode.scala 323:30]
  reg  reservedFreeList2_33; // @[decode.scala 323:30]
  reg  reservedFreeList2_34; // @[decode.scala 323:30]
  reg  reservedFreeList2_35; // @[decode.scala 323:30]
  reg  reservedFreeList2_36; // @[decode.scala 323:30]
  reg  reservedFreeList2_37; // @[decode.scala 323:30]
  reg  reservedFreeList2_38; // @[decode.scala 323:30]
  reg  reservedFreeList2_39; // @[decode.scala 323:30]
  reg  reservedFreeList2_40; // @[decode.scala 323:30]
  reg  reservedFreeList2_41; // @[decode.scala 323:30]
  reg  reservedFreeList2_42; // @[decode.scala 323:30]
  reg  reservedFreeList2_43; // @[decode.scala 323:30]
  reg  reservedFreeList2_44; // @[decode.scala 323:30]
  reg  reservedFreeList2_45; // @[decode.scala 323:30]
  reg  reservedFreeList2_46; // @[decode.scala 323:30]
  reg  reservedFreeList2_47; // @[decode.scala 323:30]
  reg  reservedFreeList2_48; // @[decode.scala 323:30]
  reg  reservedFreeList2_49; // @[decode.scala 323:30]
  reg  reservedFreeList2_50; // @[decode.scala 323:30]
  reg  reservedFreeList2_51; // @[decode.scala 323:30]
  reg  reservedFreeList2_52; // @[decode.scala 323:30]
  reg  reservedFreeList2_53; // @[decode.scala 323:30]
  reg  reservedFreeList2_54; // @[decode.scala 323:30]
  reg  reservedFreeList2_55; // @[decode.scala 323:30]
  reg  reservedFreeList2_56; // @[decode.scala 323:30]
  reg  reservedFreeList2_57; // @[decode.scala 323:30]
  reg  reservedFreeList2_58; // @[decode.scala 323:30]
  reg  reservedFreeList2_59; // @[decode.scala 323:30]
  reg  reservedFreeList2_60; // @[decode.scala 323:30]
  reg  reservedFreeList2_61; // @[decode.scala 323:30]
  reg  reservedFreeList2_62; // @[decode.scala 323:30]
  reg  reservedFreeList3_0; // @[decode.scala 324:30]
  reg  reservedFreeList3_1; // @[decode.scala 324:30]
  reg  reservedFreeList3_2; // @[decode.scala 324:30]
  reg  reservedFreeList3_3; // @[decode.scala 324:30]
  reg  reservedFreeList3_4; // @[decode.scala 324:30]
  reg  reservedFreeList3_5; // @[decode.scala 324:30]
  reg  reservedFreeList3_6; // @[decode.scala 324:30]
  reg  reservedFreeList3_7; // @[decode.scala 324:30]
  reg  reservedFreeList3_8; // @[decode.scala 324:30]
  reg  reservedFreeList3_9; // @[decode.scala 324:30]
  reg  reservedFreeList3_10; // @[decode.scala 324:30]
  reg  reservedFreeList3_11; // @[decode.scala 324:30]
  reg  reservedFreeList3_12; // @[decode.scala 324:30]
  reg  reservedFreeList3_13; // @[decode.scala 324:30]
  reg  reservedFreeList3_14; // @[decode.scala 324:30]
  reg  reservedFreeList3_15; // @[decode.scala 324:30]
  reg  reservedFreeList3_16; // @[decode.scala 324:30]
  reg  reservedFreeList3_17; // @[decode.scala 324:30]
  reg  reservedFreeList3_18; // @[decode.scala 324:30]
  reg  reservedFreeList3_19; // @[decode.scala 324:30]
  reg  reservedFreeList3_20; // @[decode.scala 324:30]
  reg  reservedFreeList3_21; // @[decode.scala 324:30]
  reg  reservedFreeList3_22; // @[decode.scala 324:30]
  reg  reservedFreeList3_23; // @[decode.scala 324:30]
  reg  reservedFreeList3_24; // @[decode.scala 324:30]
  reg  reservedFreeList3_25; // @[decode.scala 324:30]
  reg  reservedFreeList3_26; // @[decode.scala 324:30]
  reg  reservedFreeList3_27; // @[decode.scala 324:30]
  reg  reservedFreeList3_28; // @[decode.scala 324:30]
  reg  reservedFreeList3_29; // @[decode.scala 324:30]
  reg  reservedFreeList3_30; // @[decode.scala 324:30]
  reg  reservedFreeList3_31; // @[decode.scala 324:30]
  reg  reservedFreeList3_32; // @[decode.scala 324:30]
  reg  reservedFreeList3_33; // @[decode.scala 324:30]
  reg  reservedFreeList3_34; // @[decode.scala 324:30]
  reg  reservedFreeList3_35; // @[decode.scala 324:30]
  reg  reservedFreeList3_36; // @[decode.scala 324:30]
  reg  reservedFreeList3_37; // @[decode.scala 324:30]
  reg  reservedFreeList3_38; // @[decode.scala 324:30]
  reg  reservedFreeList3_39; // @[decode.scala 324:30]
  reg  reservedFreeList3_40; // @[decode.scala 324:30]
  reg  reservedFreeList3_41; // @[decode.scala 324:30]
  reg  reservedFreeList3_42; // @[decode.scala 324:30]
  reg  reservedFreeList3_43; // @[decode.scala 324:30]
  reg  reservedFreeList3_44; // @[decode.scala 324:30]
  reg  reservedFreeList3_45; // @[decode.scala 324:30]
  reg  reservedFreeList3_46; // @[decode.scala 324:30]
  reg  reservedFreeList3_47; // @[decode.scala 324:30]
  reg  reservedFreeList3_48; // @[decode.scala 324:30]
  reg  reservedFreeList3_49; // @[decode.scala 324:30]
  reg  reservedFreeList3_50; // @[decode.scala 324:30]
  reg  reservedFreeList3_51; // @[decode.scala 324:30]
  reg  reservedFreeList3_52; // @[decode.scala 324:30]
  reg  reservedFreeList3_53; // @[decode.scala 324:30]
  reg  reservedFreeList3_54; // @[decode.scala 324:30]
  reg  reservedFreeList3_55; // @[decode.scala 324:30]
  reg  reservedFreeList3_56; // @[decode.scala 324:30]
  reg  reservedFreeList3_57; // @[decode.scala 324:30]
  reg  reservedFreeList3_58; // @[decode.scala 324:30]
  reg  reservedFreeList3_59; // @[decode.scala 324:30]
  reg  reservedFreeList3_60; // @[decode.scala 324:30]
  reg  reservedFreeList3_61; // @[decode.scala 324:30]
  reg  reservedFreeList3_62; // @[decode.scala 324:30]
  reg  reservedFreeList4_0; // @[decode.scala 325:30]
  reg  reservedFreeList4_1; // @[decode.scala 325:30]
  reg  reservedFreeList4_2; // @[decode.scala 325:30]
  reg  reservedFreeList4_3; // @[decode.scala 325:30]
  reg  reservedFreeList4_4; // @[decode.scala 325:30]
  reg  reservedFreeList4_5; // @[decode.scala 325:30]
  reg  reservedFreeList4_6; // @[decode.scala 325:30]
  reg  reservedFreeList4_7; // @[decode.scala 325:30]
  reg  reservedFreeList4_8; // @[decode.scala 325:30]
  reg  reservedFreeList4_9; // @[decode.scala 325:30]
  reg  reservedFreeList4_10; // @[decode.scala 325:30]
  reg  reservedFreeList4_11; // @[decode.scala 325:30]
  reg  reservedFreeList4_12; // @[decode.scala 325:30]
  reg  reservedFreeList4_13; // @[decode.scala 325:30]
  reg  reservedFreeList4_14; // @[decode.scala 325:30]
  reg  reservedFreeList4_15; // @[decode.scala 325:30]
  reg  reservedFreeList4_16; // @[decode.scala 325:30]
  reg  reservedFreeList4_17; // @[decode.scala 325:30]
  reg  reservedFreeList4_18; // @[decode.scala 325:30]
  reg  reservedFreeList4_19; // @[decode.scala 325:30]
  reg  reservedFreeList4_20; // @[decode.scala 325:30]
  reg  reservedFreeList4_21; // @[decode.scala 325:30]
  reg  reservedFreeList4_22; // @[decode.scala 325:30]
  reg  reservedFreeList4_23; // @[decode.scala 325:30]
  reg  reservedFreeList4_24; // @[decode.scala 325:30]
  reg  reservedFreeList4_25; // @[decode.scala 325:30]
  reg  reservedFreeList4_26; // @[decode.scala 325:30]
  reg  reservedFreeList4_27; // @[decode.scala 325:30]
  reg  reservedFreeList4_28; // @[decode.scala 325:30]
  reg  reservedFreeList4_29; // @[decode.scala 325:30]
  reg  reservedFreeList4_30; // @[decode.scala 325:30]
  reg  reservedFreeList4_31; // @[decode.scala 325:30]
  reg  reservedFreeList4_32; // @[decode.scala 325:30]
  reg  reservedFreeList4_33; // @[decode.scala 325:30]
  reg  reservedFreeList4_34; // @[decode.scala 325:30]
  reg  reservedFreeList4_35; // @[decode.scala 325:30]
  reg  reservedFreeList4_36; // @[decode.scala 325:30]
  reg  reservedFreeList4_37; // @[decode.scala 325:30]
  reg  reservedFreeList4_38; // @[decode.scala 325:30]
  reg  reservedFreeList4_39; // @[decode.scala 325:30]
  reg  reservedFreeList4_40; // @[decode.scala 325:30]
  reg  reservedFreeList4_41; // @[decode.scala 325:30]
  reg  reservedFreeList4_42; // @[decode.scala 325:30]
  reg  reservedFreeList4_43; // @[decode.scala 325:30]
  reg  reservedFreeList4_44; // @[decode.scala 325:30]
  reg  reservedFreeList4_45; // @[decode.scala 325:30]
  reg  reservedFreeList4_46; // @[decode.scala 325:30]
  reg  reservedFreeList4_47; // @[decode.scala 325:30]
  reg  reservedFreeList4_48; // @[decode.scala 325:30]
  reg  reservedFreeList4_49; // @[decode.scala 325:30]
  reg  reservedFreeList4_50; // @[decode.scala 325:30]
  reg  reservedFreeList4_51; // @[decode.scala 325:30]
  reg  reservedFreeList4_52; // @[decode.scala 325:30]
  reg  reservedFreeList4_53; // @[decode.scala 325:30]
  reg  reservedFreeList4_54; // @[decode.scala 325:30]
  reg  reservedFreeList4_55; // @[decode.scala 325:30]
  reg  reservedFreeList4_56; // @[decode.scala 325:30]
  reg  reservedFreeList4_57; // @[decode.scala 325:30]
  reg  reservedFreeList4_58; // @[decode.scala 325:30]
  reg  reservedFreeList4_59; // @[decode.scala 325:30]
  reg  reservedFreeList4_60; // @[decode.scala 325:30]
  reg  reservedFreeList4_61; // @[decode.scala 325:30]
  reg  reservedFreeList4_62; // @[decode.scala 325:30]
  reg  reservedValidList1_0; // @[decode.scala 327:31]
  reg  reservedValidList1_1; // @[decode.scala 327:31]
  reg  reservedValidList1_2; // @[decode.scala 327:31]
  reg  reservedValidList1_3; // @[decode.scala 327:31]
  reg  reservedValidList1_4; // @[decode.scala 327:31]
  reg  reservedValidList1_5; // @[decode.scala 327:31]
  reg  reservedValidList1_6; // @[decode.scala 327:31]
  reg  reservedValidList1_7; // @[decode.scala 327:31]
  reg  reservedValidList1_8; // @[decode.scala 327:31]
  reg  reservedValidList1_9; // @[decode.scala 327:31]
  reg  reservedValidList1_10; // @[decode.scala 327:31]
  reg  reservedValidList1_11; // @[decode.scala 327:31]
  reg  reservedValidList1_12; // @[decode.scala 327:31]
  reg  reservedValidList1_13; // @[decode.scala 327:31]
  reg  reservedValidList1_14; // @[decode.scala 327:31]
  reg  reservedValidList1_15; // @[decode.scala 327:31]
  reg  reservedValidList1_16; // @[decode.scala 327:31]
  reg  reservedValidList1_17; // @[decode.scala 327:31]
  reg  reservedValidList1_18; // @[decode.scala 327:31]
  reg  reservedValidList1_19; // @[decode.scala 327:31]
  reg  reservedValidList1_20; // @[decode.scala 327:31]
  reg  reservedValidList1_21; // @[decode.scala 327:31]
  reg  reservedValidList1_22; // @[decode.scala 327:31]
  reg  reservedValidList1_23; // @[decode.scala 327:31]
  reg  reservedValidList1_24; // @[decode.scala 327:31]
  reg  reservedValidList1_25; // @[decode.scala 327:31]
  reg  reservedValidList1_26; // @[decode.scala 327:31]
  reg  reservedValidList1_27; // @[decode.scala 327:31]
  reg  reservedValidList1_28; // @[decode.scala 327:31]
  reg  reservedValidList1_29; // @[decode.scala 327:31]
  reg  reservedValidList1_30; // @[decode.scala 327:31]
  reg  reservedValidList1_31; // @[decode.scala 327:31]
  reg  reservedValidList1_32; // @[decode.scala 327:31]
  reg  reservedValidList1_33; // @[decode.scala 327:31]
  reg  reservedValidList1_34; // @[decode.scala 327:31]
  reg  reservedValidList1_35; // @[decode.scala 327:31]
  reg  reservedValidList1_36; // @[decode.scala 327:31]
  reg  reservedValidList1_37; // @[decode.scala 327:31]
  reg  reservedValidList1_38; // @[decode.scala 327:31]
  reg  reservedValidList1_39; // @[decode.scala 327:31]
  reg  reservedValidList1_40; // @[decode.scala 327:31]
  reg  reservedValidList1_41; // @[decode.scala 327:31]
  reg  reservedValidList1_42; // @[decode.scala 327:31]
  reg  reservedValidList1_43; // @[decode.scala 327:31]
  reg  reservedValidList1_44; // @[decode.scala 327:31]
  reg  reservedValidList1_45; // @[decode.scala 327:31]
  reg  reservedValidList1_46; // @[decode.scala 327:31]
  reg  reservedValidList1_47; // @[decode.scala 327:31]
  reg  reservedValidList1_48; // @[decode.scala 327:31]
  reg  reservedValidList1_49; // @[decode.scala 327:31]
  reg  reservedValidList1_50; // @[decode.scala 327:31]
  reg  reservedValidList1_51; // @[decode.scala 327:31]
  reg  reservedValidList1_52; // @[decode.scala 327:31]
  reg  reservedValidList1_53; // @[decode.scala 327:31]
  reg  reservedValidList1_54; // @[decode.scala 327:31]
  reg  reservedValidList1_55; // @[decode.scala 327:31]
  reg  reservedValidList1_56; // @[decode.scala 327:31]
  reg  reservedValidList1_57; // @[decode.scala 327:31]
  reg  reservedValidList1_58; // @[decode.scala 327:31]
  reg  reservedValidList1_59; // @[decode.scala 327:31]
  reg  reservedValidList1_60; // @[decode.scala 327:31]
  reg  reservedValidList1_61; // @[decode.scala 327:31]
  reg  reservedValidList1_62; // @[decode.scala 327:31]
  reg  reservedValidList1_63; // @[decode.scala 327:31]
  reg  reservedValidList2_0; // @[decode.scala 328:31]
  reg  reservedValidList2_1; // @[decode.scala 328:31]
  reg  reservedValidList2_2; // @[decode.scala 328:31]
  reg  reservedValidList2_3; // @[decode.scala 328:31]
  reg  reservedValidList2_4; // @[decode.scala 328:31]
  reg  reservedValidList2_5; // @[decode.scala 328:31]
  reg  reservedValidList2_6; // @[decode.scala 328:31]
  reg  reservedValidList2_7; // @[decode.scala 328:31]
  reg  reservedValidList2_8; // @[decode.scala 328:31]
  reg  reservedValidList2_9; // @[decode.scala 328:31]
  reg  reservedValidList2_10; // @[decode.scala 328:31]
  reg  reservedValidList2_11; // @[decode.scala 328:31]
  reg  reservedValidList2_12; // @[decode.scala 328:31]
  reg  reservedValidList2_13; // @[decode.scala 328:31]
  reg  reservedValidList2_14; // @[decode.scala 328:31]
  reg  reservedValidList2_15; // @[decode.scala 328:31]
  reg  reservedValidList2_16; // @[decode.scala 328:31]
  reg  reservedValidList2_17; // @[decode.scala 328:31]
  reg  reservedValidList2_18; // @[decode.scala 328:31]
  reg  reservedValidList2_19; // @[decode.scala 328:31]
  reg  reservedValidList2_20; // @[decode.scala 328:31]
  reg  reservedValidList2_21; // @[decode.scala 328:31]
  reg  reservedValidList2_22; // @[decode.scala 328:31]
  reg  reservedValidList2_23; // @[decode.scala 328:31]
  reg  reservedValidList2_24; // @[decode.scala 328:31]
  reg  reservedValidList2_25; // @[decode.scala 328:31]
  reg  reservedValidList2_26; // @[decode.scala 328:31]
  reg  reservedValidList2_27; // @[decode.scala 328:31]
  reg  reservedValidList2_28; // @[decode.scala 328:31]
  reg  reservedValidList2_29; // @[decode.scala 328:31]
  reg  reservedValidList2_30; // @[decode.scala 328:31]
  reg  reservedValidList2_31; // @[decode.scala 328:31]
  reg  reservedValidList2_32; // @[decode.scala 328:31]
  reg  reservedValidList2_33; // @[decode.scala 328:31]
  reg  reservedValidList2_34; // @[decode.scala 328:31]
  reg  reservedValidList2_35; // @[decode.scala 328:31]
  reg  reservedValidList2_36; // @[decode.scala 328:31]
  reg  reservedValidList2_37; // @[decode.scala 328:31]
  reg  reservedValidList2_38; // @[decode.scala 328:31]
  reg  reservedValidList2_39; // @[decode.scala 328:31]
  reg  reservedValidList2_40; // @[decode.scala 328:31]
  reg  reservedValidList2_41; // @[decode.scala 328:31]
  reg  reservedValidList2_42; // @[decode.scala 328:31]
  reg  reservedValidList2_43; // @[decode.scala 328:31]
  reg  reservedValidList2_44; // @[decode.scala 328:31]
  reg  reservedValidList2_45; // @[decode.scala 328:31]
  reg  reservedValidList2_46; // @[decode.scala 328:31]
  reg  reservedValidList2_47; // @[decode.scala 328:31]
  reg  reservedValidList2_48; // @[decode.scala 328:31]
  reg  reservedValidList2_49; // @[decode.scala 328:31]
  reg  reservedValidList2_50; // @[decode.scala 328:31]
  reg  reservedValidList2_51; // @[decode.scala 328:31]
  reg  reservedValidList2_52; // @[decode.scala 328:31]
  reg  reservedValidList2_53; // @[decode.scala 328:31]
  reg  reservedValidList2_54; // @[decode.scala 328:31]
  reg  reservedValidList2_55; // @[decode.scala 328:31]
  reg  reservedValidList2_56; // @[decode.scala 328:31]
  reg  reservedValidList2_57; // @[decode.scala 328:31]
  reg  reservedValidList2_58; // @[decode.scala 328:31]
  reg  reservedValidList2_59; // @[decode.scala 328:31]
  reg  reservedValidList2_60; // @[decode.scala 328:31]
  reg  reservedValidList2_61; // @[decode.scala 328:31]
  reg  reservedValidList2_62; // @[decode.scala 328:31]
  reg  reservedValidList2_63; // @[decode.scala 328:31]
  reg  reservedValidList3_0; // @[decode.scala 329:31]
  reg  reservedValidList3_1; // @[decode.scala 329:31]
  reg  reservedValidList3_2; // @[decode.scala 329:31]
  reg  reservedValidList3_3; // @[decode.scala 329:31]
  reg  reservedValidList3_4; // @[decode.scala 329:31]
  reg  reservedValidList3_5; // @[decode.scala 329:31]
  reg  reservedValidList3_6; // @[decode.scala 329:31]
  reg  reservedValidList3_7; // @[decode.scala 329:31]
  reg  reservedValidList3_8; // @[decode.scala 329:31]
  reg  reservedValidList3_9; // @[decode.scala 329:31]
  reg  reservedValidList3_10; // @[decode.scala 329:31]
  reg  reservedValidList3_11; // @[decode.scala 329:31]
  reg  reservedValidList3_12; // @[decode.scala 329:31]
  reg  reservedValidList3_13; // @[decode.scala 329:31]
  reg  reservedValidList3_14; // @[decode.scala 329:31]
  reg  reservedValidList3_15; // @[decode.scala 329:31]
  reg  reservedValidList3_16; // @[decode.scala 329:31]
  reg  reservedValidList3_17; // @[decode.scala 329:31]
  reg  reservedValidList3_18; // @[decode.scala 329:31]
  reg  reservedValidList3_19; // @[decode.scala 329:31]
  reg  reservedValidList3_20; // @[decode.scala 329:31]
  reg  reservedValidList3_21; // @[decode.scala 329:31]
  reg  reservedValidList3_22; // @[decode.scala 329:31]
  reg  reservedValidList3_23; // @[decode.scala 329:31]
  reg  reservedValidList3_24; // @[decode.scala 329:31]
  reg  reservedValidList3_25; // @[decode.scala 329:31]
  reg  reservedValidList3_26; // @[decode.scala 329:31]
  reg  reservedValidList3_27; // @[decode.scala 329:31]
  reg  reservedValidList3_28; // @[decode.scala 329:31]
  reg  reservedValidList3_29; // @[decode.scala 329:31]
  reg  reservedValidList3_30; // @[decode.scala 329:31]
  reg  reservedValidList3_31; // @[decode.scala 329:31]
  reg  reservedValidList3_32; // @[decode.scala 329:31]
  reg  reservedValidList3_33; // @[decode.scala 329:31]
  reg  reservedValidList3_34; // @[decode.scala 329:31]
  reg  reservedValidList3_35; // @[decode.scala 329:31]
  reg  reservedValidList3_36; // @[decode.scala 329:31]
  reg  reservedValidList3_37; // @[decode.scala 329:31]
  reg  reservedValidList3_38; // @[decode.scala 329:31]
  reg  reservedValidList3_39; // @[decode.scala 329:31]
  reg  reservedValidList3_40; // @[decode.scala 329:31]
  reg  reservedValidList3_41; // @[decode.scala 329:31]
  reg  reservedValidList3_42; // @[decode.scala 329:31]
  reg  reservedValidList3_43; // @[decode.scala 329:31]
  reg  reservedValidList3_44; // @[decode.scala 329:31]
  reg  reservedValidList3_45; // @[decode.scala 329:31]
  reg  reservedValidList3_46; // @[decode.scala 329:31]
  reg  reservedValidList3_47; // @[decode.scala 329:31]
  reg  reservedValidList3_48; // @[decode.scala 329:31]
  reg  reservedValidList3_49; // @[decode.scala 329:31]
  reg  reservedValidList3_50; // @[decode.scala 329:31]
  reg  reservedValidList3_51; // @[decode.scala 329:31]
  reg  reservedValidList3_52; // @[decode.scala 329:31]
  reg  reservedValidList3_53; // @[decode.scala 329:31]
  reg  reservedValidList3_54; // @[decode.scala 329:31]
  reg  reservedValidList3_55; // @[decode.scala 329:31]
  reg  reservedValidList3_56; // @[decode.scala 329:31]
  reg  reservedValidList3_57; // @[decode.scala 329:31]
  reg  reservedValidList3_58; // @[decode.scala 329:31]
  reg  reservedValidList3_59; // @[decode.scala 329:31]
  reg  reservedValidList3_60; // @[decode.scala 329:31]
  reg  reservedValidList3_61; // @[decode.scala 329:31]
  reg  reservedValidList3_62; // @[decode.scala 329:31]
  reg  reservedValidList3_63; // @[decode.scala 329:31]
  reg  reservedValidList4_0; // @[decode.scala 330:31]
  reg  reservedValidList4_1; // @[decode.scala 330:31]
  reg  reservedValidList4_2; // @[decode.scala 330:31]
  reg  reservedValidList4_3; // @[decode.scala 330:31]
  reg  reservedValidList4_4; // @[decode.scala 330:31]
  reg  reservedValidList4_5; // @[decode.scala 330:31]
  reg  reservedValidList4_6; // @[decode.scala 330:31]
  reg  reservedValidList4_7; // @[decode.scala 330:31]
  reg  reservedValidList4_8; // @[decode.scala 330:31]
  reg  reservedValidList4_9; // @[decode.scala 330:31]
  reg  reservedValidList4_10; // @[decode.scala 330:31]
  reg  reservedValidList4_11; // @[decode.scala 330:31]
  reg  reservedValidList4_12; // @[decode.scala 330:31]
  reg  reservedValidList4_13; // @[decode.scala 330:31]
  reg  reservedValidList4_14; // @[decode.scala 330:31]
  reg  reservedValidList4_15; // @[decode.scala 330:31]
  reg  reservedValidList4_16; // @[decode.scala 330:31]
  reg  reservedValidList4_17; // @[decode.scala 330:31]
  reg  reservedValidList4_18; // @[decode.scala 330:31]
  reg  reservedValidList4_19; // @[decode.scala 330:31]
  reg  reservedValidList4_20; // @[decode.scala 330:31]
  reg  reservedValidList4_21; // @[decode.scala 330:31]
  reg  reservedValidList4_22; // @[decode.scala 330:31]
  reg  reservedValidList4_23; // @[decode.scala 330:31]
  reg  reservedValidList4_24; // @[decode.scala 330:31]
  reg  reservedValidList4_25; // @[decode.scala 330:31]
  reg  reservedValidList4_26; // @[decode.scala 330:31]
  reg  reservedValidList4_27; // @[decode.scala 330:31]
  reg  reservedValidList4_28; // @[decode.scala 330:31]
  reg  reservedValidList4_29; // @[decode.scala 330:31]
  reg  reservedValidList4_30; // @[decode.scala 330:31]
  reg  reservedValidList4_31; // @[decode.scala 330:31]
  reg  reservedValidList4_32; // @[decode.scala 330:31]
  reg  reservedValidList4_33; // @[decode.scala 330:31]
  reg  reservedValidList4_34; // @[decode.scala 330:31]
  reg  reservedValidList4_35; // @[decode.scala 330:31]
  reg  reservedValidList4_36; // @[decode.scala 330:31]
  reg  reservedValidList4_37; // @[decode.scala 330:31]
  reg  reservedValidList4_38; // @[decode.scala 330:31]
  reg  reservedValidList4_39; // @[decode.scala 330:31]
  reg  reservedValidList4_40; // @[decode.scala 330:31]
  reg  reservedValidList4_41; // @[decode.scala 330:31]
  reg  reservedValidList4_42; // @[decode.scala 330:31]
  reg  reservedValidList4_43; // @[decode.scala 330:31]
  reg  reservedValidList4_44; // @[decode.scala 330:31]
  reg  reservedValidList4_45; // @[decode.scala 330:31]
  reg  reservedValidList4_46; // @[decode.scala 330:31]
  reg  reservedValidList4_47; // @[decode.scala 330:31]
  reg  reservedValidList4_48; // @[decode.scala 330:31]
  reg  reservedValidList4_49; // @[decode.scala 330:31]
  reg  reservedValidList4_50; // @[decode.scala 330:31]
  reg  reservedValidList4_51; // @[decode.scala 330:31]
  reg  reservedValidList4_52; // @[decode.scala 330:31]
  reg  reservedValidList4_53; // @[decode.scala 330:31]
  reg  reservedValidList4_54; // @[decode.scala 330:31]
  reg  reservedValidList4_55; // @[decode.scala 330:31]
  reg  reservedValidList4_56; // @[decode.scala 330:31]
  reg  reservedValidList4_57; // @[decode.scala 330:31]
  reg  reservedValidList4_58; // @[decode.scala 330:31]
  reg  reservedValidList4_59; // @[decode.scala 330:31]
  reg  reservedValidList4_60; // @[decode.scala 330:31]
  reg  reservedValidList4_61; // @[decode.scala 330:31]
  reg  reservedValidList4_62; // @[decode.scala 330:31]
  reg  reservedValidList4_63; // @[decode.scala 330:31]
  wire  _GEN_273 = 6'h0 == rs1Addr ? 1'h0 : PRFFreeList_0; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_274 = 6'h1 == rs1Addr ? 1'h0 : PRFFreeList_1; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_275 = 6'h2 == rs1Addr ? 1'h0 : PRFFreeList_2; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_276 = 6'h3 == rs1Addr ? 1'h0 : PRFFreeList_3; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_277 = 6'h4 == rs1Addr ? 1'h0 : PRFFreeList_4; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_278 = 6'h5 == rs1Addr ? 1'h0 : PRFFreeList_5; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_279 = 6'h6 == rs1Addr ? 1'h0 : PRFFreeList_6; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_280 = 6'h7 == rs1Addr ? 1'h0 : PRFFreeList_7; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_281 = 6'h8 == rs1Addr ? 1'h0 : PRFFreeList_8; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_282 = 6'h9 == rs1Addr ? 1'h0 : PRFFreeList_9; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_283 = 6'ha == rs1Addr ? 1'h0 : PRFFreeList_10; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_284 = 6'hb == rs1Addr ? 1'h0 : PRFFreeList_11; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_285 = 6'hc == rs1Addr ? 1'h0 : PRFFreeList_12; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_286 = 6'hd == rs1Addr ? 1'h0 : PRFFreeList_13; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_287 = 6'he == rs1Addr ? 1'h0 : PRFFreeList_14; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_288 = 6'hf == rs1Addr ? 1'h0 : PRFFreeList_15; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_289 = 6'h10 == rs1Addr ? 1'h0 : PRFFreeList_16; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_290 = 6'h11 == rs1Addr ? 1'h0 : PRFFreeList_17; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_291 = 6'h12 == rs1Addr ? 1'h0 : PRFFreeList_18; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_292 = 6'h13 == rs1Addr ? 1'h0 : PRFFreeList_19; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_293 = 6'h14 == rs1Addr ? 1'h0 : PRFFreeList_20; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_294 = 6'h15 == rs1Addr ? 1'h0 : PRFFreeList_21; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_295 = 6'h16 == rs1Addr ? 1'h0 : PRFFreeList_22; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_296 = 6'h17 == rs1Addr ? 1'h0 : PRFFreeList_23; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_297 = 6'h18 == rs1Addr ? 1'h0 : PRFFreeList_24; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_298 = 6'h19 == rs1Addr ? 1'h0 : PRFFreeList_25; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_299 = 6'h1a == rs1Addr ? 1'h0 : PRFFreeList_26; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_300 = 6'h1b == rs1Addr ? 1'h0 : PRFFreeList_27; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_301 = 6'h1c == rs1Addr ? 1'h0 : PRFFreeList_28; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_302 = 6'h1d == rs1Addr ? 1'h0 : PRFFreeList_29; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_303 = 6'h1e == rs1Addr ? 1'h0 : PRFFreeList_30; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_304 = 6'h1f == rs1Addr ? 1'h0 : PRFFreeList_31; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_305 = 6'h20 == rs1Addr ? 1'h0 : PRFFreeList_32; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_306 = 6'h21 == rs1Addr ? 1'h0 : PRFFreeList_33; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_307 = 6'h22 == rs1Addr ? 1'h0 : PRFFreeList_34; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_308 = 6'h23 == rs1Addr ? 1'h0 : PRFFreeList_35; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_309 = 6'h24 == rs1Addr ? 1'h0 : PRFFreeList_36; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_310 = 6'h25 == rs1Addr ? 1'h0 : PRFFreeList_37; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_311 = 6'h26 == rs1Addr ? 1'h0 : PRFFreeList_38; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_312 = 6'h27 == rs1Addr ? 1'h0 : PRFFreeList_39; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_313 = 6'h28 == rs1Addr ? 1'h0 : PRFFreeList_40; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_314 = 6'h29 == rs1Addr ? 1'h0 : PRFFreeList_41; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_315 = 6'h2a == rs1Addr ? 1'h0 : PRFFreeList_42; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_316 = 6'h2b == rs1Addr ? 1'h0 : PRFFreeList_43; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_317 = 6'h2c == rs1Addr ? 1'h0 : PRFFreeList_44; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_318 = 6'h2d == rs1Addr ? 1'h0 : PRFFreeList_45; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_319 = 6'h2e == rs1Addr ? 1'h0 : PRFFreeList_46; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_320 = 6'h2f == rs1Addr ? 1'h0 : PRFFreeList_47; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_321 = 6'h30 == rs1Addr ? 1'h0 : PRFFreeList_48; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_322 = 6'h31 == rs1Addr ? 1'h0 : PRFFreeList_49; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_323 = 6'h32 == rs1Addr ? 1'h0 : PRFFreeList_50; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_324 = 6'h33 == rs1Addr ? 1'h0 : PRFFreeList_51; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_325 = 6'h34 == rs1Addr ? 1'h0 : PRFFreeList_52; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_326 = 6'h35 == rs1Addr ? 1'h0 : PRFFreeList_53; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_327 = 6'h36 == rs1Addr ? 1'h0 : PRFFreeList_54; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_328 = 6'h37 == rs1Addr ? 1'h0 : PRFFreeList_55; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_329 = 6'h38 == rs1Addr ? 1'h0 : PRFFreeList_56; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_330 = 6'h39 == rs1Addr ? 1'h0 : PRFFreeList_57; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_331 = 6'h3a == rs1Addr ? 1'h0 : PRFFreeList_58; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_332 = 6'h3b == rs1Addr ? 1'h0 : PRFFreeList_59; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_333 = 6'h3c == rs1Addr ? 1'h0 : PRFFreeList_60; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_334 = 6'h3d == rs1Addr ? 1'h0 : PRFFreeList_61; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_335 = 6'h3e == rs1Addr ? 1'h0 : PRFFreeList_62; // @[decode.scala 345:{28,28} 310:36]
  wire  _GEN_337 = 6'h0 == rs2Addr ? 1'h0 : PRFFreeList_0; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_338 = 6'h1 == rs2Addr ? 1'h0 : PRFFreeList_1; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_339 = 6'h2 == rs2Addr ? 1'h0 : PRFFreeList_2; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_340 = 6'h3 == rs2Addr ? 1'h0 : PRFFreeList_3; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_341 = 6'h4 == rs2Addr ? 1'h0 : PRFFreeList_4; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_342 = 6'h5 == rs2Addr ? 1'h0 : PRFFreeList_5; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_343 = 6'h6 == rs2Addr ? 1'h0 : PRFFreeList_6; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_344 = 6'h7 == rs2Addr ? 1'h0 : PRFFreeList_7; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_345 = 6'h8 == rs2Addr ? 1'h0 : PRFFreeList_8; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_346 = 6'h9 == rs2Addr ? 1'h0 : PRFFreeList_9; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_347 = 6'ha == rs2Addr ? 1'h0 : PRFFreeList_10; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_348 = 6'hb == rs2Addr ? 1'h0 : PRFFreeList_11; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_349 = 6'hc == rs2Addr ? 1'h0 : PRFFreeList_12; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_350 = 6'hd == rs2Addr ? 1'h0 : PRFFreeList_13; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_351 = 6'he == rs2Addr ? 1'h0 : PRFFreeList_14; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_352 = 6'hf == rs2Addr ? 1'h0 : PRFFreeList_15; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_353 = 6'h10 == rs2Addr ? 1'h0 : PRFFreeList_16; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_354 = 6'h11 == rs2Addr ? 1'h0 : PRFFreeList_17; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_355 = 6'h12 == rs2Addr ? 1'h0 : PRFFreeList_18; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_356 = 6'h13 == rs2Addr ? 1'h0 : PRFFreeList_19; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_357 = 6'h14 == rs2Addr ? 1'h0 : PRFFreeList_20; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_358 = 6'h15 == rs2Addr ? 1'h0 : PRFFreeList_21; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_359 = 6'h16 == rs2Addr ? 1'h0 : PRFFreeList_22; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_360 = 6'h17 == rs2Addr ? 1'h0 : PRFFreeList_23; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_361 = 6'h18 == rs2Addr ? 1'h0 : PRFFreeList_24; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_362 = 6'h19 == rs2Addr ? 1'h0 : PRFFreeList_25; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_363 = 6'h1a == rs2Addr ? 1'h0 : PRFFreeList_26; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_364 = 6'h1b == rs2Addr ? 1'h0 : PRFFreeList_27; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_365 = 6'h1c == rs2Addr ? 1'h0 : PRFFreeList_28; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_366 = 6'h1d == rs2Addr ? 1'h0 : PRFFreeList_29; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_367 = 6'h1e == rs2Addr ? 1'h0 : PRFFreeList_30; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_368 = 6'h1f == rs2Addr ? 1'h0 : PRFFreeList_31; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_369 = 6'h20 == rs2Addr ? 1'h0 : PRFFreeList_32; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_370 = 6'h21 == rs2Addr ? 1'h0 : PRFFreeList_33; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_371 = 6'h22 == rs2Addr ? 1'h0 : PRFFreeList_34; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_372 = 6'h23 == rs2Addr ? 1'h0 : PRFFreeList_35; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_373 = 6'h24 == rs2Addr ? 1'h0 : PRFFreeList_36; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_374 = 6'h25 == rs2Addr ? 1'h0 : PRFFreeList_37; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_375 = 6'h26 == rs2Addr ? 1'h0 : PRFFreeList_38; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_376 = 6'h27 == rs2Addr ? 1'h0 : PRFFreeList_39; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_377 = 6'h28 == rs2Addr ? 1'h0 : PRFFreeList_40; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_378 = 6'h29 == rs2Addr ? 1'h0 : PRFFreeList_41; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_379 = 6'h2a == rs2Addr ? 1'h0 : PRFFreeList_42; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_380 = 6'h2b == rs2Addr ? 1'h0 : PRFFreeList_43; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_381 = 6'h2c == rs2Addr ? 1'h0 : PRFFreeList_44; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_382 = 6'h2d == rs2Addr ? 1'h0 : PRFFreeList_45; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_383 = 6'h2e == rs2Addr ? 1'h0 : PRFFreeList_46; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_384 = 6'h2f == rs2Addr ? 1'h0 : PRFFreeList_47; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_385 = 6'h30 == rs2Addr ? 1'h0 : PRFFreeList_48; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_386 = 6'h31 == rs2Addr ? 1'h0 : PRFFreeList_49; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_387 = 6'h32 == rs2Addr ? 1'h0 : PRFFreeList_50; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_388 = 6'h33 == rs2Addr ? 1'h0 : PRFFreeList_51; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_389 = 6'h34 == rs2Addr ? 1'h0 : PRFFreeList_52; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_390 = 6'h35 == rs2Addr ? 1'h0 : PRFFreeList_53; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_391 = 6'h36 == rs2Addr ? 1'h0 : PRFFreeList_54; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_392 = 6'h37 == rs2Addr ? 1'h0 : PRFFreeList_55; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_393 = 6'h38 == rs2Addr ? 1'h0 : PRFFreeList_56; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_394 = 6'h39 == rs2Addr ? 1'h0 : PRFFreeList_57; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_395 = 6'h3a == rs2Addr ? 1'h0 : PRFFreeList_58; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_396 = 6'h3b == rs2Addr ? 1'h0 : PRFFreeList_59; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_397 = 6'h3c == rs2Addr ? 1'h0 : PRFFreeList_60; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_398 = 6'h3d == rs2Addr ? 1'h0 : PRFFreeList_61; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_399 = 6'h3e == rs2Addr ? 1'h0 : PRFFreeList_62; // @[decode.scala 347:{28,28} 310:36]
  wire  _GEN_401 = _T_22 ? _GEN_337 : PRFFreeList_0; // @[decode.scala 310:36 346:41]
  wire  _GEN_402 = _T_22 ? _GEN_338 : PRFFreeList_1; // @[decode.scala 310:36 346:41]
  wire  _GEN_403 = _T_22 ? _GEN_339 : PRFFreeList_2; // @[decode.scala 310:36 346:41]
  wire  _GEN_404 = _T_22 ? _GEN_340 : PRFFreeList_3; // @[decode.scala 310:36 346:41]
  wire  _GEN_405 = _T_22 ? _GEN_341 : PRFFreeList_4; // @[decode.scala 310:36 346:41]
  wire  _GEN_406 = _T_22 ? _GEN_342 : PRFFreeList_5; // @[decode.scala 310:36 346:41]
  wire  _GEN_407 = _T_22 ? _GEN_343 : PRFFreeList_6; // @[decode.scala 310:36 346:41]
  wire  _GEN_408 = _T_22 ? _GEN_344 : PRFFreeList_7; // @[decode.scala 310:36 346:41]
  wire  _GEN_409 = _T_22 ? _GEN_345 : PRFFreeList_8; // @[decode.scala 310:36 346:41]
  wire  _GEN_410 = _T_22 ? _GEN_346 : PRFFreeList_9; // @[decode.scala 310:36 346:41]
  wire  _GEN_411 = _T_22 ? _GEN_347 : PRFFreeList_10; // @[decode.scala 310:36 346:41]
  wire  _GEN_412 = _T_22 ? _GEN_348 : PRFFreeList_11; // @[decode.scala 310:36 346:41]
  wire  _GEN_413 = _T_22 ? _GEN_349 : PRFFreeList_12; // @[decode.scala 310:36 346:41]
  wire  _GEN_414 = _T_22 ? _GEN_350 : PRFFreeList_13; // @[decode.scala 310:36 346:41]
  wire  _GEN_415 = _T_22 ? _GEN_351 : PRFFreeList_14; // @[decode.scala 310:36 346:41]
  wire  _GEN_416 = _T_22 ? _GEN_352 : PRFFreeList_15; // @[decode.scala 310:36 346:41]
  wire  _GEN_417 = _T_22 ? _GEN_353 : PRFFreeList_16; // @[decode.scala 310:36 346:41]
  wire  _GEN_418 = _T_22 ? _GEN_354 : PRFFreeList_17; // @[decode.scala 310:36 346:41]
  wire  _GEN_419 = _T_22 ? _GEN_355 : PRFFreeList_18; // @[decode.scala 310:36 346:41]
  wire  _GEN_420 = _T_22 ? _GEN_356 : PRFFreeList_19; // @[decode.scala 310:36 346:41]
  wire  _GEN_421 = _T_22 ? _GEN_357 : PRFFreeList_20; // @[decode.scala 310:36 346:41]
  wire  _GEN_422 = _T_22 ? _GEN_358 : PRFFreeList_21; // @[decode.scala 310:36 346:41]
  wire  _GEN_423 = _T_22 ? _GEN_359 : PRFFreeList_22; // @[decode.scala 310:36 346:41]
  wire  _GEN_424 = _T_22 ? _GEN_360 : PRFFreeList_23; // @[decode.scala 310:36 346:41]
  wire  _GEN_425 = _T_22 ? _GEN_361 : PRFFreeList_24; // @[decode.scala 310:36 346:41]
  wire  _GEN_426 = _T_22 ? _GEN_362 : PRFFreeList_25; // @[decode.scala 310:36 346:41]
  wire  _GEN_427 = _T_22 ? _GEN_363 : PRFFreeList_26; // @[decode.scala 310:36 346:41]
  wire  _GEN_428 = _T_22 ? _GEN_364 : PRFFreeList_27; // @[decode.scala 310:36 346:41]
  wire  _GEN_429 = _T_22 ? _GEN_365 : PRFFreeList_28; // @[decode.scala 310:36 346:41]
  wire  _GEN_430 = _T_22 ? _GEN_366 : PRFFreeList_29; // @[decode.scala 310:36 346:41]
  wire  _GEN_431 = _T_22 ? _GEN_367 : PRFFreeList_30; // @[decode.scala 310:36 346:41]
  wire  _GEN_432 = _T_22 ? _GEN_368 : PRFFreeList_31; // @[decode.scala 310:36 346:41]
  wire  _GEN_433 = _T_22 ? _GEN_369 : PRFFreeList_32; // @[decode.scala 310:36 346:41]
  wire  _GEN_434 = _T_22 ? _GEN_370 : PRFFreeList_33; // @[decode.scala 310:36 346:41]
  wire  _GEN_435 = _T_22 ? _GEN_371 : PRFFreeList_34; // @[decode.scala 310:36 346:41]
  wire  _GEN_436 = _T_22 ? _GEN_372 : PRFFreeList_35; // @[decode.scala 310:36 346:41]
  wire  _GEN_437 = _T_22 ? _GEN_373 : PRFFreeList_36; // @[decode.scala 310:36 346:41]
  wire  _GEN_438 = _T_22 ? _GEN_374 : PRFFreeList_37; // @[decode.scala 310:36 346:41]
  wire  _GEN_439 = _T_22 ? _GEN_375 : PRFFreeList_38; // @[decode.scala 310:36 346:41]
  wire  _GEN_440 = _T_22 ? _GEN_376 : PRFFreeList_39; // @[decode.scala 310:36 346:41]
  wire  _GEN_441 = _T_22 ? _GEN_377 : PRFFreeList_40; // @[decode.scala 310:36 346:41]
  wire  _GEN_442 = _T_22 ? _GEN_378 : PRFFreeList_41; // @[decode.scala 310:36 346:41]
  wire  _GEN_443 = _T_22 ? _GEN_379 : PRFFreeList_42; // @[decode.scala 310:36 346:41]
  wire  _GEN_444 = _T_22 ? _GEN_380 : PRFFreeList_43; // @[decode.scala 310:36 346:41]
  wire  _GEN_445 = _T_22 ? _GEN_381 : PRFFreeList_44; // @[decode.scala 310:36 346:41]
  wire  _GEN_446 = _T_22 ? _GEN_382 : PRFFreeList_45; // @[decode.scala 310:36 346:41]
  wire  _GEN_447 = _T_22 ? _GEN_383 : PRFFreeList_46; // @[decode.scala 310:36 346:41]
  wire  _GEN_448 = _T_22 ? _GEN_384 : PRFFreeList_47; // @[decode.scala 310:36 346:41]
  wire  _GEN_449 = _T_22 ? _GEN_385 : PRFFreeList_48; // @[decode.scala 310:36 346:41]
  wire  _GEN_450 = _T_22 ? _GEN_386 : PRFFreeList_49; // @[decode.scala 310:36 346:41]
  wire  _GEN_451 = _T_22 ? _GEN_387 : PRFFreeList_50; // @[decode.scala 310:36 346:41]
  wire  _GEN_452 = _T_22 ? _GEN_388 : PRFFreeList_51; // @[decode.scala 310:36 346:41]
  wire  _GEN_453 = _T_22 ? _GEN_389 : PRFFreeList_52; // @[decode.scala 310:36 346:41]
  wire  _GEN_454 = _T_22 ? _GEN_390 : PRFFreeList_53; // @[decode.scala 310:36 346:41]
  wire  _GEN_455 = _T_22 ? _GEN_391 : PRFFreeList_54; // @[decode.scala 310:36 346:41]
  wire  _GEN_456 = _T_22 ? _GEN_392 : PRFFreeList_55; // @[decode.scala 310:36 346:41]
  wire  _GEN_457 = _T_22 ? _GEN_393 : PRFFreeList_56; // @[decode.scala 310:36 346:41]
  wire  _GEN_458 = _T_22 ? _GEN_394 : PRFFreeList_57; // @[decode.scala 310:36 346:41]
  wire  _GEN_459 = _T_22 ? _GEN_395 : PRFFreeList_58; // @[decode.scala 310:36 346:41]
  wire  _GEN_460 = _T_22 ? _GEN_396 : PRFFreeList_59; // @[decode.scala 310:36 346:41]
  wire  _GEN_461 = _T_22 ? _GEN_397 : PRFFreeList_60; // @[decode.scala 310:36 346:41]
  wire  _GEN_462 = _T_22 ? _GEN_398 : PRFFreeList_61; // @[decode.scala 310:36 346:41]
  wire  _GEN_463 = _T_22 ? _GEN_399 : PRFFreeList_62; // @[decode.scala 310:36 346:41]
  wire  _GEN_465 = _T_21 ? _GEN_273 : _GEN_401; // @[decode.scala 344:35]
  wire  _GEN_466 = _T_21 ? _GEN_274 : _GEN_402; // @[decode.scala 344:35]
  wire  _GEN_467 = _T_21 ? _GEN_275 : _GEN_403; // @[decode.scala 344:35]
  wire  _GEN_468 = _T_21 ? _GEN_276 : _GEN_404; // @[decode.scala 344:35]
  wire  _GEN_469 = _T_21 ? _GEN_277 : _GEN_405; // @[decode.scala 344:35]
  wire  _GEN_470 = _T_21 ? _GEN_278 : _GEN_406; // @[decode.scala 344:35]
  wire  _GEN_471 = _T_21 ? _GEN_279 : _GEN_407; // @[decode.scala 344:35]
  wire  _GEN_472 = _T_21 ? _GEN_280 : _GEN_408; // @[decode.scala 344:35]
  wire  _GEN_473 = _T_21 ? _GEN_281 : _GEN_409; // @[decode.scala 344:35]
  wire  _GEN_474 = _T_21 ? _GEN_282 : _GEN_410; // @[decode.scala 344:35]
  wire  _GEN_475 = _T_21 ? _GEN_283 : _GEN_411; // @[decode.scala 344:35]
  wire  _GEN_476 = _T_21 ? _GEN_284 : _GEN_412; // @[decode.scala 344:35]
  wire  _GEN_477 = _T_21 ? _GEN_285 : _GEN_413; // @[decode.scala 344:35]
  wire  _GEN_478 = _T_21 ? _GEN_286 : _GEN_414; // @[decode.scala 344:35]
  wire  _GEN_479 = _T_21 ? _GEN_287 : _GEN_415; // @[decode.scala 344:35]
  wire  _GEN_480 = _T_21 ? _GEN_288 : _GEN_416; // @[decode.scala 344:35]
  wire  _GEN_481 = _T_21 ? _GEN_289 : _GEN_417; // @[decode.scala 344:35]
  wire  _GEN_482 = _T_21 ? _GEN_290 : _GEN_418; // @[decode.scala 344:35]
  wire  _GEN_483 = _T_21 ? _GEN_291 : _GEN_419; // @[decode.scala 344:35]
  wire  _GEN_484 = _T_21 ? _GEN_292 : _GEN_420; // @[decode.scala 344:35]
  wire  _GEN_485 = _T_21 ? _GEN_293 : _GEN_421; // @[decode.scala 344:35]
  wire  _GEN_486 = _T_21 ? _GEN_294 : _GEN_422; // @[decode.scala 344:35]
  wire  _GEN_487 = _T_21 ? _GEN_295 : _GEN_423; // @[decode.scala 344:35]
  wire  _GEN_488 = _T_21 ? _GEN_296 : _GEN_424; // @[decode.scala 344:35]
  wire  _GEN_489 = _T_21 ? _GEN_297 : _GEN_425; // @[decode.scala 344:35]
  wire  _GEN_490 = _T_21 ? _GEN_298 : _GEN_426; // @[decode.scala 344:35]
  wire  _GEN_491 = _T_21 ? _GEN_299 : _GEN_427; // @[decode.scala 344:35]
  wire  _GEN_492 = _T_21 ? _GEN_300 : _GEN_428; // @[decode.scala 344:35]
  wire  _GEN_493 = _T_21 ? _GEN_301 : _GEN_429; // @[decode.scala 344:35]
  wire  _GEN_494 = _T_21 ? _GEN_302 : _GEN_430; // @[decode.scala 344:35]
  wire  _GEN_495 = _T_21 ? _GEN_303 : _GEN_431; // @[decode.scala 344:35]
  wire  _GEN_496 = _T_21 ? _GEN_304 : _GEN_432; // @[decode.scala 344:35]
  wire  _GEN_497 = _T_21 ? _GEN_305 : _GEN_433; // @[decode.scala 344:35]
  wire  _GEN_498 = _T_21 ? _GEN_306 : _GEN_434; // @[decode.scala 344:35]
  wire  _GEN_499 = _T_21 ? _GEN_307 : _GEN_435; // @[decode.scala 344:35]
  wire  _GEN_500 = _T_21 ? _GEN_308 : _GEN_436; // @[decode.scala 344:35]
  wire  _GEN_501 = _T_21 ? _GEN_309 : _GEN_437; // @[decode.scala 344:35]
  wire  _GEN_502 = _T_21 ? _GEN_310 : _GEN_438; // @[decode.scala 344:35]
  wire  _GEN_503 = _T_21 ? _GEN_311 : _GEN_439; // @[decode.scala 344:35]
  wire  _GEN_504 = _T_21 ? _GEN_312 : _GEN_440; // @[decode.scala 344:35]
  wire  _GEN_505 = _T_21 ? _GEN_313 : _GEN_441; // @[decode.scala 344:35]
  wire  _GEN_506 = _T_21 ? _GEN_314 : _GEN_442; // @[decode.scala 344:35]
  wire  _GEN_507 = _T_21 ? _GEN_315 : _GEN_443; // @[decode.scala 344:35]
  wire  _GEN_508 = _T_21 ? _GEN_316 : _GEN_444; // @[decode.scala 344:35]
  wire  _GEN_509 = _T_21 ? _GEN_317 : _GEN_445; // @[decode.scala 344:35]
  wire  _GEN_510 = _T_21 ? _GEN_318 : _GEN_446; // @[decode.scala 344:35]
  wire  _GEN_511 = _T_21 ? _GEN_319 : _GEN_447; // @[decode.scala 344:35]
  wire  _GEN_512 = _T_21 ? _GEN_320 : _GEN_448; // @[decode.scala 344:35]
  wire  _GEN_513 = _T_21 ? _GEN_321 : _GEN_449; // @[decode.scala 344:35]
  wire  _GEN_514 = _T_21 ? _GEN_322 : _GEN_450; // @[decode.scala 344:35]
  wire  _GEN_515 = _T_21 ? _GEN_323 : _GEN_451; // @[decode.scala 344:35]
  wire  _GEN_516 = _T_21 ? _GEN_324 : _GEN_452; // @[decode.scala 344:35]
  wire  _GEN_517 = _T_21 ? _GEN_325 : _GEN_453; // @[decode.scala 344:35]
  wire  _GEN_518 = _T_21 ? _GEN_326 : _GEN_454; // @[decode.scala 344:35]
  wire  _GEN_519 = _T_21 ? _GEN_327 : _GEN_455; // @[decode.scala 344:35]
  wire  _GEN_520 = _T_21 ? _GEN_328 : _GEN_456; // @[decode.scala 344:35]
  wire  _GEN_521 = _T_21 ? _GEN_329 : _GEN_457; // @[decode.scala 344:35]
  wire  _GEN_522 = _T_21 ? _GEN_330 : _GEN_458; // @[decode.scala 344:35]
  wire  _GEN_523 = _T_21 ? _GEN_331 : _GEN_459; // @[decode.scala 344:35]
  wire  _GEN_524 = _T_21 ? _GEN_332 : _GEN_460; // @[decode.scala 344:35]
  wire  _GEN_525 = _T_21 ? _GEN_333 : _GEN_461; // @[decode.scala 344:35]
  wire  _GEN_526 = _T_21 ? _GEN_334 : _GEN_462; // @[decode.scala 344:35]
  wire  _GEN_527 = _T_21 ? _GEN_335 : _GEN_463; // @[decode.scala 344:35]
  wire  _GEN_530 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_465 : PRFFreeList_0; // @[decode.scala 310:36 342:60]
  wire  _GEN_531 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_466 : PRFFreeList_1; // @[decode.scala 310:36 342:60]
  wire  _GEN_532 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_467 : PRFFreeList_2; // @[decode.scala 310:36 342:60]
  wire  _GEN_533 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_468 : PRFFreeList_3; // @[decode.scala 310:36 342:60]
  wire  _GEN_534 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_469 : PRFFreeList_4; // @[decode.scala 310:36 342:60]
  wire  _GEN_535 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_470 : PRFFreeList_5; // @[decode.scala 310:36 342:60]
  wire  _GEN_536 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_471 : PRFFreeList_6; // @[decode.scala 310:36 342:60]
  wire  _GEN_537 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_472 : PRFFreeList_7; // @[decode.scala 310:36 342:60]
  wire  _GEN_538 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_473 : PRFFreeList_8; // @[decode.scala 310:36 342:60]
  wire  _GEN_539 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_474 : PRFFreeList_9; // @[decode.scala 310:36 342:60]
  wire  _GEN_540 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_475 : PRFFreeList_10; // @[decode.scala 310:36 342:60]
  wire  _GEN_541 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_476 : PRFFreeList_11; // @[decode.scala 310:36 342:60]
  wire  _GEN_542 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_477 : PRFFreeList_12; // @[decode.scala 310:36 342:60]
  wire  _GEN_543 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_478 : PRFFreeList_13; // @[decode.scala 310:36 342:60]
  wire  _GEN_544 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_479 : PRFFreeList_14; // @[decode.scala 310:36 342:60]
  wire  _GEN_545 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_480 : PRFFreeList_15; // @[decode.scala 310:36 342:60]
  wire  _GEN_546 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_481 : PRFFreeList_16; // @[decode.scala 310:36 342:60]
  wire  _GEN_547 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_482 : PRFFreeList_17; // @[decode.scala 310:36 342:60]
  wire  _GEN_548 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_483 : PRFFreeList_18; // @[decode.scala 310:36 342:60]
  wire  _GEN_549 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_484 : PRFFreeList_19; // @[decode.scala 310:36 342:60]
  wire  _GEN_550 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_485 : PRFFreeList_20; // @[decode.scala 310:36 342:60]
  wire  _GEN_551 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_486 : PRFFreeList_21; // @[decode.scala 310:36 342:60]
  wire  _GEN_552 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_487 : PRFFreeList_22; // @[decode.scala 310:36 342:60]
  wire  _GEN_553 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_488 : PRFFreeList_23; // @[decode.scala 310:36 342:60]
  wire  _GEN_554 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_489 : PRFFreeList_24; // @[decode.scala 310:36 342:60]
  wire  _GEN_555 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_490 : PRFFreeList_25; // @[decode.scala 310:36 342:60]
  wire  _GEN_556 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_491 : PRFFreeList_26; // @[decode.scala 310:36 342:60]
  wire  _GEN_557 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_492 : PRFFreeList_27; // @[decode.scala 310:36 342:60]
  wire  _GEN_558 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_493 : PRFFreeList_28; // @[decode.scala 310:36 342:60]
  wire  _GEN_559 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_494 : PRFFreeList_29; // @[decode.scala 310:36 342:60]
  wire  _GEN_560 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_495 : PRFFreeList_30; // @[decode.scala 310:36 342:60]
  wire  _GEN_561 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_496 : PRFFreeList_31; // @[decode.scala 310:36 342:60]
  wire  _GEN_562 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_497 : PRFFreeList_32; // @[decode.scala 310:36 342:60]
  wire  _GEN_563 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_498 : PRFFreeList_33; // @[decode.scala 310:36 342:60]
  wire  _GEN_564 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_499 : PRFFreeList_34; // @[decode.scala 310:36 342:60]
  wire  _GEN_565 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_500 : PRFFreeList_35; // @[decode.scala 310:36 342:60]
  wire  _GEN_566 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_501 : PRFFreeList_36; // @[decode.scala 310:36 342:60]
  wire  _GEN_567 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_502 : PRFFreeList_37; // @[decode.scala 310:36 342:60]
  wire  _GEN_568 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_503 : PRFFreeList_38; // @[decode.scala 310:36 342:60]
  wire  _GEN_569 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_504 : PRFFreeList_39; // @[decode.scala 310:36 342:60]
  wire  _GEN_570 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_505 : PRFFreeList_40; // @[decode.scala 310:36 342:60]
  wire  _GEN_571 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_506 : PRFFreeList_41; // @[decode.scala 310:36 342:60]
  wire  _GEN_572 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_507 : PRFFreeList_42; // @[decode.scala 310:36 342:60]
  wire  _GEN_573 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_508 : PRFFreeList_43; // @[decode.scala 310:36 342:60]
  wire  _GEN_574 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_509 : PRFFreeList_44; // @[decode.scala 310:36 342:60]
  wire  _GEN_575 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_510 : PRFFreeList_45; // @[decode.scala 310:36 342:60]
  wire  _GEN_576 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_511 : PRFFreeList_46; // @[decode.scala 310:36 342:60]
  wire  _GEN_577 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_512 : PRFFreeList_47; // @[decode.scala 310:36 342:60]
  wire  _GEN_578 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_513 : PRFFreeList_48; // @[decode.scala 310:36 342:60]
  wire  _GEN_579 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_514 : PRFFreeList_49; // @[decode.scala 310:36 342:60]
  wire  _GEN_580 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_515 : PRFFreeList_50; // @[decode.scala 310:36 342:60]
  wire  _GEN_581 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_516 : PRFFreeList_51; // @[decode.scala 310:36 342:60]
  wire  _GEN_582 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_517 : PRFFreeList_52; // @[decode.scala 310:36 342:60]
  wire  _GEN_583 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_518 : PRFFreeList_53; // @[decode.scala 310:36 342:60]
  wire  _GEN_584 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_519 : PRFFreeList_54; // @[decode.scala 310:36 342:60]
  wire  _GEN_585 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_520 : PRFFreeList_55; // @[decode.scala 310:36 342:60]
  wire  _GEN_586 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_521 : PRFFreeList_56; // @[decode.scala 310:36 342:60]
  wire  _GEN_587 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_522 : PRFFreeList_57; // @[decode.scala 310:36 342:60]
  wire  _GEN_588 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_523 : PRFFreeList_58; // @[decode.scala 310:36 342:60]
  wire  _GEN_589 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_524 : PRFFreeList_59; // @[decode.scala 310:36 342:60]
  wire  _GEN_590 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_525 : PRFFreeList_60; // @[decode.scala 310:36 342:60]
  wire  _GEN_591 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_526 : PRFFreeList_61; // @[decode.scala 310:36 342:60]
  wire  _GEN_592 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_527 : PRFFreeList_62; // @[decode.scala 310:36 342:60]
  wire  _GEN_658 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h0 == outputBuffer_PRFDest |
    PRFValidList_0 : PRFValidList_0; // @[decode.scala 199:29 351:71]
  wire  _GEN_659 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h1 == outputBuffer_PRFDest |
    PRFValidList_1 : PRFValidList_1; // @[decode.scala 199:29 351:71]
  wire  _GEN_660 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h2 == outputBuffer_PRFDest |
    PRFValidList_2 : PRFValidList_2; // @[decode.scala 199:29 351:71]
  wire  _GEN_661 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h3 == outputBuffer_PRFDest |
    PRFValidList_3 : PRFValidList_3; // @[decode.scala 199:29 351:71]
  wire  _GEN_662 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h4 == outputBuffer_PRFDest |
    PRFValidList_4 : PRFValidList_4; // @[decode.scala 199:29 351:71]
  wire  _GEN_663 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h5 == outputBuffer_PRFDest |
    PRFValidList_5 : PRFValidList_5; // @[decode.scala 199:29 351:71]
  wire  _GEN_664 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h6 == outputBuffer_PRFDest |
    PRFValidList_6 : PRFValidList_6; // @[decode.scala 199:29 351:71]
  wire  _GEN_665 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h7 == outputBuffer_PRFDest |
    PRFValidList_7 : PRFValidList_7; // @[decode.scala 199:29 351:71]
  wire  _GEN_666 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h8 == outputBuffer_PRFDest |
    PRFValidList_8 : PRFValidList_8; // @[decode.scala 199:29 351:71]
  wire  _GEN_667 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h9 == outputBuffer_PRFDest |
    PRFValidList_9 : PRFValidList_9; // @[decode.scala 199:29 351:71]
  wire  _GEN_668 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'ha == outputBuffer_PRFDest |
    PRFValidList_10 : PRFValidList_10; // @[decode.scala 199:29 351:71]
  wire  _GEN_669 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'hb == outputBuffer_PRFDest |
    PRFValidList_11 : PRFValidList_11; // @[decode.scala 199:29 351:71]
  wire  _GEN_670 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'hc == outputBuffer_PRFDest |
    PRFValidList_12 : PRFValidList_12; // @[decode.scala 199:29 351:71]
  wire  _GEN_671 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'hd == outputBuffer_PRFDest |
    PRFValidList_13 : PRFValidList_13; // @[decode.scala 199:29 351:71]
  wire  _GEN_672 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'he == outputBuffer_PRFDest |
    PRFValidList_14 : PRFValidList_14; // @[decode.scala 199:29 351:71]
  wire  _GEN_673 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'hf == outputBuffer_PRFDest |
    PRFValidList_15 : PRFValidList_15; // @[decode.scala 199:29 351:71]
  wire  _GEN_674 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h10 == outputBuffer_PRFDest |
    PRFValidList_16 : PRFValidList_16; // @[decode.scala 199:29 351:71]
  wire  _GEN_675 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h11 == outputBuffer_PRFDest |
    PRFValidList_17 : PRFValidList_17; // @[decode.scala 199:29 351:71]
  wire  _GEN_676 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h12 == outputBuffer_PRFDest |
    PRFValidList_18 : PRFValidList_18; // @[decode.scala 199:29 351:71]
  wire  _GEN_677 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h13 == outputBuffer_PRFDest |
    PRFValidList_19 : PRFValidList_19; // @[decode.scala 199:29 351:71]
  wire  _GEN_678 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h14 == outputBuffer_PRFDest |
    PRFValidList_20 : PRFValidList_20; // @[decode.scala 199:29 351:71]
  wire  _GEN_679 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h15 == outputBuffer_PRFDest |
    PRFValidList_21 : PRFValidList_21; // @[decode.scala 199:29 351:71]
  wire  _GEN_680 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h16 == outputBuffer_PRFDest |
    PRFValidList_22 : PRFValidList_22; // @[decode.scala 199:29 351:71]
  wire  _GEN_681 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h17 == outputBuffer_PRFDest |
    PRFValidList_23 : PRFValidList_23; // @[decode.scala 199:29 351:71]
  wire  _GEN_682 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h18 == outputBuffer_PRFDest |
    PRFValidList_24 : PRFValidList_24; // @[decode.scala 199:29 351:71]
  wire  _GEN_683 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h19 == outputBuffer_PRFDest |
    PRFValidList_25 : PRFValidList_25; // @[decode.scala 199:29 351:71]
  wire  _GEN_684 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h1a == outputBuffer_PRFDest |
    PRFValidList_26 : PRFValidList_26; // @[decode.scala 199:29 351:71]
  wire  _GEN_685 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h1b == outputBuffer_PRFDest |
    PRFValidList_27 : PRFValidList_27; // @[decode.scala 199:29 351:71]
  wire  _GEN_686 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h1c == outputBuffer_PRFDest |
    PRFValidList_28 : PRFValidList_28; // @[decode.scala 199:29 351:71]
  wire  _GEN_687 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h1d == outputBuffer_PRFDest |
    PRFValidList_29 : PRFValidList_29; // @[decode.scala 199:29 351:71]
  wire  _GEN_688 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h1e == outputBuffer_PRFDest |
    PRFValidList_30 : PRFValidList_30; // @[decode.scala 199:29 351:71]
  wire  _GEN_689 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h1f == outputBuffer_PRFDest |
    PRFValidList_31 : PRFValidList_31; // @[decode.scala 199:29 351:71]
  wire  _GEN_690 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h20 == outputBuffer_PRFDest |
    PRFValidList_32 : PRFValidList_32; // @[decode.scala 199:29 351:71]
  wire  _GEN_691 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h21 == outputBuffer_PRFDest |
    PRFValidList_33 : PRFValidList_33; // @[decode.scala 199:29 351:71]
  wire  _GEN_692 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h22 == outputBuffer_PRFDest |
    PRFValidList_34 : PRFValidList_34; // @[decode.scala 199:29 351:71]
  wire  _GEN_693 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h23 == outputBuffer_PRFDest |
    PRFValidList_35 : PRFValidList_35; // @[decode.scala 199:29 351:71]
  wire  _GEN_694 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h24 == outputBuffer_PRFDest |
    PRFValidList_36 : PRFValidList_36; // @[decode.scala 199:29 351:71]
  wire  _GEN_695 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h25 == outputBuffer_PRFDest |
    PRFValidList_37 : PRFValidList_37; // @[decode.scala 199:29 351:71]
  wire  _GEN_696 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h26 == outputBuffer_PRFDest |
    PRFValidList_38 : PRFValidList_38; // @[decode.scala 199:29 351:71]
  wire  _GEN_697 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h27 == outputBuffer_PRFDest |
    PRFValidList_39 : PRFValidList_39; // @[decode.scala 199:29 351:71]
  wire  _GEN_698 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h28 == outputBuffer_PRFDest |
    PRFValidList_40 : PRFValidList_40; // @[decode.scala 199:29 351:71]
  wire  _GEN_699 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h29 == outputBuffer_PRFDest |
    PRFValidList_41 : PRFValidList_41; // @[decode.scala 199:29 351:71]
  wire  _GEN_700 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h2a == outputBuffer_PRFDest |
    PRFValidList_42 : PRFValidList_42; // @[decode.scala 199:29 351:71]
  wire  _GEN_701 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h2b == outputBuffer_PRFDest |
    PRFValidList_43 : PRFValidList_43; // @[decode.scala 199:29 351:71]
  wire  _GEN_702 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h2c == outputBuffer_PRFDest |
    PRFValidList_44 : PRFValidList_44; // @[decode.scala 199:29 351:71]
  wire  _GEN_703 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h2d == outputBuffer_PRFDest |
    PRFValidList_45 : PRFValidList_45; // @[decode.scala 199:29 351:71]
  wire  _GEN_704 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h2e == outputBuffer_PRFDest |
    PRFValidList_46 : PRFValidList_46; // @[decode.scala 199:29 351:71]
  wire  _GEN_705 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h2f == outputBuffer_PRFDest |
    PRFValidList_47 : PRFValidList_47; // @[decode.scala 199:29 351:71]
  wire  _GEN_706 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h30 == outputBuffer_PRFDest |
    PRFValidList_48 : PRFValidList_48; // @[decode.scala 199:29 351:71]
  wire  _GEN_707 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h31 == outputBuffer_PRFDest |
    PRFValidList_49 : PRFValidList_49; // @[decode.scala 199:29 351:71]
  wire  _GEN_708 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h32 == outputBuffer_PRFDest |
    PRFValidList_50 : PRFValidList_50; // @[decode.scala 199:29 351:71]
  wire  _GEN_709 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h33 == outputBuffer_PRFDest |
    PRFValidList_51 : PRFValidList_51; // @[decode.scala 199:29 351:71]
  wire  _GEN_710 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h34 == outputBuffer_PRFDest |
    PRFValidList_52 : PRFValidList_52; // @[decode.scala 199:29 351:71]
  wire  _GEN_711 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h35 == outputBuffer_PRFDest |
    PRFValidList_53 : PRFValidList_53; // @[decode.scala 199:29 351:71]
  wire  _GEN_712 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h36 == outputBuffer_PRFDest |
    PRFValidList_54 : PRFValidList_54; // @[decode.scala 199:29 351:71]
  wire  _GEN_713 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h37 == outputBuffer_PRFDest |
    PRFValidList_55 : PRFValidList_55; // @[decode.scala 199:29 351:71]
  wire  _GEN_714 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h38 == outputBuffer_PRFDest |
    PRFValidList_56 : PRFValidList_56; // @[decode.scala 199:29 351:71]
  wire  _GEN_715 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h39 == outputBuffer_PRFDest |
    PRFValidList_57 : PRFValidList_57; // @[decode.scala 199:29 351:71]
  wire  _GEN_716 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h3a == outputBuffer_PRFDest |
    PRFValidList_58 : PRFValidList_58; // @[decode.scala 199:29 351:71]
  wire  _GEN_717 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h3b == outputBuffer_PRFDest |
    PRFValidList_59 : PRFValidList_59; // @[decode.scala 199:29 351:71]
  wire  _GEN_718 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h3c == outputBuffer_PRFDest |
    PRFValidList_60 : PRFValidList_60; // @[decode.scala 199:29 351:71]
  wire  _GEN_719 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h3d == outputBuffer_PRFDest |
    PRFValidList_61 : PRFValidList_61; // @[decode.scala 199:29 351:71]
  wire  _GEN_720 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h3e == outputBuffer_PRFDest |
    PRFValidList_62 : PRFValidList_62; // @[decode.scala 199:29 351:71]
  wire  _GEN_721 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h3f == outputBuffer_PRFDest |
    PRFValidList_63 : PRFValidList_63; // @[decode.scala 199:29 351:71]
  wire  _GEN_722 = 6'h0 == freeRegAddr ? 1'h0 : _GEN_530; // @[decode.scala 355:{33,33}]
  wire  _GEN_723 = 6'h1 == freeRegAddr ? 1'h0 : _GEN_531; // @[decode.scala 355:{33,33}]
  wire  _GEN_724 = 6'h2 == freeRegAddr ? 1'h0 : _GEN_532; // @[decode.scala 355:{33,33}]
  wire  _GEN_725 = 6'h3 == freeRegAddr ? 1'h0 : _GEN_533; // @[decode.scala 355:{33,33}]
  wire  _GEN_726 = 6'h4 == freeRegAddr ? 1'h0 : _GEN_534; // @[decode.scala 355:{33,33}]
  wire  _GEN_727 = 6'h5 == freeRegAddr ? 1'h0 : _GEN_535; // @[decode.scala 355:{33,33}]
  wire  _GEN_728 = 6'h6 == freeRegAddr ? 1'h0 : _GEN_536; // @[decode.scala 355:{33,33}]
  wire  _GEN_729 = 6'h7 == freeRegAddr ? 1'h0 : _GEN_537; // @[decode.scala 355:{33,33}]
  wire  _GEN_730 = 6'h8 == freeRegAddr ? 1'h0 : _GEN_538; // @[decode.scala 355:{33,33}]
  wire  _GEN_731 = 6'h9 == freeRegAddr ? 1'h0 : _GEN_539; // @[decode.scala 355:{33,33}]
  wire  _GEN_732 = 6'ha == freeRegAddr ? 1'h0 : _GEN_540; // @[decode.scala 355:{33,33}]
  wire  _GEN_733 = 6'hb == freeRegAddr ? 1'h0 : _GEN_541; // @[decode.scala 355:{33,33}]
  wire  _GEN_734 = 6'hc == freeRegAddr ? 1'h0 : _GEN_542; // @[decode.scala 355:{33,33}]
  wire  _GEN_735 = 6'hd == freeRegAddr ? 1'h0 : _GEN_543; // @[decode.scala 355:{33,33}]
  wire  _GEN_736 = 6'he == freeRegAddr ? 1'h0 : _GEN_544; // @[decode.scala 355:{33,33}]
  wire  _GEN_737 = 6'hf == freeRegAddr ? 1'h0 : _GEN_545; // @[decode.scala 355:{33,33}]
  wire  _GEN_738 = 6'h10 == freeRegAddr ? 1'h0 : _GEN_546; // @[decode.scala 355:{33,33}]
  wire  _GEN_739 = 6'h11 == freeRegAddr ? 1'h0 : _GEN_547; // @[decode.scala 355:{33,33}]
  wire  _GEN_740 = 6'h12 == freeRegAddr ? 1'h0 : _GEN_548; // @[decode.scala 355:{33,33}]
  wire  _GEN_741 = 6'h13 == freeRegAddr ? 1'h0 : _GEN_549; // @[decode.scala 355:{33,33}]
  wire  _GEN_742 = 6'h14 == freeRegAddr ? 1'h0 : _GEN_550; // @[decode.scala 355:{33,33}]
  wire  _GEN_743 = 6'h15 == freeRegAddr ? 1'h0 : _GEN_551; // @[decode.scala 355:{33,33}]
  wire  _GEN_744 = 6'h16 == freeRegAddr ? 1'h0 : _GEN_552; // @[decode.scala 355:{33,33}]
  wire  _GEN_745 = 6'h17 == freeRegAddr ? 1'h0 : _GEN_553; // @[decode.scala 355:{33,33}]
  wire  _GEN_746 = 6'h18 == freeRegAddr ? 1'h0 : _GEN_554; // @[decode.scala 355:{33,33}]
  wire  _GEN_747 = 6'h19 == freeRegAddr ? 1'h0 : _GEN_555; // @[decode.scala 355:{33,33}]
  wire  _GEN_748 = 6'h1a == freeRegAddr ? 1'h0 : _GEN_556; // @[decode.scala 355:{33,33}]
  wire  _GEN_749 = 6'h1b == freeRegAddr ? 1'h0 : _GEN_557; // @[decode.scala 355:{33,33}]
  wire  _GEN_750 = 6'h1c == freeRegAddr ? 1'h0 : _GEN_558; // @[decode.scala 355:{33,33}]
  wire  _GEN_751 = 6'h1d == freeRegAddr ? 1'h0 : _GEN_559; // @[decode.scala 355:{33,33}]
  wire  _GEN_752 = 6'h1e == freeRegAddr ? 1'h0 : _GEN_560; // @[decode.scala 355:{33,33}]
  wire  _GEN_753 = 6'h1f == freeRegAddr ? 1'h0 : _GEN_561; // @[decode.scala 355:{33,33}]
  wire  _GEN_754 = 6'h20 == freeRegAddr ? 1'h0 : _GEN_562; // @[decode.scala 355:{33,33}]
  wire  _GEN_755 = 6'h21 == freeRegAddr ? 1'h0 : _GEN_563; // @[decode.scala 355:{33,33}]
  wire  _GEN_756 = 6'h22 == freeRegAddr ? 1'h0 : _GEN_564; // @[decode.scala 355:{33,33}]
  wire  _GEN_757 = 6'h23 == freeRegAddr ? 1'h0 : _GEN_565; // @[decode.scala 355:{33,33}]
  wire  _GEN_758 = 6'h24 == freeRegAddr ? 1'h0 : _GEN_566; // @[decode.scala 355:{33,33}]
  wire  _GEN_759 = 6'h25 == freeRegAddr ? 1'h0 : _GEN_567; // @[decode.scala 355:{33,33}]
  wire  _GEN_760 = 6'h26 == freeRegAddr ? 1'h0 : _GEN_568; // @[decode.scala 355:{33,33}]
  wire  _GEN_761 = 6'h27 == freeRegAddr ? 1'h0 : _GEN_569; // @[decode.scala 355:{33,33}]
  wire  _GEN_762 = 6'h28 == freeRegAddr ? 1'h0 : _GEN_570; // @[decode.scala 355:{33,33}]
  wire  _GEN_763 = 6'h29 == freeRegAddr ? 1'h0 : _GEN_571; // @[decode.scala 355:{33,33}]
  wire  _GEN_764 = 6'h2a == freeRegAddr ? 1'h0 : _GEN_572; // @[decode.scala 355:{33,33}]
  wire  _GEN_765 = 6'h2b == freeRegAddr ? 1'h0 : _GEN_573; // @[decode.scala 355:{33,33}]
  wire  _GEN_766 = 6'h2c == freeRegAddr ? 1'h0 : _GEN_574; // @[decode.scala 355:{33,33}]
  wire  _GEN_767 = 6'h2d == freeRegAddr ? 1'h0 : _GEN_575; // @[decode.scala 355:{33,33}]
  wire  _GEN_768 = 6'h2e == freeRegAddr ? 1'h0 : _GEN_576; // @[decode.scala 355:{33,33}]
  wire  _GEN_769 = 6'h2f == freeRegAddr ? 1'h0 : _GEN_577; // @[decode.scala 355:{33,33}]
  wire  _GEN_770 = 6'h30 == freeRegAddr ? 1'h0 : _GEN_578; // @[decode.scala 355:{33,33}]
  wire  _GEN_771 = 6'h31 == freeRegAddr ? 1'h0 : _GEN_579; // @[decode.scala 355:{33,33}]
  wire  _GEN_772 = 6'h32 == freeRegAddr ? 1'h0 : _GEN_580; // @[decode.scala 355:{33,33}]
  wire  _GEN_773 = 6'h33 == freeRegAddr ? 1'h0 : _GEN_581; // @[decode.scala 355:{33,33}]
  wire  _GEN_774 = 6'h34 == freeRegAddr ? 1'h0 : _GEN_582; // @[decode.scala 355:{33,33}]
  wire  _GEN_775 = 6'h35 == freeRegAddr ? 1'h0 : _GEN_583; // @[decode.scala 355:{33,33}]
  wire  _GEN_776 = 6'h36 == freeRegAddr ? 1'h0 : _GEN_584; // @[decode.scala 355:{33,33}]
  wire  _GEN_777 = 6'h37 == freeRegAddr ? 1'h0 : _GEN_585; // @[decode.scala 355:{33,33}]
  wire  _GEN_778 = 6'h38 == freeRegAddr ? 1'h0 : _GEN_586; // @[decode.scala 355:{33,33}]
  wire  _GEN_779 = 6'h39 == freeRegAddr ? 1'h0 : _GEN_587; // @[decode.scala 355:{33,33}]
  wire  _GEN_780 = 6'h3a == freeRegAddr ? 1'h0 : _GEN_588; // @[decode.scala 355:{33,33}]
  wire  _GEN_781 = 6'h3b == freeRegAddr ? 1'h0 : _GEN_589; // @[decode.scala 355:{33,33}]
  wire  _GEN_782 = 6'h3c == freeRegAddr ? 1'h0 : _GEN_590; // @[decode.scala 355:{33,33}]
  wire  _GEN_783 = 6'h3d == freeRegAddr ? 1'h0 : _GEN_591; // @[decode.scala 355:{33,33}]
  wire  _GEN_784 = 6'h3e == freeRegAddr ? 1'h0 : _GEN_592; // @[decode.scala 355:{33,33}]
  wire  _GEN_786 = 6'h0 == freeRegAddr ? 1'h0 : _GEN_658; // @[decode.scala 356:{33,33}]
  wire  _GEN_787 = 6'h1 == freeRegAddr ? 1'h0 : _GEN_659; // @[decode.scala 356:{33,33}]
  wire  _GEN_788 = 6'h2 == freeRegAddr ? 1'h0 : _GEN_660; // @[decode.scala 356:{33,33}]
  wire  _GEN_789 = 6'h3 == freeRegAddr ? 1'h0 : _GEN_661; // @[decode.scala 356:{33,33}]
  wire  _GEN_790 = 6'h4 == freeRegAddr ? 1'h0 : _GEN_662; // @[decode.scala 356:{33,33}]
  wire  _GEN_791 = 6'h5 == freeRegAddr ? 1'h0 : _GEN_663; // @[decode.scala 356:{33,33}]
  wire  _GEN_792 = 6'h6 == freeRegAddr ? 1'h0 : _GEN_664; // @[decode.scala 356:{33,33}]
  wire  _GEN_793 = 6'h7 == freeRegAddr ? 1'h0 : _GEN_665; // @[decode.scala 356:{33,33}]
  wire  _GEN_794 = 6'h8 == freeRegAddr ? 1'h0 : _GEN_666; // @[decode.scala 356:{33,33}]
  wire  _GEN_795 = 6'h9 == freeRegAddr ? 1'h0 : _GEN_667; // @[decode.scala 356:{33,33}]
  wire  _GEN_796 = 6'ha == freeRegAddr ? 1'h0 : _GEN_668; // @[decode.scala 356:{33,33}]
  wire  _GEN_797 = 6'hb == freeRegAddr ? 1'h0 : _GEN_669; // @[decode.scala 356:{33,33}]
  wire  _GEN_798 = 6'hc == freeRegAddr ? 1'h0 : _GEN_670; // @[decode.scala 356:{33,33}]
  wire  _GEN_799 = 6'hd == freeRegAddr ? 1'h0 : _GEN_671; // @[decode.scala 356:{33,33}]
  wire  _GEN_800 = 6'he == freeRegAddr ? 1'h0 : _GEN_672; // @[decode.scala 356:{33,33}]
  wire  _GEN_801 = 6'hf == freeRegAddr ? 1'h0 : _GEN_673; // @[decode.scala 356:{33,33}]
  wire  _GEN_802 = 6'h10 == freeRegAddr ? 1'h0 : _GEN_674; // @[decode.scala 356:{33,33}]
  wire  _GEN_803 = 6'h11 == freeRegAddr ? 1'h0 : _GEN_675; // @[decode.scala 356:{33,33}]
  wire  _GEN_804 = 6'h12 == freeRegAddr ? 1'h0 : _GEN_676; // @[decode.scala 356:{33,33}]
  wire  _GEN_805 = 6'h13 == freeRegAddr ? 1'h0 : _GEN_677; // @[decode.scala 356:{33,33}]
  wire  _GEN_806 = 6'h14 == freeRegAddr ? 1'h0 : _GEN_678; // @[decode.scala 356:{33,33}]
  wire  _GEN_807 = 6'h15 == freeRegAddr ? 1'h0 : _GEN_679; // @[decode.scala 356:{33,33}]
  wire  _GEN_808 = 6'h16 == freeRegAddr ? 1'h0 : _GEN_680; // @[decode.scala 356:{33,33}]
  wire  _GEN_809 = 6'h17 == freeRegAddr ? 1'h0 : _GEN_681; // @[decode.scala 356:{33,33}]
  wire  _GEN_810 = 6'h18 == freeRegAddr ? 1'h0 : _GEN_682; // @[decode.scala 356:{33,33}]
  wire  _GEN_811 = 6'h19 == freeRegAddr ? 1'h0 : _GEN_683; // @[decode.scala 356:{33,33}]
  wire  _GEN_812 = 6'h1a == freeRegAddr ? 1'h0 : _GEN_684; // @[decode.scala 356:{33,33}]
  wire  _GEN_813 = 6'h1b == freeRegAddr ? 1'h0 : _GEN_685; // @[decode.scala 356:{33,33}]
  wire  _GEN_814 = 6'h1c == freeRegAddr ? 1'h0 : _GEN_686; // @[decode.scala 356:{33,33}]
  wire  _GEN_815 = 6'h1d == freeRegAddr ? 1'h0 : _GEN_687; // @[decode.scala 356:{33,33}]
  wire  _GEN_816 = 6'h1e == freeRegAddr ? 1'h0 : _GEN_688; // @[decode.scala 356:{33,33}]
  wire  _GEN_817 = 6'h1f == freeRegAddr ? 1'h0 : _GEN_689; // @[decode.scala 356:{33,33}]
  wire  _GEN_818 = 6'h20 == freeRegAddr ? 1'h0 : _GEN_690; // @[decode.scala 356:{33,33}]
  wire  _GEN_819 = 6'h21 == freeRegAddr ? 1'h0 : _GEN_691; // @[decode.scala 356:{33,33}]
  wire  _GEN_820 = 6'h22 == freeRegAddr ? 1'h0 : _GEN_692; // @[decode.scala 356:{33,33}]
  wire  _GEN_821 = 6'h23 == freeRegAddr ? 1'h0 : _GEN_693; // @[decode.scala 356:{33,33}]
  wire  _GEN_822 = 6'h24 == freeRegAddr ? 1'h0 : _GEN_694; // @[decode.scala 356:{33,33}]
  wire  _GEN_823 = 6'h25 == freeRegAddr ? 1'h0 : _GEN_695; // @[decode.scala 356:{33,33}]
  wire  _GEN_824 = 6'h26 == freeRegAddr ? 1'h0 : _GEN_696; // @[decode.scala 356:{33,33}]
  wire  _GEN_825 = 6'h27 == freeRegAddr ? 1'h0 : _GEN_697; // @[decode.scala 356:{33,33}]
  wire  _GEN_826 = 6'h28 == freeRegAddr ? 1'h0 : _GEN_698; // @[decode.scala 356:{33,33}]
  wire  _GEN_827 = 6'h29 == freeRegAddr ? 1'h0 : _GEN_699; // @[decode.scala 356:{33,33}]
  wire  _GEN_828 = 6'h2a == freeRegAddr ? 1'h0 : _GEN_700; // @[decode.scala 356:{33,33}]
  wire  _GEN_829 = 6'h2b == freeRegAddr ? 1'h0 : _GEN_701; // @[decode.scala 356:{33,33}]
  wire  _GEN_830 = 6'h2c == freeRegAddr ? 1'h0 : _GEN_702; // @[decode.scala 356:{33,33}]
  wire  _GEN_831 = 6'h2d == freeRegAddr ? 1'h0 : _GEN_703; // @[decode.scala 356:{33,33}]
  wire  _GEN_832 = 6'h2e == freeRegAddr ? 1'h0 : _GEN_704; // @[decode.scala 356:{33,33}]
  wire  _GEN_833 = 6'h2f == freeRegAddr ? 1'h0 : _GEN_705; // @[decode.scala 356:{33,33}]
  wire  _GEN_834 = 6'h30 == freeRegAddr ? 1'h0 : _GEN_706; // @[decode.scala 356:{33,33}]
  wire  _GEN_835 = 6'h31 == freeRegAddr ? 1'h0 : _GEN_707; // @[decode.scala 356:{33,33}]
  wire  _GEN_836 = 6'h32 == freeRegAddr ? 1'h0 : _GEN_708; // @[decode.scala 356:{33,33}]
  wire  _GEN_837 = 6'h33 == freeRegAddr ? 1'h0 : _GEN_709; // @[decode.scala 356:{33,33}]
  wire  _GEN_838 = 6'h34 == freeRegAddr ? 1'h0 : _GEN_710; // @[decode.scala 356:{33,33}]
  wire  _GEN_839 = 6'h35 == freeRegAddr ? 1'h0 : _GEN_711; // @[decode.scala 356:{33,33}]
  wire  _GEN_840 = 6'h36 == freeRegAddr ? 1'h0 : _GEN_712; // @[decode.scala 356:{33,33}]
  wire  _GEN_841 = 6'h37 == freeRegAddr ? 1'h0 : _GEN_713; // @[decode.scala 356:{33,33}]
  wire  _GEN_842 = 6'h38 == freeRegAddr ? 1'h0 : _GEN_714; // @[decode.scala 356:{33,33}]
  wire  _GEN_843 = 6'h39 == freeRegAddr ? 1'h0 : _GEN_715; // @[decode.scala 356:{33,33}]
  wire  _GEN_844 = 6'h3a == freeRegAddr ? 1'h0 : _GEN_716; // @[decode.scala 356:{33,33}]
  wire  _GEN_845 = 6'h3b == freeRegAddr ? 1'h0 : _GEN_717; // @[decode.scala 356:{33,33}]
  wire  _GEN_846 = 6'h3c == freeRegAddr ? 1'h0 : _GEN_718; // @[decode.scala 356:{33,33}]
  wire  _GEN_847 = 6'h3d == freeRegAddr ? 1'h0 : _GEN_719; // @[decode.scala 356:{33,33}]
  wire  _GEN_848 = 6'h3e == freeRegAddr ? 1'h0 : _GEN_720; // @[decode.scala 356:{33,33}]
  wire  _GEN_849 = 6'h3f == freeRegAddr ? 1'h0 : _GEN_721; // @[decode.scala 356:{33,33}]
  wire [5:0] _GEN_850 = 5'h0 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_0; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_851 = 5'h1 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_1; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_852 = 5'h2 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_2; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_853 = 5'h3 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_3; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_854 = 5'h4 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_4; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_855 = 5'h5 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_5; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_856 = 5'h6 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_6; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_857 = 5'h7 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_7; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_858 = 5'h8 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_8; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_859 = 5'h9 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_9; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_860 = 5'ha == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_10; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_861 = 5'hb == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_11; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_862 = 5'hc == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_12; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_863 = 5'hd == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_13; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_864 = 5'he == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_14; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_865 = 5'hf == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_15; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_866 = 5'h10 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_16; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_867 = 5'h11 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_17; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_868 = 5'h12 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_18; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_869 = 5'h13 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_19; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_870 = 5'h14 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_20; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_871 = 5'h15 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_21; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_872 = 5'h16 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_22; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_873 = 5'h17 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_23; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_874 = 5'h18 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_24; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_875 = 5'h19 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_25; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_876 = 5'h1a == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_26; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_877 = 5'h1b == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_27; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_878 = 5'h1c == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_28; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_879 = 5'h1d == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_29; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_880 = 5'h1e == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_30; // @[decode.scala 357:{33,33} 308:36]
  wire [5:0] _GEN_881 = 5'h1f == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_31; // @[decode.scala 357:{33,33} 308:36]
  wire  _GEN_882 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_722 : _GEN_530; // @[decode.scala 354:55]
  wire  _GEN_883 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_723 : _GEN_531; // @[decode.scala 354:55]
  wire  _GEN_884 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_724 : _GEN_532; // @[decode.scala 354:55]
  wire  _GEN_885 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_725 : _GEN_533; // @[decode.scala 354:55]
  wire  _GEN_886 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_726 : _GEN_534; // @[decode.scala 354:55]
  wire  _GEN_887 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_727 : _GEN_535; // @[decode.scala 354:55]
  wire  _GEN_888 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_728 : _GEN_536; // @[decode.scala 354:55]
  wire  _GEN_889 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_729 : _GEN_537; // @[decode.scala 354:55]
  wire  _GEN_890 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_730 : _GEN_538; // @[decode.scala 354:55]
  wire  _GEN_891 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_731 : _GEN_539; // @[decode.scala 354:55]
  wire  _GEN_892 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_732 : _GEN_540; // @[decode.scala 354:55]
  wire  _GEN_893 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_733 : _GEN_541; // @[decode.scala 354:55]
  wire  _GEN_894 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_734 : _GEN_542; // @[decode.scala 354:55]
  wire  _GEN_895 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_735 : _GEN_543; // @[decode.scala 354:55]
  wire  _GEN_896 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_736 : _GEN_544; // @[decode.scala 354:55]
  wire  _GEN_897 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_737 : _GEN_545; // @[decode.scala 354:55]
  wire  _GEN_898 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_738 : _GEN_546; // @[decode.scala 354:55]
  wire  _GEN_899 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_739 : _GEN_547; // @[decode.scala 354:55]
  wire  _GEN_900 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_740 : _GEN_548; // @[decode.scala 354:55]
  wire  _GEN_901 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_741 : _GEN_549; // @[decode.scala 354:55]
  wire  _GEN_902 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_742 : _GEN_550; // @[decode.scala 354:55]
  wire  _GEN_903 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_743 : _GEN_551; // @[decode.scala 354:55]
  wire  _GEN_904 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_744 : _GEN_552; // @[decode.scala 354:55]
  wire  _GEN_905 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_745 : _GEN_553; // @[decode.scala 354:55]
  wire  _GEN_906 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_746 : _GEN_554; // @[decode.scala 354:55]
  wire  _GEN_907 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_747 : _GEN_555; // @[decode.scala 354:55]
  wire  _GEN_908 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_748 : _GEN_556; // @[decode.scala 354:55]
  wire  _GEN_909 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_749 : _GEN_557; // @[decode.scala 354:55]
  wire  _GEN_910 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_750 : _GEN_558; // @[decode.scala 354:55]
  wire  _GEN_911 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_751 : _GEN_559; // @[decode.scala 354:55]
  wire  _GEN_912 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_752 : _GEN_560; // @[decode.scala 354:55]
  wire  _GEN_913 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_753 : _GEN_561; // @[decode.scala 354:55]
  wire  _GEN_914 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_754 : _GEN_562; // @[decode.scala 354:55]
  wire  _GEN_915 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_755 : _GEN_563; // @[decode.scala 354:55]
  wire  _GEN_916 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_756 : _GEN_564; // @[decode.scala 354:55]
  wire  _GEN_917 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_757 : _GEN_565; // @[decode.scala 354:55]
  wire  _GEN_918 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_758 : _GEN_566; // @[decode.scala 354:55]
  wire  _GEN_919 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_759 : _GEN_567; // @[decode.scala 354:55]
  wire  _GEN_920 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_760 : _GEN_568; // @[decode.scala 354:55]
  wire  _GEN_921 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_761 : _GEN_569; // @[decode.scala 354:55]
  wire  _GEN_922 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_762 : _GEN_570; // @[decode.scala 354:55]
  wire  _GEN_923 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_763 : _GEN_571; // @[decode.scala 354:55]
  wire  _GEN_924 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_764 : _GEN_572; // @[decode.scala 354:55]
  wire  _GEN_925 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_765 : _GEN_573; // @[decode.scala 354:55]
  wire  _GEN_926 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_766 : _GEN_574; // @[decode.scala 354:55]
  wire  _GEN_927 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_767 : _GEN_575; // @[decode.scala 354:55]
  wire  _GEN_928 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_768 : _GEN_576; // @[decode.scala 354:55]
  wire  _GEN_929 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_769 : _GEN_577; // @[decode.scala 354:55]
  wire  _GEN_930 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_770 : _GEN_578; // @[decode.scala 354:55]
  wire  _GEN_931 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_771 : _GEN_579; // @[decode.scala 354:55]
  wire  _GEN_932 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_772 : _GEN_580; // @[decode.scala 354:55]
  wire  _GEN_933 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_773 : _GEN_581; // @[decode.scala 354:55]
  wire  _GEN_934 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_774 : _GEN_582; // @[decode.scala 354:55]
  wire  _GEN_935 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_775 : _GEN_583; // @[decode.scala 354:55]
  wire  _GEN_936 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_776 : _GEN_584; // @[decode.scala 354:55]
  wire  _GEN_937 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_777 : _GEN_585; // @[decode.scala 354:55]
  wire  _GEN_938 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_778 : _GEN_586; // @[decode.scala 354:55]
  wire  _GEN_939 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_779 : _GEN_587; // @[decode.scala 354:55]
  wire  _GEN_940 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_780 : _GEN_588; // @[decode.scala 354:55]
  wire  _GEN_941 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_781 : _GEN_589; // @[decode.scala 354:55]
  wire  _GEN_942 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_782 : _GEN_590; // @[decode.scala 354:55]
  wire  _GEN_943 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_783 : _GEN_591; // @[decode.scala 354:55]
  wire  _GEN_944 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_784 : _GEN_592; // @[decode.scala 354:55]
  wire  _GEN_946 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_786 : _GEN_658; // @[decode.scala 354:55]
  wire  _GEN_947 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_787 : _GEN_659; // @[decode.scala 354:55]
  wire  _GEN_948 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_788 : _GEN_660; // @[decode.scala 354:55]
  wire  _GEN_949 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_789 : _GEN_661; // @[decode.scala 354:55]
  wire  _GEN_950 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_790 : _GEN_662; // @[decode.scala 354:55]
  wire  _GEN_951 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_791 : _GEN_663; // @[decode.scala 354:55]
  wire  _GEN_952 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_792 : _GEN_664; // @[decode.scala 354:55]
  wire  _GEN_953 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_793 : _GEN_665; // @[decode.scala 354:55]
  wire  _GEN_954 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_794 : _GEN_666; // @[decode.scala 354:55]
  wire  _GEN_955 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_795 : _GEN_667; // @[decode.scala 354:55]
  wire  _GEN_956 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_796 : _GEN_668; // @[decode.scala 354:55]
  wire  _GEN_957 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_797 : _GEN_669; // @[decode.scala 354:55]
  wire  _GEN_958 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_798 : _GEN_670; // @[decode.scala 354:55]
  wire  _GEN_959 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_799 : _GEN_671; // @[decode.scala 354:55]
  wire  _GEN_960 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_800 : _GEN_672; // @[decode.scala 354:55]
  wire  _GEN_961 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_801 : _GEN_673; // @[decode.scala 354:55]
  wire  _GEN_962 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_802 : _GEN_674; // @[decode.scala 354:55]
  wire  _GEN_963 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_803 : _GEN_675; // @[decode.scala 354:55]
  wire  _GEN_964 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_804 : _GEN_676; // @[decode.scala 354:55]
  wire  _GEN_965 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_805 : _GEN_677; // @[decode.scala 354:55]
  wire  _GEN_966 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_806 : _GEN_678; // @[decode.scala 354:55]
  wire  _GEN_967 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_807 : _GEN_679; // @[decode.scala 354:55]
  wire  _GEN_968 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_808 : _GEN_680; // @[decode.scala 354:55]
  wire  _GEN_969 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_809 : _GEN_681; // @[decode.scala 354:55]
  wire  _GEN_970 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_810 : _GEN_682; // @[decode.scala 354:55]
  wire  _GEN_971 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_811 : _GEN_683; // @[decode.scala 354:55]
  wire  _GEN_972 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_812 : _GEN_684; // @[decode.scala 354:55]
  wire  _GEN_973 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_813 : _GEN_685; // @[decode.scala 354:55]
  wire  _GEN_974 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_814 : _GEN_686; // @[decode.scala 354:55]
  wire  _GEN_975 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_815 : _GEN_687; // @[decode.scala 354:55]
  wire  _GEN_976 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_816 : _GEN_688; // @[decode.scala 354:55]
  wire  _GEN_977 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_817 : _GEN_689; // @[decode.scala 354:55]
  wire  _GEN_978 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_818 : _GEN_690; // @[decode.scala 354:55]
  wire  _GEN_979 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_819 : _GEN_691; // @[decode.scala 354:55]
  wire  _GEN_980 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_820 : _GEN_692; // @[decode.scala 354:55]
  wire  _GEN_981 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_821 : _GEN_693; // @[decode.scala 354:55]
  wire  _GEN_982 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_822 : _GEN_694; // @[decode.scala 354:55]
  wire  _GEN_983 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_823 : _GEN_695; // @[decode.scala 354:55]
  wire  _GEN_984 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_824 : _GEN_696; // @[decode.scala 354:55]
  wire  _GEN_985 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_825 : _GEN_697; // @[decode.scala 354:55]
  wire  _GEN_986 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_826 : _GEN_698; // @[decode.scala 354:55]
  wire  _GEN_987 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_827 : _GEN_699; // @[decode.scala 354:55]
  wire  _GEN_988 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_828 : _GEN_700; // @[decode.scala 354:55]
  wire  _GEN_989 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_829 : _GEN_701; // @[decode.scala 354:55]
  wire  _GEN_990 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_830 : _GEN_702; // @[decode.scala 354:55]
  wire  _GEN_991 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_831 : _GEN_703; // @[decode.scala 354:55]
  wire  _GEN_992 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_832 : _GEN_704; // @[decode.scala 354:55]
  wire  _GEN_993 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_833 : _GEN_705; // @[decode.scala 354:55]
  wire  _GEN_994 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_834 : _GEN_706; // @[decode.scala 354:55]
  wire  _GEN_995 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_835 : _GEN_707; // @[decode.scala 354:55]
  wire  _GEN_996 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_836 : _GEN_708; // @[decode.scala 354:55]
  wire  _GEN_997 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_837 : _GEN_709; // @[decode.scala 354:55]
  wire  _GEN_998 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_838 : _GEN_710; // @[decode.scala 354:55]
  wire  _GEN_999 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_839 : _GEN_711; // @[decode.scala 354:55]
  wire  _GEN_1000 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_840 : _GEN_712; // @[decode.scala 354:55]
  wire  _GEN_1001 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_841 : _GEN_713; // @[decode.scala 354:55]
  wire  _GEN_1002 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_842 : _GEN_714; // @[decode.scala 354:55]
  wire  _GEN_1003 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_843 : _GEN_715; // @[decode.scala 354:55]
  wire  _GEN_1004 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_844 : _GEN_716; // @[decode.scala 354:55]
  wire  _GEN_1005 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_845 : _GEN_717; // @[decode.scala 354:55]
  wire  _GEN_1006 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_846 : _GEN_718; // @[decode.scala 354:55]
  wire  _GEN_1007 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_847 : _GEN_719; // @[decode.scala 354:55]
  wire  _GEN_1008 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_848 : _GEN_720; // @[decode.scala 354:55]
  wire  _GEN_1009 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_849 : _GEN_721; // @[decode.scala 354:55]
  wire [5:0] _GEN_1010 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_850 : frontEndRegMap_0; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1011 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_851 : frontEndRegMap_1; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1012 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_852 : frontEndRegMap_2; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1013 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_853 : frontEndRegMap_3; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1014 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_854 : frontEndRegMap_4; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1015 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_855 : frontEndRegMap_5; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1016 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_856 : frontEndRegMap_6; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1017 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_857 : frontEndRegMap_7; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1018 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_858 : frontEndRegMap_8; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1019 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_859 : frontEndRegMap_9; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1020 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_860 : frontEndRegMap_10; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1021 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_861 : frontEndRegMap_11; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1022 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_862 : frontEndRegMap_12; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1023 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_863 : frontEndRegMap_13; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1024 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_864 : frontEndRegMap_14; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1025 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_865 : frontEndRegMap_15; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1026 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_866 : frontEndRegMap_16; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1027 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_867 : frontEndRegMap_17; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1028 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_868 : frontEndRegMap_18; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1029 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_869 : frontEndRegMap_19; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1030 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_870 : frontEndRegMap_20; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1031 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_871 : frontEndRegMap_21; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1032 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_872 : frontEndRegMap_22; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1033 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_873 : frontEndRegMap_23; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1034 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_874 : frontEndRegMap_24; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1035 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_875 : frontEndRegMap_25; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1036 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_876 : frontEndRegMap_26; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1037 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_877 : frontEndRegMap_27; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1038 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_878 : frontEndRegMap_28; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1039 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_879 : frontEndRegMap_29; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1040 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_880 : frontEndRegMap_30; // @[decode.scala 308:36 354:55]
  wire [5:0] _GEN_1041 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_881 : frontEndRegMap_31; // @[decode.scala 308:36 354:55]
  wire  _GEN_1042 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_882 : _GEN_530; // @[decode.scala 353:149]
  wire  _GEN_1043 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_883 : _GEN_531; // @[decode.scala 353:149]
  wire  _GEN_1044 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_884 : _GEN_532; // @[decode.scala 353:149]
  wire  _GEN_1045 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_885 : _GEN_533; // @[decode.scala 353:149]
  wire  _GEN_1046 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_886 : _GEN_534; // @[decode.scala 353:149]
  wire  _GEN_1047 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_887 : _GEN_535; // @[decode.scala 353:149]
  wire  _GEN_1048 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_888 : _GEN_536; // @[decode.scala 353:149]
  wire  _GEN_1049 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_889 : _GEN_537; // @[decode.scala 353:149]
  wire  _GEN_1050 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_890 : _GEN_538; // @[decode.scala 353:149]
  wire  _GEN_1051 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_891 : _GEN_539; // @[decode.scala 353:149]
  wire  _GEN_1052 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_892 : _GEN_540; // @[decode.scala 353:149]
  wire  _GEN_1053 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_893 : _GEN_541; // @[decode.scala 353:149]
  wire  _GEN_1054 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_894 : _GEN_542; // @[decode.scala 353:149]
  wire  _GEN_1055 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_895 : _GEN_543; // @[decode.scala 353:149]
  wire  _GEN_1056 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_896 : _GEN_544; // @[decode.scala 353:149]
  wire  _GEN_1057 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_897 : _GEN_545; // @[decode.scala 353:149]
  wire  _GEN_1058 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_898 : _GEN_546; // @[decode.scala 353:149]
  wire  _GEN_1059 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_899 : _GEN_547; // @[decode.scala 353:149]
  wire  _GEN_1060 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_900 : _GEN_548; // @[decode.scala 353:149]
  wire  _GEN_1061 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_901 : _GEN_549; // @[decode.scala 353:149]
  wire  _GEN_1062 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_902 : _GEN_550; // @[decode.scala 353:149]
  wire  _GEN_1063 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_903 : _GEN_551; // @[decode.scala 353:149]
  wire  _GEN_1064 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_904 : _GEN_552; // @[decode.scala 353:149]
  wire  _GEN_1065 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_905 : _GEN_553; // @[decode.scala 353:149]
  wire  _GEN_1066 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_906 : _GEN_554; // @[decode.scala 353:149]
  wire  _GEN_1067 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_907 : _GEN_555; // @[decode.scala 353:149]
  wire  _GEN_1068 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_908 : _GEN_556; // @[decode.scala 353:149]
  wire  _GEN_1069 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_909 : _GEN_557; // @[decode.scala 353:149]
  wire  _GEN_1070 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_910 : _GEN_558; // @[decode.scala 353:149]
  wire  _GEN_1071 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_911 : _GEN_559; // @[decode.scala 353:149]
  wire  _GEN_1072 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_912 : _GEN_560; // @[decode.scala 353:149]
  wire  _GEN_1073 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_913 : _GEN_561; // @[decode.scala 353:149]
  wire  _GEN_1074 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_914 : _GEN_562; // @[decode.scala 353:149]
  wire  _GEN_1075 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_915 : _GEN_563; // @[decode.scala 353:149]
  wire  _GEN_1076 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_916 : _GEN_564; // @[decode.scala 353:149]
  wire  _GEN_1077 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_917 : _GEN_565; // @[decode.scala 353:149]
  wire  _GEN_1078 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_918 : _GEN_566; // @[decode.scala 353:149]
  wire  _GEN_1079 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_919 : _GEN_567; // @[decode.scala 353:149]
  wire  _GEN_1080 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_920 : _GEN_568; // @[decode.scala 353:149]
  wire  _GEN_1081 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_921 : _GEN_569; // @[decode.scala 353:149]
  wire  _GEN_1082 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_922 : _GEN_570; // @[decode.scala 353:149]
  wire  _GEN_1083 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_923 : _GEN_571; // @[decode.scala 353:149]
  wire  _GEN_1084 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_924 : _GEN_572; // @[decode.scala 353:149]
  wire  _GEN_1085 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_925 : _GEN_573; // @[decode.scala 353:149]
  wire  _GEN_1086 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_926 : _GEN_574; // @[decode.scala 353:149]
  wire  _GEN_1087 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_927 : _GEN_575; // @[decode.scala 353:149]
  wire  _GEN_1088 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_928 : _GEN_576; // @[decode.scala 353:149]
  wire  _GEN_1089 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_929 : _GEN_577; // @[decode.scala 353:149]
  wire  _GEN_1090 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_930 : _GEN_578; // @[decode.scala 353:149]
  wire  _GEN_1091 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_931 : _GEN_579; // @[decode.scala 353:149]
  wire  _GEN_1092 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_932 : _GEN_580; // @[decode.scala 353:149]
  wire  _GEN_1093 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_933 : _GEN_581; // @[decode.scala 353:149]
  wire  _GEN_1094 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_934 : _GEN_582; // @[decode.scala 353:149]
  wire  _GEN_1095 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_935 : _GEN_583; // @[decode.scala 353:149]
  wire  _GEN_1096 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_936 : _GEN_584; // @[decode.scala 353:149]
  wire  _GEN_1097 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_937 : _GEN_585; // @[decode.scala 353:149]
  wire  _GEN_1098 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_938 : _GEN_586; // @[decode.scala 353:149]
  wire  _GEN_1099 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_939 : _GEN_587; // @[decode.scala 353:149]
  wire  _GEN_1100 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_940 : _GEN_588; // @[decode.scala 353:149]
  wire  _GEN_1101 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_941 : _GEN_589; // @[decode.scala 353:149]
  wire  _GEN_1102 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_942 : _GEN_590; // @[decode.scala 353:149]
  wire  _GEN_1103 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_943 : _GEN_591; // @[decode.scala 353:149]
  wire  _GEN_1104 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_944 : _GEN_592; // @[decode.scala 353:149]
  wire  _GEN_1106 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_946 : _GEN_658; // @[decode.scala 353:149]
  wire  _GEN_1107 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_947 : _GEN_659; // @[decode.scala 353:149]
  wire  _GEN_1108 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_948 : _GEN_660; // @[decode.scala 353:149]
  wire  _GEN_1109 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_949 : _GEN_661; // @[decode.scala 353:149]
  wire  _GEN_1110 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_950 : _GEN_662; // @[decode.scala 353:149]
  wire  _GEN_1111 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_951 : _GEN_663; // @[decode.scala 353:149]
  wire  _GEN_1112 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_952 : _GEN_664; // @[decode.scala 353:149]
  wire  _GEN_1113 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_953 : _GEN_665; // @[decode.scala 353:149]
  wire  _GEN_1114 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_954 : _GEN_666; // @[decode.scala 353:149]
  wire  _GEN_1115 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_955 : _GEN_667; // @[decode.scala 353:149]
  wire  _GEN_1116 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_956 : _GEN_668; // @[decode.scala 353:149]
  wire  _GEN_1117 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_957 : _GEN_669; // @[decode.scala 353:149]
  wire  _GEN_1118 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_958 : _GEN_670; // @[decode.scala 353:149]
  wire  _GEN_1119 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_959 : _GEN_671; // @[decode.scala 353:149]
  wire  _GEN_1120 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_960 : _GEN_672; // @[decode.scala 353:149]
  wire  _GEN_1121 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_961 : _GEN_673; // @[decode.scala 353:149]
  wire  _GEN_1122 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_962 : _GEN_674; // @[decode.scala 353:149]
  wire  _GEN_1123 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_963 : _GEN_675; // @[decode.scala 353:149]
  wire  _GEN_1124 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_964 : _GEN_676; // @[decode.scala 353:149]
  wire  _GEN_1125 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_965 : _GEN_677; // @[decode.scala 353:149]
  wire  _GEN_1126 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_966 : _GEN_678; // @[decode.scala 353:149]
  wire  _GEN_1127 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_967 : _GEN_679; // @[decode.scala 353:149]
  wire  _GEN_1128 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_968 : _GEN_680; // @[decode.scala 353:149]
  wire  _GEN_1129 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_969 : _GEN_681; // @[decode.scala 353:149]
  wire  _GEN_1130 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_970 : _GEN_682; // @[decode.scala 353:149]
  wire  _GEN_1131 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_971 : _GEN_683; // @[decode.scala 353:149]
  wire  _GEN_1132 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_972 : _GEN_684; // @[decode.scala 353:149]
  wire  _GEN_1133 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_973 : _GEN_685; // @[decode.scala 353:149]
  wire  _GEN_1134 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_974 : _GEN_686; // @[decode.scala 353:149]
  wire  _GEN_1135 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_975 : _GEN_687; // @[decode.scala 353:149]
  wire  _GEN_1136 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_976 : _GEN_688; // @[decode.scala 353:149]
  wire  _GEN_1137 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_977 : _GEN_689; // @[decode.scala 353:149]
  wire  _GEN_1138 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_978 : _GEN_690; // @[decode.scala 353:149]
  wire  _GEN_1139 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_979 : _GEN_691; // @[decode.scala 353:149]
  wire  _GEN_1140 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_980 : _GEN_692; // @[decode.scala 353:149]
  wire  _GEN_1141 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_981 : _GEN_693; // @[decode.scala 353:149]
  wire  _GEN_1142 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_982 : _GEN_694; // @[decode.scala 353:149]
  wire  _GEN_1143 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_983 : _GEN_695; // @[decode.scala 353:149]
  wire  _GEN_1144 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_984 : _GEN_696; // @[decode.scala 353:149]
  wire  _GEN_1145 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_985 : _GEN_697; // @[decode.scala 353:149]
  wire  _GEN_1146 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_986 : _GEN_698; // @[decode.scala 353:149]
  wire  _GEN_1147 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_987 : _GEN_699; // @[decode.scala 353:149]
  wire  _GEN_1148 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_988 : _GEN_700; // @[decode.scala 353:149]
  wire  _GEN_1149 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_989 : _GEN_701; // @[decode.scala 353:149]
  wire  _GEN_1150 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_990 : _GEN_702; // @[decode.scala 353:149]
  wire  _GEN_1151 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_991 : _GEN_703; // @[decode.scala 353:149]
  wire  _GEN_1152 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_992 : _GEN_704; // @[decode.scala 353:149]
  wire  _GEN_1153 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_993 : _GEN_705; // @[decode.scala 353:149]
  wire  _GEN_1154 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_994 : _GEN_706; // @[decode.scala 353:149]
  wire  _GEN_1155 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_995 : _GEN_707; // @[decode.scala 353:149]
  wire  _GEN_1156 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_996 : _GEN_708; // @[decode.scala 353:149]
  wire  _GEN_1157 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_997 : _GEN_709; // @[decode.scala 353:149]
  wire  _GEN_1158 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_998 : _GEN_710; // @[decode.scala 353:149]
  wire  _GEN_1159 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_999 : _GEN_711; // @[decode.scala 353:149]
  wire  _GEN_1160 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1000 : _GEN_712; // @[decode.scala 353:149]
  wire  _GEN_1161 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1001 : _GEN_713; // @[decode.scala 353:149]
  wire  _GEN_1162 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1002 : _GEN_714; // @[decode.scala 353:149]
  wire  _GEN_1163 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1003 : _GEN_715; // @[decode.scala 353:149]
  wire  _GEN_1164 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1004 : _GEN_716; // @[decode.scala 353:149]
  wire  _GEN_1165 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1005 : _GEN_717; // @[decode.scala 353:149]
  wire  _GEN_1166 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1006 : _GEN_718; // @[decode.scala 353:149]
  wire  _GEN_1167 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1007 : _GEN_719; // @[decode.scala 353:149]
  wire  _GEN_1168 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1008 : _GEN_720; // @[decode.scala 353:149]
  wire  _GEN_1169 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1009 : _GEN_721; // @[decode.scala 353:149]
  wire [5:0] _GEN_1170 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1010 : frontEndRegMap_0; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1171 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1011 : frontEndRegMap_1; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1172 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1012 : frontEndRegMap_2; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1173 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1013 : frontEndRegMap_3; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1174 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1014 : frontEndRegMap_4; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1175 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1015 : frontEndRegMap_5; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1176 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1016 : frontEndRegMap_6; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1177 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1017 : frontEndRegMap_7; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1178 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1018 : frontEndRegMap_8; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1179 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1019 : frontEndRegMap_9; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1180 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1020 : frontEndRegMap_10; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1181 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1021 : frontEndRegMap_11; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1182 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1022 : frontEndRegMap_12; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1183 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1023 : frontEndRegMap_13; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1184 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1024 : frontEndRegMap_14; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1185 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1025 : frontEndRegMap_15; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1186 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1026 : frontEndRegMap_16; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1187 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1027 : frontEndRegMap_17; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1188 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1028 : frontEndRegMap_18; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1189 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1029 : frontEndRegMap_19; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1190 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1030 : frontEndRegMap_20; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1191 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1031 : frontEndRegMap_21; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1192 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1032 : frontEndRegMap_22; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1193 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1033 : frontEndRegMap_23; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1194 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1034 : frontEndRegMap_24; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1195 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1035 : frontEndRegMap_25; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1196 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1036 : frontEndRegMap_26; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1197 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1037 : frontEndRegMap_27; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1198 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1038 : frontEndRegMap_28; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1199 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1039 : frontEndRegMap_29; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1200 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1040 : frontEndRegMap_30; // @[decode.scala 353:149 308:36]
  wire [5:0] _GEN_1201 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1041 : frontEndRegMap_31; // @[decode.scala 353:149 308:36]
  wire [2:0] _branchTracker_T_1 = branchTracker - 3'h1; // @[decode.scala 364:36]
  wire [4:0] _T_44 = _toExec_branchMask_T & 5'h10; // @[decode.scala 367:73]
  wire [4:0] _T_46 = ~branchEvalIn_branchMask; // @[decode.scala 367:124]
  wire [4:0] _T_47 = _toExec_branchMask_T & _T_46; // @[decode.scala 367:121]
  wire [4:0] _T_48 = _T_47 & 5'hf; // @[decode.scala 367:151]
  wire [4:0] _T_49 = _T_44 | _T_48; // @[decode.scala 367:86]
  wire  _GEN_1202 = 6'h0 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1203 = 6'h1 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1204 = 6'h2 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1205 = 6'h3 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1206 = 6'h4 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1207 = 6'h5 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1208 = 6'h6 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1209 = 6'h7 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1210 = 6'h8 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1211 = 6'h9 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1212 = 6'ha == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1213 = 6'hb == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1214 = 6'hc == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1215 = 6'hd == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1216 = 6'he == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1217 = 6'hf == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1218 = 6'h10 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1219 = 6'h11 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1220 = 6'h12 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1221 = 6'h13 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1222 = 6'h14 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1223 = 6'h15 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1224 = 6'h16 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1225 = 6'h17 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1226 = 6'h18 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1227 = 6'h19 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1228 = 6'h1a == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1229 = 6'h1b == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1230 = 6'h1c == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1231 = 6'h1d == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1232 = 6'h1e == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1233 = 6'h1f == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1234 = 6'h20 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1235 = 6'h21 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1236 = 6'h22 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1237 = 6'h23 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1238 = 6'h24 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1239 = 6'h25 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1240 = 6'h26 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1241 = 6'h27 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1242 = 6'h28 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1243 = 6'h29 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1244 = 6'h2a == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1245 = 6'h2b == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1246 = 6'h2c == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1247 = 6'h2d == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1248 = 6'h2e == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1249 = 6'h2f == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1250 = 6'h30 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1251 = 6'h31 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1252 = 6'h32 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1253 = 6'h33 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1254 = 6'h34 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1255 = 6'h35 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1256 = 6'h36 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1257 = 6'h37 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1258 = 6'h38 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1259 = 6'h39 == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1260 = 6'h3a == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1261 = 6'h3b == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1262 = 6'h3c == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1263 = 6'h3d == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1264 = 6'h3e == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1265 = 6'h3f == architecturalRegMap_0; // @[decode.scala 388:24 392:{47,47}]
  wire  _GEN_1266 = 6'h0 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1267 = 6'h1 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1268 = 6'h2 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1269 = 6'h3 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1270 = 6'h4 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1271 = 6'h5 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1272 = 6'h6 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1273 = 6'h7 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1274 = 6'h8 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1275 = 6'h9 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1276 = 6'ha == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1277 = 6'hb == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1278 = 6'hc == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1279 = 6'hd == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1280 = 6'he == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1281 = 6'hf == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1282 = 6'h10 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1283 = 6'h11 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1284 = 6'h12 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1285 = 6'h13 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1286 = 6'h14 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1287 = 6'h15 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1288 = 6'h16 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1289 = 6'h17 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1290 = 6'h18 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1291 = 6'h19 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1292 = 6'h1a == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1293 = 6'h1b == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1294 = 6'h1c == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1295 = 6'h1d == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1296 = 6'h1e == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1297 = 6'h1f == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1298 = 6'h20 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1299 = 6'h21 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1300 = 6'h22 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1301 = 6'h23 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1302 = 6'h24 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1303 = 6'h25 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1304 = 6'h26 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1305 = 6'h27 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1306 = 6'h28 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1307 = 6'h29 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1308 = 6'h2a == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1309 = 6'h2b == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1310 = 6'h2c == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1311 = 6'h2d == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1312 = 6'h2e == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1313 = 6'h2f == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1314 = 6'h30 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1315 = 6'h31 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1316 = 6'h32 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1317 = 6'h33 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1318 = 6'h34 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1319 = 6'h35 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1320 = 6'h36 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1321 = 6'h37 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1322 = 6'h38 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1323 = 6'h39 == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1324 = 6'h3a == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1325 = 6'h3b == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1326 = 6'h3c == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1327 = 6'h3d == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1328 = 6'h3e == architecturalRegMap_0 ? 1'h0 : 1'h1; // @[decode.scala 387:24 393:{46,46}]
  wire  _GEN_1394 = 6'h0 == architecturalRegMap_1 ? 1'h0 : _GEN_1266; // @[decode.scala 393:{46,46}]
  wire  _GEN_1395 = 6'h1 == architecturalRegMap_1 ? 1'h0 : _GEN_1267; // @[decode.scala 393:{46,46}]
  wire  _GEN_1396 = 6'h2 == architecturalRegMap_1 ? 1'h0 : _GEN_1268; // @[decode.scala 393:{46,46}]
  wire  _GEN_1397 = 6'h3 == architecturalRegMap_1 ? 1'h0 : _GEN_1269; // @[decode.scala 393:{46,46}]
  wire  _GEN_1398 = 6'h4 == architecturalRegMap_1 ? 1'h0 : _GEN_1270; // @[decode.scala 393:{46,46}]
  wire  _GEN_1399 = 6'h5 == architecturalRegMap_1 ? 1'h0 : _GEN_1271; // @[decode.scala 393:{46,46}]
  wire  _GEN_1400 = 6'h6 == architecturalRegMap_1 ? 1'h0 : _GEN_1272; // @[decode.scala 393:{46,46}]
  wire  _GEN_1401 = 6'h7 == architecturalRegMap_1 ? 1'h0 : _GEN_1273; // @[decode.scala 393:{46,46}]
  wire  _GEN_1402 = 6'h8 == architecturalRegMap_1 ? 1'h0 : _GEN_1274; // @[decode.scala 393:{46,46}]
  wire  _GEN_1403 = 6'h9 == architecturalRegMap_1 ? 1'h0 : _GEN_1275; // @[decode.scala 393:{46,46}]
  wire  _GEN_1404 = 6'ha == architecturalRegMap_1 ? 1'h0 : _GEN_1276; // @[decode.scala 393:{46,46}]
  wire  _GEN_1405 = 6'hb == architecturalRegMap_1 ? 1'h0 : _GEN_1277; // @[decode.scala 393:{46,46}]
  wire  _GEN_1406 = 6'hc == architecturalRegMap_1 ? 1'h0 : _GEN_1278; // @[decode.scala 393:{46,46}]
  wire  _GEN_1407 = 6'hd == architecturalRegMap_1 ? 1'h0 : _GEN_1279; // @[decode.scala 393:{46,46}]
  wire  _GEN_1408 = 6'he == architecturalRegMap_1 ? 1'h0 : _GEN_1280; // @[decode.scala 393:{46,46}]
  wire  _GEN_1409 = 6'hf == architecturalRegMap_1 ? 1'h0 : _GEN_1281; // @[decode.scala 393:{46,46}]
  wire  _GEN_1410 = 6'h10 == architecturalRegMap_1 ? 1'h0 : _GEN_1282; // @[decode.scala 393:{46,46}]
  wire  _GEN_1411 = 6'h11 == architecturalRegMap_1 ? 1'h0 : _GEN_1283; // @[decode.scala 393:{46,46}]
  wire  _GEN_1412 = 6'h12 == architecturalRegMap_1 ? 1'h0 : _GEN_1284; // @[decode.scala 393:{46,46}]
  wire  _GEN_1413 = 6'h13 == architecturalRegMap_1 ? 1'h0 : _GEN_1285; // @[decode.scala 393:{46,46}]
  wire  _GEN_1414 = 6'h14 == architecturalRegMap_1 ? 1'h0 : _GEN_1286; // @[decode.scala 393:{46,46}]
  wire  _GEN_1415 = 6'h15 == architecturalRegMap_1 ? 1'h0 : _GEN_1287; // @[decode.scala 393:{46,46}]
  wire  _GEN_1416 = 6'h16 == architecturalRegMap_1 ? 1'h0 : _GEN_1288; // @[decode.scala 393:{46,46}]
  wire  _GEN_1417 = 6'h17 == architecturalRegMap_1 ? 1'h0 : _GEN_1289; // @[decode.scala 393:{46,46}]
  wire  _GEN_1418 = 6'h18 == architecturalRegMap_1 ? 1'h0 : _GEN_1290; // @[decode.scala 393:{46,46}]
  wire  _GEN_1419 = 6'h19 == architecturalRegMap_1 ? 1'h0 : _GEN_1291; // @[decode.scala 393:{46,46}]
  wire  _GEN_1420 = 6'h1a == architecturalRegMap_1 ? 1'h0 : _GEN_1292; // @[decode.scala 393:{46,46}]
  wire  _GEN_1421 = 6'h1b == architecturalRegMap_1 ? 1'h0 : _GEN_1293; // @[decode.scala 393:{46,46}]
  wire  _GEN_1422 = 6'h1c == architecturalRegMap_1 ? 1'h0 : _GEN_1294; // @[decode.scala 393:{46,46}]
  wire  _GEN_1423 = 6'h1d == architecturalRegMap_1 ? 1'h0 : _GEN_1295; // @[decode.scala 393:{46,46}]
  wire  _GEN_1424 = 6'h1e == architecturalRegMap_1 ? 1'h0 : _GEN_1296; // @[decode.scala 393:{46,46}]
  wire  _GEN_1425 = 6'h1f == architecturalRegMap_1 ? 1'h0 : _GEN_1297; // @[decode.scala 393:{46,46}]
  wire  _GEN_1426 = 6'h20 == architecturalRegMap_1 ? 1'h0 : _GEN_1298; // @[decode.scala 393:{46,46}]
  wire  _GEN_1427 = 6'h21 == architecturalRegMap_1 ? 1'h0 : _GEN_1299; // @[decode.scala 393:{46,46}]
  wire  _GEN_1428 = 6'h22 == architecturalRegMap_1 ? 1'h0 : _GEN_1300; // @[decode.scala 393:{46,46}]
  wire  _GEN_1429 = 6'h23 == architecturalRegMap_1 ? 1'h0 : _GEN_1301; // @[decode.scala 393:{46,46}]
  wire  _GEN_1430 = 6'h24 == architecturalRegMap_1 ? 1'h0 : _GEN_1302; // @[decode.scala 393:{46,46}]
  wire  _GEN_1431 = 6'h25 == architecturalRegMap_1 ? 1'h0 : _GEN_1303; // @[decode.scala 393:{46,46}]
  wire  _GEN_1432 = 6'h26 == architecturalRegMap_1 ? 1'h0 : _GEN_1304; // @[decode.scala 393:{46,46}]
  wire  _GEN_1433 = 6'h27 == architecturalRegMap_1 ? 1'h0 : _GEN_1305; // @[decode.scala 393:{46,46}]
  wire  _GEN_1434 = 6'h28 == architecturalRegMap_1 ? 1'h0 : _GEN_1306; // @[decode.scala 393:{46,46}]
  wire  _GEN_1435 = 6'h29 == architecturalRegMap_1 ? 1'h0 : _GEN_1307; // @[decode.scala 393:{46,46}]
  wire  _GEN_1436 = 6'h2a == architecturalRegMap_1 ? 1'h0 : _GEN_1308; // @[decode.scala 393:{46,46}]
  wire  _GEN_1437 = 6'h2b == architecturalRegMap_1 ? 1'h0 : _GEN_1309; // @[decode.scala 393:{46,46}]
  wire  _GEN_1438 = 6'h2c == architecturalRegMap_1 ? 1'h0 : _GEN_1310; // @[decode.scala 393:{46,46}]
  wire  _GEN_1439 = 6'h2d == architecturalRegMap_1 ? 1'h0 : _GEN_1311; // @[decode.scala 393:{46,46}]
  wire  _GEN_1440 = 6'h2e == architecturalRegMap_1 ? 1'h0 : _GEN_1312; // @[decode.scala 393:{46,46}]
  wire  _GEN_1441 = 6'h2f == architecturalRegMap_1 ? 1'h0 : _GEN_1313; // @[decode.scala 393:{46,46}]
  wire  _GEN_1442 = 6'h30 == architecturalRegMap_1 ? 1'h0 : _GEN_1314; // @[decode.scala 393:{46,46}]
  wire  _GEN_1443 = 6'h31 == architecturalRegMap_1 ? 1'h0 : _GEN_1315; // @[decode.scala 393:{46,46}]
  wire  _GEN_1444 = 6'h32 == architecturalRegMap_1 ? 1'h0 : _GEN_1316; // @[decode.scala 393:{46,46}]
  wire  _GEN_1445 = 6'h33 == architecturalRegMap_1 ? 1'h0 : _GEN_1317; // @[decode.scala 393:{46,46}]
  wire  _GEN_1446 = 6'h34 == architecturalRegMap_1 ? 1'h0 : _GEN_1318; // @[decode.scala 393:{46,46}]
  wire  _GEN_1447 = 6'h35 == architecturalRegMap_1 ? 1'h0 : _GEN_1319; // @[decode.scala 393:{46,46}]
  wire  _GEN_1448 = 6'h36 == architecturalRegMap_1 ? 1'h0 : _GEN_1320; // @[decode.scala 393:{46,46}]
  wire  _GEN_1449 = 6'h37 == architecturalRegMap_1 ? 1'h0 : _GEN_1321; // @[decode.scala 393:{46,46}]
  wire  _GEN_1450 = 6'h38 == architecturalRegMap_1 ? 1'h0 : _GEN_1322; // @[decode.scala 393:{46,46}]
  wire  _GEN_1451 = 6'h39 == architecturalRegMap_1 ? 1'h0 : _GEN_1323; // @[decode.scala 393:{46,46}]
  wire  _GEN_1452 = 6'h3a == architecturalRegMap_1 ? 1'h0 : _GEN_1324; // @[decode.scala 393:{46,46}]
  wire  _GEN_1453 = 6'h3b == architecturalRegMap_1 ? 1'h0 : _GEN_1325; // @[decode.scala 393:{46,46}]
  wire  _GEN_1454 = 6'h3c == architecturalRegMap_1 ? 1'h0 : _GEN_1326; // @[decode.scala 393:{46,46}]
  wire  _GEN_1455 = 6'h3d == architecturalRegMap_1 ? 1'h0 : _GEN_1327; // @[decode.scala 393:{46,46}]
  wire  _GEN_1456 = 6'h3e == architecturalRegMap_1 ? 1'h0 : _GEN_1328; // @[decode.scala 393:{46,46}]
  wire  _GEN_1522 = 6'h0 == architecturalRegMap_2 ? 1'h0 : _GEN_1394; // @[decode.scala 393:{46,46}]
  wire  _GEN_1523 = 6'h1 == architecturalRegMap_2 ? 1'h0 : _GEN_1395; // @[decode.scala 393:{46,46}]
  wire  _GEN_1524 = 6'h2 == architecturalRegMap_2 ? 1'h0 : _GEN_1396; // @[decode.scala 393:{46,46}]
  wire  _GEN_1525 = 6'h3 == architecturalRegMap_2 ? 1'h0 : _GEN_1397; // @[decode.scala 393:{46,46}]
  wire  _GEN_1526 = 6'h4 == architecturalRegMap_2 ? 1'h0 : _GEN_1398; // @[decode.scala 393:{46,46}]
  wire  _GEN_1527 = 6'h5 == architecturalRegMap_2 ? 1'h0 : _GEN_1399; // @[decode.scala 393:{46,46}]
  wire  _GEN_1528 = 6'h6 == architecturalRegMap_2 ? 1'h0 : _GEN_1400; // @[decode.scala 393:{46,46}]
  wire  _GEN_1529 = 6'h7 == architecturalRegMap_2 ? 1'h0 : _GEN_1401; // @[decode.scala 393:{46,46}]
  wire  _GEN_1530 = 6'h8 == architecturalRegMap_2 ? 1'h0 : _GEN_1402; // @[decode.scala 393:{46,46}]
  wire  _GEN_1531 = 6'h9 == architecturalRegMap_2 ? 1'h0 : _GEN_1403; // @[decode.scala 393:{46,46}]
  wire  _GEN_1532 = 6'ha == architecturalRegMap_2 ? 1'h0 : _GEN_1404; // @[decode.scala 393:{46,46}]
  wire  _GEN_1533 = 6'hb == architecturalRegMap_2 ? 1'h0 : _GEN_1405; // @[decode.scala 393:{46,46}]
  wire  _GEN_1534 = 6'hc == architecturalRegMap_2 ? 1'h0 : _GEN_1406; // @[decode.scala 393:{46,46}]
  wire  _GEN_1535 = 6'hd == architecturalRegMap_2 ? 1'h0 : _GEN_1407; // @[decode.scala 393:{46,46}]
  wire  _GEN_1536 = 6'he == architecturalRegMap_2 ? 1'h0 : _GEN_1408; // @[decode.scala 393:{46,46}]
  wire  _GEN_1537 = 6'hf == architecturalRegMap_2 ? 1'h0 : _GEN_1409; // @[decode.scala 393:{46,46}]
  wire  _GEN_1538 = 6'h10 == architecturalRegMap_2 ? 1'h0 : _GEN_1410; // @[decode.scala 393:{46,46}]
  wire  _GEN_1539 = 6'h11 == architecturalRegMap_2 ? 1'h0 : _GEN_1411; // @[decode.scala 393:{46,46}]
  wire  _GEN_1540 = 6'h12 == architecturalRegMap_2 ? 1'h0 : _GEN_1412; // @[decode.scala 393:{46,46}]
  wire  _GEN_1541 = 6'h13 == architecturalRegMap_2 ? 1'h0 : _GEN_1413; // @[decode.scala 393:{46,46}]
  wire  _GEN_1542 = 6'h14 == architecturalRegMap_2 ? 1'h0 : _GEN_1414; // @[decode.scala 393:{46,46}]
  wire  _GEN_1543 = 6'h15 == architecturalRegMap_2 ? 1'h0 : _GEN_1415; // @[decode.scala 393:{46,46}]
  wire  _GEN_1544 = 6'h16 == architecturalRegMap_2 ? 1'h0 : _GEN_1416; // @[decode.scala 393:{46,46}]
  wire  _GEN_1545 = 6'h17 == architecturalRegMap_2 ? 1'h0 : _GEN_1417; // @[decode.scala 393:{46,46}]
  wire  _GEN_1546 = 6'h18 == architecturalRegMap_2 ? 1'h0 : _GEN_1418; // @[decode.scala 393:{46,46}]
  wire  _GEN_1547 = 6'h19 == architecturalRegMap_2 ? 1'h0 : _GEN_1419; // @[decode.scala 393:{46,46}]
  wire  _GEN_1548 = 6'h1a == architecturalRegMap_2 ? 1'h0 : _GEN_1420; // @[decode.scala 393:{46,46}]
  wire  _GEN_1549 = 6'h1b == architecturalRegMap_2 ? 1'h0 : _GEN_1421; // @[decode.scala 393:{46,46}]
  wire  _GEN_1550 = 6'h1c == architecturalRegMap_2 ? 1'h0 : _GEN_1422; // @[decode.scala 393:{46,46}]
  wire  _GEN_1551 = 6'h1d == architecturalRegMap_2 ? 1'h0 : _GEN_1423; // @[decode.scala 393:{46,46}]
  wire  _GEN_1552 = 6'h1e == architecturalRegMap_2 ? 1'h0 : _GEN_1424; // @[decode.scala 393:{46,46}]
  wire  _GEN_1553 = 6'h1f == architecturalRegMap_2 ? 1'h0 : _GEN_1425; // @[decode.scala 393:{46,46}]
  wire  _GEN_1554 = 6'h20 == architecturalRegMap_2 ? 1'h0 : _GEN_1426; // @[decode.scala 393:{46,46}]
  wire  _GEN_1555 = 6'h21 == architecturalRegMap_2 ? 1'h0 : _GEN_1427; // @[decode.scala 393:{46,46}]
  wire  _GEN_1556 = 6'h22 == architecturalRegMap_2 ? 1'h0 : _GEN_1428; // @[decode.scala 393:{46,46}]
  wire  _GEN_1557 = 6'h23 == architecturalRegMap_2 ? 1'h0 : _GEN_1429; // @[decode.scala 393:{46,46}]
  wire  _GEN_1558 = 6'h24 == architecturalRegMap_2 ? 1'h0 : _GEN_1430; // @[decode.scala 393:{46,46}]
  wire  _GEN_1559 = 6'h25 == architecturalRegMap_2 ? 1'h0 : _GEN_1431; // @[decode.scala 393:{46,46}]
  wire  _GEN_1560 = 6'h26 == architecturalRegMap_2 ? 1'h0 : _GEN_1432; // @[decode.scala 393:{46,46}]
  wire  _GEN_1561 = 6'h27 == architecturalRegMap_2 ? 1'h0 : _GEN_1433; // @[decode.scala 393:{46,46}]
  wire  _GEN_1562 = 6'h28 == architecturalRegMap_2 ? 1'h0 : _GEN_1434; // @[decode.scala 393:{46,46}]
  wire  _GEN_1563 = 6'h29 == architecturalRegMap_2 ? 1'h0 : _GEN_1435; // @[decode.scala 393:{46,46}]
  wire  _GEN_1564 = 6'h2a == architecturalRegMap_2 ? 1'h0 : _GEN_1436; // @[decode.scala 393:{46,46}]
  wire  _GEN_1565 = 6'h2b == architecturalRegMap_2 ? 1'h0 : _GEN_1437; // @[decode.scala 393:{46,46}]
  wire  _GEN_1566 = 6'h2c == architecturalRegMap_2 ? 1'h0 : _GEN_1438; // @[decode.scala 393:{46,46}]
  wire  _GEN_1567 = 6'h2d == architecturalRegMap_2 ? 1'h0 : _GEN_1439; // @[decode.scala 393:{46,46}]
  wire  _GEN_1568 = 6'h2e == architecturalRegMap_2 ? 1'h0 : _GEN_1440; // @[decode.scala 393:{46,46}]
  wire  _GEN_1569 = 6'h2f == architecturalRegMap_2 ? 1'h0 : _GEN_1441; // @[decode.scala 393:{46,46}]
  wire  _GEN_1570 = 6'h30 == architecturalRegMap_2 ? 1'h0 : _GEN_1442; // @[decode.scala 393:{46,46}]
  wire  _GEN_1571 = 6'h31 == architecturalRegMap_2 ? 1'h0 : _GEN_1443; // @[decode.scala 393:{46,46}]
  wire  _GEN_1572 = 6'h32 == architecturalRegMap_2 ? 1'h0 : _GEN_1444; // @[decode.scala 393:{46,46}]
  wire  _GEN_1573 = 6'h33 == architecturalRegMap_2 ? 1'h0 : _GEN_1445; // @[decode.scala 393:{46,46}]
  wire  _GEN_1574 = 6'h34 == architecturalRegMap_2 ? 1'h0 : _GEN_1446; // @[decode.scala 393:{46,46}]
  wire  _GEN_1575 = 6'h35 == architecturalRegMap_2 ? 1'h0 : _GEN_1447; // @[decode.scala 393:{46,46}]
  wire  _GEN_1576 = 6'h36 == architecturalRegMap_2 ? 1'h0 : _GEN_1448; // @[decode.scala 393:{46,46}]
  wire  _GEN_1577 = 6'h37 == architecturalRegMap_2 ? 1'h0 : _GEN_1449; // @[decode.scala 393:{46,46}]
  wire  _GEN_1578 = 6'h38 == architecturalRegMap_2 ? 1'h0 : _GEN_1450; // @[decode.scala 393:{46,46}]
  wire  _GEN_1579 = 6'h39 == architecturalRegMap_2 ? 1'h0 : _GEN_1451; // @[decode.scala 393:{46,46}]
  wire  _GEN_1580 = 6'h3a == architecturalRegMap_2 ? 1'h0 : _GEN_1452; // @[decode.scala 393:{46,46}]
  wire  _GEN_1581 = 6'h3b == architecturalRegMap_2 ? 1'h0 : _GEN_1453; // @[decode.scala 393:{46,46}]
  wire  _GEN_1582 = 6'h3c == architecturalRegMap_2 ? 1'h0 : _GEN_1454; // @[decode.scala 393:{46,46}]
  wire  _GEN_1583 = 6'h3d == architecturalRegMap_2 ? 1'h0 : _GEN_1455; // @[decode.scala 393:{46,46}]
  wire  _GEN_1584 = 6'h3e == architecturalRegMap_2 ? 1'h0 : _GEN_1456; // @[decode.scala 393:{46,46}]
  wire  _GEN_1650 = 6'h0 == architecturalRegMap_3 ? 1'h0 : _GEN_1522; // @[decode.scala 393:{46,46}]
  wire  _GEN_1651 = 6'h1 == architecturalRegMap_3 ? 1'h0 : _GEN_1523; // @[decode.scala 393:{46,46}]
  wire  _GEN_1652 = 6'h2 == architecturalRegMap_3 ? 1'h0 : _GEN_1524; // @[decode.scala 393:{46,46}]
  wire  _GEN_1653 = 6'h3 == architecturalRegMap_3 ? 1'h0 : _GEN_1525; // @[decode.scala 393:{46,46}]
  wire  _GEN_1654 = 6'h4 == architecturalRegMap_3 ? 1'h0 : _GEN_1526; // @[decode.scala 393:{46,46}]
  wire  _GEN_1655 = 6'h5 == architecturalRegMap_3 ? 1'h0 : _GEN_1527; // @[decode.scala 393:{46,46}]
  wire  _GEN_1656 = 6'h6 == architecturalRegMap_3 ? 1'h0 : _GEN_1528; // @[decode.scala 393:{46,46}]
  wire  _GEN_1657 = 6'h7 == architecturalRegMap_3 ? 1'h0 : _GEN_1529; // @[decode.scala 393:{46,46}]
  wire  _GEN_1658 = 6'h8 == architecturalRegMap_3 ? 1'h0 : _GEN_1530; // @[decode.scala 393:{46,46}]
  wire  _GEN_1659 = 6'h9 == architecturalRegMap_3 ? 1'h0 : _GEN_1531; // @[decode.scala 393:{46,46}]
  wire  _GEN_1660 = 6'ha == architecturalRegMap_3 ? 1'h0 : _GEN_1532; // @[decode.scala 393:{46,46}]
  wire  _GEN_1661 = 6'hb == architecturalRegMap_3 ? 1'h0 : _GEN_1533; // @[decode.scala 393:{46,46}]
  wire  _GEN_1662 = 6'hc == architecturalRegMap_3 ? 1'h0 : _GEN_1534; // @[decode.scala 393:{46,46}]
  wire  _GEN_1663 = 6'hd == architecturalRegMap_3 ? 1'h0 : _GEN_1535; // @[decode.scala 393:{46,46}]
  wire  _GEN_1664 = 6'he == architecturalRegMap_3 ? 1'h0 : _GEN_1536; // @[decode.scala 393:{46,46}]
  wire  _GEN_1665 = 6'hf == architecturalRegMap_3 ? 1'h0 : _GEN_1537; // @[decode.scala 393:{46,46}]
  wire  _GEN_1666 = 6'h10 == architecturalRegMap_3 ? 1'h0 : _GEN_1538; // @[decode.scala 393:{46,46}]
  wire  _GEN_1667 = 6'h11 == architecturalRegMap_3 ? 1'h0 : _GEN_1539; // @[decode.scala 393:{46,46}]
  wire  _GEN_1668 = 6'h12 == architecturalRegMap_3 ? 1'h0 : _GEN_1540; // @[decode.scala 393:{46,46}]
  wire  _GEN_1669 = 6'h13 == architecturalRegMap_3 ? 1'h0 : _GEN_1541; // @[decode.scala 393:{46,46}]
  wire  _GEN_1670 = 6'h14 == architecturalRegMap_3 ? 1'h0 : _GEN_1542; // @[decode.scala 393:{46,46}]
  wire  _GEN_1671 = 6'h15 == architecturalRegMap_3 ? 1'h0 : _GEN_1543; // @[decode.scala 393:{46,46}]
  wire  _GEN_1672 = 6'h16 == architecturalRegMap_3 ? 1'h0 : _GEN_1544; // @[decode.scala 393:{46,46}]
  wire  _GEN_1673 = 6'h17 == architecturalRegMap_3 ? 1'h0 : _GEN_1545; // @[decode.scala 393:{46,46}]
  wire  _GEN_1674 = 6'h18 == architecturalRegMap_3 ? 1'h0 : _GEN_1546; // @[decode.scala 393:{46,46}]
  wire  _GEN_1675 = 6'h19 == architecturalRegMap_3 ? 1'h0 : _GEN_1547; // @[decode.scala 393:{46,46}]
  wire  _GEN_1676 = 6'h1a == architecturalRegMap_3 ? 1'h0 : _GEN_1548; // @[decode.scala 393:{46,46}]
  wire  _GEN_1677 = 6'h1b == architecturalRegMap_3 ? 1'h0 : _GEN_1549; // @[decode.scala 393:{46,46}]
  wire  _GEN_1678 = 6'h1c == architecturalRegMap_3 ? 1'h0 : _GEN_1550; // @[decode.scala 393:{46,46}]
  wire  _GEN_1679 = 6'h1d == architecturalRegMap_3 ? 1'h0 : _GEN_1551; // @[decode.scala 393:{46,46}]
  wire  _GEN_1680 = 6'h1e == architecturalRegMap_3 ? 1'h0 : _GEN_1552; // @[decode.scala 393:{46,46}]
  wire  _GEN_1681 = 6'h1f == architecturalRegMap_3 ? 1'h0 : _GEN_1553; // @[decode.scala 393:{46,46}]
  wire  _GEN_1682 = 6'h20 == architecturalRegMap_3 ? 1'h0 : _GEN_1554; // @[decode.scala 393:{46,46}]
  wire  _GEN_1683 = 6'h21 == architecturalRegMap_3 ? 1'h0 : _GEN_1555; // @[decode.scala 393:{46,46}]
  wire  _GEN_1684 = 6'h22 == architecturalRegMap_3 ? 1'h0 : _GEN_1556; // @[decode.scala 393:{46,46}]
  wire  _GEN_1685 = 6'h23 == architecturalRegMap_3 ? 1'h0 : _GEN_1557; // @[decode.scala 393:{46,46}]
  wire  _GEN_1686 = 6'h24 == architecturalRegMap_3 ? 1'h0 : _GEN_1558; // @[decode.scala 393:{46,46}]
  wire  _GEN_1687 = 6'h25 == architecturalRegMap_3 ? 1'h0 : _GEN_1559; // @[decode.scala 393:{46,46}]
  wire  _GEN_1688 = 6'h26 == architecturalRegMap_3 ? 1'h0 : _GEN_1560; // @[decode.scala 393:{46,46}]
  wire  _GEN_1689 = 6'h27 == architecturalRegMap_3 ? 1'h0 : _GEN_1561; // @[decode.scala 393:{46,46}]
  wire  _GEN_1690 = 6'h28 == architecturalRegMap_3 ? 1'h0 : _GEN_1562; // @[decode.scala 393:{46,46}]
  wire  _GEN_1691 = 6'h29 == architecturalRegMap_3 ? 1'h0 : _GEN_1563; // @[decode.scala 393:{46,46}]
  wire  _GEN_1692 = 6'h2a == architecturalRegMap_3 ? 1'h0 : _GEN_1564; // @[decode.scala 393:{46,46}]
  wire  _GEN_1693 = 6'h2b == architecturalRegMap_3 ? 1'h0 : _GEN_1565; // @[decode.scala 393:{46,46}]
  wire  _GEN_1694 = 6'h2c == architecturalRegMap_3 ? 1'h0 : _GEN_1566; // @[decode.scala 393:{46,46}]
  wire  _GEN_1695 = 6'h2d == architecturalRegMap_3 ? 1'h0 : _GEN_1567; // @[decode.scala 393:{46,46}]
  wire  _GEN_1696 = 6'h2e == architecturalRegMap_3 ? 1'h0 : _GEN_1568; // @[decode.scala 393:{46,46}]
  wire  _GEN_1697 = 6'h2f == architecturalRegMap_3 ? 1'h0 : _GEN_1569; // @[decode.scala 393:{46,46}]
  wire  _GEN_1698 = 6'h30 == architecturalRegMap_3 ? 1'h0 : _GEN_1570; // @[decode.scala 393:{46,46}]
  wire  _GEN_1699 = 6'h31 == architecturalRegMap_3 ? 1'h0 : _GEN_1571; // @[decode.scala 393:{46,46}]
  wire  _GEN_1700 = 6'h32 == architecturalRegMap_3 ? 1'h0 : _GEN_1572; // @[decode.scala 393:{46,46}]
  wire  _GEN_1701 = 6'h33 == architecturalRegMap_3 ? 1'h0 : _GEN_1573; // @[decode.scala 393:{46,46}]
  wire  _GEN_1702 = 6'h34 == architecturalRegMap_3 ? 1'h0 : _GEN_1574; // @[decode.scala 393:{46,46}]
  wire  _GEN_1703 = 6'h35 == architecturalRegMap_3 ? 1'h0 : _GEN_1575; // @[decode.scala 393:{46,46}]
  wire  _GEN_1704 = 6'h36 == architecturalRegMap_3 ? 1'h0 : _GEN_1576; // @[decode.scala 393:{46,46}]
  wire  _GEN_1705 = 6'h37 == architecturalRegMap_3 ? 1'h0 : _GEN_1577; // @[decode.scala 393:{46,46}]
  wire  _GEN_1706 = 6'h38 == architecturalRegMap_3 ? 1'h0 : _GEN_1578; // @[decode.scala 393:{46,46}]
  wire  _GEN_1707 = 6'h39 == architecturalRegMap_3 ? 1'h0 : _GEN_1579; // @[decode.scala 393:{46,46}]
  wire  _GEN_1708 = 6'h3a == architecturalRegMap_3 ? 1'h0 : _GEN_1580; // @[decode.scala 393:{46,46}]
  wire  _GEN_1709 = 6'h3b == architecturalRegMap_3 ? 1'h0 : _GEN_1581; // @[decode.scala 393:{46,46}]
  wire  _GEN_1710 = 6'h3c == architecturalRegMap_3 ? 1'h0 : _GEN_1582; // @[decode.scala 393:{46,46}]
  wire  _GEN_1711 = 6'h3d == architecturalRegMap_3 ? 1'h0 : _GEN_1583; // @[decode.scala 393:{46,46}]
  wire  _GEN_1712 = 6'h3e == architecturalRegMap_3 ? 1'h0 : _GEN_1584; // @[decode.scala 393:{46,46}]
  wire  _GEN_1778 = 6'h0 == architecturalRegMap_4 ? 1'h0 : _GEN_1650; // @[decode.scala 393:{46,46}]
  wire  _GEN_1779 = 6'h1 == architecturalRegMap_4 ? 1'h0 : _GEN_1651; // @[decode.scala 393:{46,46}]
  wire  _GEN_1780 = 6'h2 == architecturalRegMap_4 ? 1'h0 : _GEN_1652; // @[decode.scala 393:{46,46}]
  wire  _GEN_1781 = 6'h3 == architecturalRegMap_4 ? 1'h0 : _GEN_1653; // @[decode.scala 393:{46,46}]
  wire  _GEN_1782 = 6'h4 == architecturalRegMap_4 ? 1'h0 : _GEN_1654; // @[decode.scala 393:{46,46}]
  wire  _GEN_1783 = 6'h5 == architecturalRegMap_4 ? 1'h0 : _GEN_1655; // @[decode.scala 393:{46,46}]
  wire  _GEN_1784 = 6'h6 == architecturalRegMap_4 ? 1'h0 : _GEN_1656; // @[decode.scala 393:{46,46}]
  wire  _GEN_1785 = 6'h7 == architecturalRegMap_4 ? 1'h0 : _GEN_1657; // @[decode.scala 393:{46,46}]
  wire  _GEN_1786 = 6'h8 == architecturalRegMap_4 ? 1'h0 : _GEN_1658; // @[decode.scala 393:{46,46}]
  wire  _GEN_1787 = 6'h9 == architecturalRegMap_4 ? 1'h0 : _GEN_1659; // @[decode.scala 393:{46,46}]
  wire  _GEN_1788 = 6'ha == architecturalRegMap_4 ? 1'h0 : _GEN_1660; // @[decode.scala 393:{46,46}]
  wire  _GEN_1789 = 6'hb == architecturalRegMap_4 ? 1'h0 : _GEN_1661; // @[decode.scala 393:{46,46}]
  wire  _GEN_1790 = 6'hc == architecturalRegMap_4 ? 1'h0 : _GEN_1662; // @[decode.scala 393:{46,46}]
  wire  _GEN_1791 = 6'hd == architecturalRegMap_4 ? 1'h0 : _GEN_1663; // @[decode.scala 393:{46,46}]
  wire  _GEN_1792 = 6'he == architecturalRegMap_4 ? 1'h0 : _GEN_1664; // @[decode.scala 393:{46,46}]
  wire  _GEN_1793 = 6'hf == architecturalRegMap_4 ? 1'h0 : _GEN_1665; // @[decode.scala 393:{46,46}]
  wire  _GEN_1794 = 6'h10 == architecturalRegMap_4 ? 1'h0 : _GEN_1666; // @[decode.scala 393:{46,46}]
  wire  _GEN_1795 = 6'h11 == architecturalRegMap_4 ? 1'h0 : _GEN_1667; // @[decode.scala 393:{46,46}]
  wire  _GEN_1796 = 6'h12 == architecturalRegMap_4 ? 1'h0 : _GEN_1668; // @[decode.scala 393:{46,46}]
  wire  _GEN_1797 = 6'h13 == architecturalRegMap_4 ? 1'h0 : _GEN_1669; // @[decode.scala 393:{46,46}]
  wire  _GEN_1798 = 6'h14 == architecturalRegMap_4 ? 1'h0 : _GEN_1670; // @[decode.scala 393:{46,46}]
  wire  _GEN_1799 = 6'h15 == architecturalRegMap_4 ? 1'h0 : _GEN_1671; // @[decode.scala 393:{46,46}]
  wire  _GEN_1800 = 6'h16 == architecturalRegMap_4 ? 1'h0 : _GEN_1672; // @[decode.scala 393:{46,46}]
  wire  _GEN_1801 = 6'h17 == architecturalRegMap_4 ? 1'h0 : _GEN_1673; // @[decode.scala 393:{46,46}]
  wire  _GEN_1802 = 6'h18 == architecturalRegMap_4 ? 1'h0 : _GEN_1674; // @[decode.scala 393:{46,46}]
  wire  _GEN_1803 = 6'h19 == architecturalRegMap_4 ? 1'h0 : _GEN_1675; // @[decode.scala 393:{46,46}]
  wire  _GEN_1804 = 6'h1a == architecturalRegMap_4 ? 1'h0 : _GEN_1676; // @[decode.scala 393:{46,46}]
  wire  _GEN_1805 = 6'h1b == architecturalRegMap_4 ? 1'h0 : _GEN_1677; // @[decode.scala 393:{46,46}]
  wire  _GEN_1806 = 6'h1c == architecturalRegMap_4 ? 1'h0 : _GEN_1678; // @[decode.scala 393:{46,46}]
  wire  _GEN_1807 = 6'h1d == architecturalRegMap_4 ? 1'h0 : _GEN_1679; // @[decode.scala 393:{46,46}]
  wire  _GEN_1808 = 6'h1e == architecturalRegMap_4 ? 1'h0 : _GEN_1680; // @[decode.scala 393:{46,46}]
  wire  _GEN_1809 = 6'h1f == architecturalRegMap_4 ? 1'h0 : _GEN_1681; // @[decode.scala 393:{46,46}]
  wire  _GEN_1810 = 6'h20 == architecturalRegMap_4 ? 1'h0 : _GEN_1682; // @[decode.scala 393:{46,46}]
  wire  _GEN_1811 = 6'h21 == architecturalRegMap_4 ? 1'h0 : _GEN_1683; // @[decode.scala 393:{46,46}]
  wire  _GEN_1812 = 6'h22 == architecturalRegMap_4 ? 1'h0 : _GEN_1684; // @[decode.scala 393:{46,46}]
  wire  _GEN_1813 = 6'h23 == architecturalRegMap_4 ? 1'h0 : _GEN_1685; // @[decode.scala 393:{46,46}]
  wire  _GEN_1814 = 6'h24 == architecturalRegMap_4 ? 1'h0 : _GEN_1686; // @[decode.scala 393:{46,46}]
  wire  _GEN_1815 = 6'h25 == architecturalRegMap_4 ? 1'h0 : _GEN_1687; // @[decode.scala 393:{46,46}]
  wire  _GEN_1816 = 6'h26 == architecturalRegMap_4 ? 1'h0 : _GEN_1688; // @[decode.scala 393:{46,46}]
  wire  _GEN_1817 = 6'h27 == architecturalRegMap_4 ? 1'h0 : _GEN_1689; // @[decode.scala 393:{46,46}]
  wire  _GEN_1818 = 6'h28 == architecturalRegMap_4 ? 1'h0 : _GEN_1690; // @[decode.scala 393:{46,46}]
  wire  _GEN_1819 = 6'h29 == architecturalRegMap_4 ? 1'h0 : _GEN_1691; // @[decode.scala 393:{46,46}]
  wire  _GEN_1820 = 6'h2a == architecturalRegMap_4 ? 1'h0 : _GEN_1692; // @[decode.scala 393:{46,46}]
  wire  _GEN_1821 = 6'h2b == architecturalRegMap_4 ? 1'h0 : _GEN_1693; // @[decode.scala 393:{46,46}]
  wire  _GEN_1822 = 6'h2c == architecturalRegMap_4 ? 1'h0 : _GEN_1694; // @[decode.scala 393:{46,46}]
  wire  _GEN_1823 = 6'h2d == architecturalRegMap_4 ? 1'h0 : _GEN_1695; // @[decode.scala 393:{46,46}]
  wire  _GEN_1824 = 6'h2e == architecturalRegMap_4 ? 1'h0 : _GEN_1696; // @[decode.scala 393:{46,46}]
  wire  _GEN_1825 = 6'h2f == architecturalRegMap_4 ? 1'h0 : _GEN_1697; // @[decode.scala 393:{46,46}]
  wire  _GEN_1826 = 6'h30 == architecturalRegMap_4 ? 1'h0 : _GEN_1698; // @[decode.scala 393:{46,46}]
  wire  _GEN_1827 = 6'h31 == architecturalRegMap_4 ? 1'h0 : _GEN_1699; // @[decode.scala 393:{46,46}]
  wire  _GEN_1828 = 6'h32 == architecturalRegMap_4 ? 1'h0 : _GEN_1700; // @[decode.scala 393:{46,46}]
  wire  _GEN_1829 = 6'h33 == architecturalRegMap_4 ? 1'h0 : _GEN_1701; // @[decode.scala 393:{46,46}]
  wire  _GEN_1830 = 6'h34 == architecturalRegMap_4 ? 1'h0 : _GEN_1702; // @[decode.scala 393:{46,46}]
  wire  _GEN_1831 = 6'h35 == architecturalRegMap_4 ? 1'h0 : _GEN_1703; // @[decode.scala 393:{46,46}]
  wire  _GEN_1832 = 6'h36 == architecturalRegMap_4 ? 1'h0 : _GEN_1704; // @[decode.scala 393:{46,46}]
  wire  _GEN_1833 = 6'h37 == architecturalRegMap_4 ? 1'h0 : _GEN_1705; // @[decode.scala 393:{46,46}]
  wire  _GEN_1834 = 6'h38 == architecturalRegMap_4 ? 1'h0 : _GEN_1706; // @[decode.scala 393:{46,46}]
  wire  _GEN_1835 = 6'h39 == architecturalRegMap_4 ? 1'h0 : _GEN_1707; // @[decode.scala 393:{46,46}]
  wire  _GEN_1836 = 6'h3a == architecturalRegMap_4 ? 1'h0 : _GEN_1708; // @[decode.scala 393:{46,46}]
  wire  _GEN_1837 = 6'h3b == architecturalRegMap_4 ? 1'h0 : _GEN_1709; // @[decode.scala 393:{46,46}]
  wire  _GEN_1838 = 6'h3c == architecturalRegMap_4 ? 1'h0 : _GEN_1710; // @[decode.scala 393:{46,46}]
  wire  _GEN_1839 = 6'h3d == architecturalRegMap_4 ? 1'h0 : _GEN_1711; // @[decode.scala 393:{46,46}]
  wire  _GEN_1840 = 6'h3e == architecturalRegMap_4 ? 1'h0 : _GEN_1712; // @[decode.scala 393:{46,46}]
  wire  _GEN_1906 = 6'h0 == architecturalRegMap_5 ? 1'h0 : _GEN_1778; // @[decode.scala 393:{46,46}]
  wire  _GEN_1907 = 6'h1 == architecturalRegMap_5 ? 1'h0 : _GEN_1779; // @[decode.scala 393:{46,46}]
  wire  _GEN_1908 = 6'h2 == architecturalRegMap_5 ? 1'h0 : _GEN_1780; // @[decode.scala 393:{46,46}]
  wire  _GEN_1909 = 6'h3 == architecturalRegMap_5 ? 1'h0 : _GEN_1781; // @[decode.scala 393:{46,46}]
  wire  _GEN_1910 = 6'h4 == architecturalRegMap_5 ? 1'h0 : _GEN_1782; // @[decode.scala 393:{46,46}]
  wire  _GEN_1911 = 6'h5 == architecturalRegMap_5 ? 1'h0 : _GEN_1783; // @[decode.scala 393:{46,46}]
  wire  _GEN_1912 = 6'h6 == architecturalRegMap_5 ? 1'h0 : _GEN_1784; // @[decode.scala 393:{46,46}]
  wire  _GEN_1913 = 6'h7 == architecturalRegMap_5 ? 1'h0 : _GEN_1785; // @[decode.scala 393:{46,46}]
  wire  _GEN_1914 = 6'h8 == architecturalRegMap_5 ? 1'h0 : _GEN_1786; // @[decode.scala 393:{46,46}]
  wire  _GEN_1915 = 6'h9 == architecturalRegMap_5 ? 1'h0 : _GEN_1787; // @[decode.scala 393:{46,46}]
  wire  _GEN_1916 = 6'ha == architecturalRegMap_5 ? 1'h0 : _GEN_1788; // @[decode.scala 393:{46,46}]
  wire  _GEN_1917 = 6'hb == architecturalRegMap_5 ? 1'h0 : _GEN_1789; // @[decode.scala 393:{46,46}]
  wire  _GEN_1918 = 6'hc == architecturalRegMap_5 ? 1'h0 : _GEN_1790; // @[decode.scala 393:{46,46}]
  wire  _GEN_1919 = 6'hd == architecturalRegMap_5 ? 1'h0 : _GEN_1791; // @[decode.scala 393:{46,46}]
  wire  _GEN_1920 = 6'he == architecturalRegMap_5 ? 1'h0 : _GEN_1792; // @[decode.scala 393:{46,46}]
  wire  _GEN_1921 = 6'hf == architecturalRegMap_5 ? 1'h0 : _GEN_1793; // @[decode.scala 393:{46,46}]
  wire  _GEN_1922 = 6'h10 == architecturalRegMap_5 ? 1'h0 : _GEN_1794; // @[decode.scala 393:{46,46}]
  wire  _GEN_1923 = 6'h11 == architecturalRegMap_5 ? 1'h0 : _GEN_1795; // @[decode.scala 393:{46,46}]
  wire  _GEN_1924 = 6'h12 == architecturalRegMap_5 ? 1'h0 : _GEN_1796; // @[decode.scala 393:{46,46}]
  wire  _GEN_1925 = 6'h13 == architecturalRegMap_5 ? 1'h0 : _GEN_1797; // @[decode.scala 393:{46,46}]
  wire  _GEN_1926 = 6'h14 == architecturalRegMap_5 ? 1'h0 : _GEN_1798; // @[decode.scala 393:{46,46}]
  wire  _GEN_1927 = 6'h15 == architecturalRegMap_5 ? 1'h0 : _GEN_1799; // @[decode.scala 393:{46,46}]
  wire  _GEN_1928 = 6'h16 == architecturalRegMap_5 ? 1'h0 : _GEN_1800; // @[decode.scala 393:{46,46}]
  wire  _GEN_1929 = 6'h17 == architecturalRegMap_5 ? 1'h0 : _GEN_1801; // @[decode.scala 393:{46,46}]
  wire  _GEN_1930 = 6'h18 == architecturalRegMap_5 ? 1'h0 : _GEN_1802; // @[decode.scala 393:{46,46}]
  wire  _GEN_1931 = 6'h19 == architecturalRegMap_5 ? 1'h0 : _GEN_1803; // @[decode.scala 393:{46,46}]
  wire  _GEN_1932 = 6'h1a == architecturalRegMap_5 ? 1'h0 : _GEN_1804; // @[decode.scala 393:{46,46}]
  wire  _GEN_1933 = 6'h1b == architecturalRegMap_5 ? 1'h0 : _GEN_1805; // @[decode.scala 393:{46,46}]
  wire  _GEN_1934 = 6'h1c == architecturalRegMap_5 ? 1'h0 : _GEN_1806; // @[decode.scala 393:{46,46}]
  wire  _GEN_1935 = 6'h1d == architecturalRegMap_5 ? 1'h0 : _GEN_1807; // @[decode.scala 393:{46,46}]
  wire  _GEN_1936 = 6'h1e == architecturalRegMap_5 ? 1'h0 : _GEN_1808; // @[decode.scala 393:{46,46}]
  wire  _GEN_1937 = 6'h1f == architecturalRegMap_5 ? 1'h0 : _GEN_1809; // @[decode.scala 393:{46,46}]
  wire  _GEN_1938 = 6'h20 == architecturalRegMap_5 ? 1'h0 : _GEN_1810; // @[decode.scala 393:{46,46}]
  wire  _GEN_1939 = 6'h21 == architecturalRegMap_5 ? 1'h0 : _GEN_1811; // @[decode.scala 393:{46,46}]
  wire  _GEN_1940 = 6'h22 == architecturalRegMap_5 ? 1'h0 : _GEN_1812; // @[decode.scala 393:{46,46}]
  wire  _GEN_1941 = 6'h23 == architecturalRegMap_5 ? 1'h0 : _GEN_1813; // @[decode.scala 393:{46,46}]
  wire  _GEN_1942 = 6'h24 == architecturalRegMap_5 ? 1'h0 : _GEN_1814; // @[decode.scala 393:{46,46}]
  wire  _GEN_1943 = 6'h25 == architecturalRegMap_5 ? 1'h0 : _GEN_1815; // @[decode.scala 393:{46,46}]
  wire  _GEN_1944 = 6'h26 == architecturalRegMap_5 ? 1'h0 : _GEN_1816; // @[decode.scala 393:{46,46}]
  wire  _GEN_1945 = 6'h27 == architecturalRegMap_5 ? 1'h0 : _GEN_1817; // @[decode.scala 393:{46,46}]
  wire  _GEN_1946 = 6'h28 == architecturalRegMap_5 ? 1'h0 : _GEN_1818; // @[decode.scala 393:{46,46}]
  wire  _GEN_1947 = 6'h29 == architecturalRegMap_5 ? 1'h0 : _GEN_1819; // @[decode.scala 393:{46,46}]
  wire  _GEN_1948 = 6'h2a == architecturalRegMap_5 ? 1'h0 : _GEN_1820; // @[decode.scala 393:{46,46}]
  wire  _GEN_1949 = 6'h2b == architecturalRegMap_5 ? 1'h0 : _GEN_1821; // @[decode.scala 393:{46,46}]
  wire  _GEN_1950 = 6'h2c == architecturalRegMap_5 ? 1'h0 : _GEN_1822; // @[decode.scala 393:{46,46}]
  wire  _GEN_1951 = 6'h2d == architecturalRegMap_5 ? 1'h0 : _GEN_1823; // @[decode.scala 393:{46,46}]
  wire  _GEN_1952 = 6'h2e == architecturalRegMap_5 ? 1'h0 : _GEN_1824; // @[decode.scala 393:{46,46}]
  wire  _GEN_1953 = 6'h2f == architecturalRegMap_5 ? 1'h0 : _GEN_1825; // @[decode.scala 393:{46,46}]
  wire  _GEN_1954 = 6'h30 == architecturalRegMap_5 ? 1'h0 : _GEN_1826; // @[decode.scala 393:{46,46}]
  wire  _GEN_1955 = 6'h31 == architecturalRegMap_5 ? 1'h0 : _GEN_1827; // @[decode.scala 393:{46,46}]
  wire  _GEN_1956 = 6'h32 == architecturalRegMap_5 ? 1'h0 : _GEN_1828; // @[decode.scala 393:{46,46}]
  wire  _GEN_1957 = 6'h33 == architecturalRegMap_5 ? 1'h0 : _GEN_1829; // @[decode.scala 393:{46,46}]
  wire  _GEN_1958 = 6'h34 == architecturalRegMap_5 ? 1'h0 : _GEN_1830; // @[decode.scala 393:{46,46}]
  wire  _GEN_1959 = 6'h35 == architecturalRegMap_5 ? 1'h0 : _GEN_1831; // @[decode.scala 393:{46,46}]
  wire  _GEN_1960 = 6'h36 == architecturalRegMap_5 ? 1'h0 : _GEN_1832; // @[decode.scala 393:{46,46}]
  wire  _GEN_1961 = 6'h37 == architecturalRegMap_5 ? 1'h0 : _GEN_1833; // @[decode.scala 393:{46,46}]
  wire  _GEN_1962 = 6'h38 == architecturalRegMap_5 ? 1'h0 : _GEN_1834; // @[decode.scala 393:{46,46}]
  wire  _GEN_1963 = 6'h39 == architecturalRegMap_5 ? 1'h0 : _GEN_1835; // @[decode.scala 393:{46,46}]
  wire  _GEN_1964 = 6'h3a == architecturalRegMap_5 ? 1'h0 : _GEN_1836; // @[decode.scala 393:{46,46}]
  wire  _GEN_1965 = 6'h3b == architecturalRegMap_5 ? 1'h0 : _GEN_1837; // @[decode.scala 393:{46,46}]
  wire  _GEN_1966 = 6'h3c == architecturalRegMap_5 ? 1'h0 : _GEN_1838; // @[decode.scala 393:{46,46}]
  wire  _GEN_1967 = 6'h3d == architecturalRegMap_5 ? 1'h0 : _GEN_1839; // @[decode.scala 393:{46,46}]
  wire  _GEN_1968 = 6'h3e == architecturalRegMap_5 ? 1'h0 : _GEN_1840; // @[decode.scala 393:{46,46}]
  wire  _GEN_2034 = 6'h0 == architecturalRegMap_6 ? 1'h0 : _GEN_1906; // @[decode.scala 393:{46,46}]
  wire  _GEN_2035 = 6'h1 == architecturalRegMap_6 ? 1'h0 : _GEN_1907; // @[decode.scala 393:{46,46}]
  wire  _GEN_2036 = 6'h2 == architecturalRegMap_6 ? 1'h0 : _GEN_1908; // @[decode.scala 393:{46,46}]
  wire  _GEN_2037 = 6'h3 == architecturalRegMap_6 ? 1'h0 : _GEN_1909; // @[decode.scala 393:{46,46}]
  wire  _GEN_2038 = 6'h4 == architecturalRegMap_6 ? 1'h0 : _GEN_1910; // @[decode.scala 393:{46,46}]
  wire  _GEN_2039 = 6'h5 == architecturalRegMap_6 ? 1'h0 : _GEN_1911; // @[decode.scala 393:{46,46}]
  wire  _GEN_2040 = 6'h6 == architecturalRegMap_6 ? 1'h0 : _GEN_1912; // @[decode.scala 393:{46,46}]
  wire  _GEN_2041 = 6'h7 == architecturalRegMap_6 ? 1'h0 : _GEN_1913; // @[decode.scala 393:{46,46}]
  wire  _GEN_2042 = 6'h8 == architecturalRegMap_6 ? 1'h0 : _GEN_1914; // @[decode.scala 393:{46,46}]
  wire  _GEN_2043 = 6'h9 == architecturalRegMap_6 ? 1'h0 : _GEN_1915; // @[decode.scala 393:{46,46}]
  wire  _GEN_2044 = 6'ha == architecturalRegMap_6 ? 1'h0 : _GEN_1916; // @[decode.scala 393:{46,46}]
  wire  _GEN_2045 = 6'hb == architecturalRegMap_6 ? 1'h0 : _GEN_1917; // @[decode.scala 393:{46,46}]
  wire  _GEN_2046 = 6'hc == architecturalRegMap_6 ? 1'h0 : _GEN_1918; // @[decode.scala 393:{46,46}]
  wire  _GEN_2047 = 6'hd == architecturalRegMap_6 ? 1'h0 : _GEN_1919; // @[decode.scala 393:{46,46}]
  wire  _GEN_2048 = 6'he == architecturalRegMap_6 ? 1'h0 : _GEN_1920; // @[decode.scala 393:{46,46}]
  wire  _GEN_2049 = 6'hf == architecturalRegMap_6 ? 1'h0 : _GEN_1921; // @[decode.scala 393:{46,46}]
  wire  _GEN_2050 = 6'h10 == architecturalRegMap_6 ? 1'h0 : _GEN_1922; // @[decode.scala 393:{46,46}]
  wire  _GEN_2051 = 6'h11 == architecturalRegMap_6 ? 1'h0 : _GEN_1923; // @[decode.scala 393:{46,46}]
  wire  _GEN_2052 = 6'h12 == architecturalRegMap_6 ? 1'h0 : _GEN_1924; // @[decode.scala 393:{46,46}]
  wire  _GEN_2053 = 6'h13 == architecturalRegMap_6 ? 1'h0 : _GEN_1925; // @[decode.scala 393:{46,46}]
  wire  _GEN_2054 = 6'h14 == architecturalRegMap_6 ? 1'h0 : _GEN_1926; // @[decode.scala 393:{46,46}]
  wire  _GEN_2055 = 6'h15 == architecturalRegMap_6 ? 1'h0 : _GEN_1927; // @[decode.scala 393:{46,46}]
  wire  _GEN_2056 = 6'h16 == architecturalRegMap_6 ? 1'h0 : _GEN_1928; // @[decode.scala 393:{46,46}]
  wire  _GEN_2057 = 6'h17 == architecturalRegMap_6 ? 1'h0 : _GEN_1929; // @[decode.scala 393:{46,46}]
  wire  _GEN_2058 = 6'h18 == architecturalRegMap_6 ? 1'h0 : _GEN_1930; // @[decode.scala 393:{46,46}]
  wire  _GEN_2059 = 6'h19 == architecturalRegMap_6 ? 1'h0 : _GEN_1931; // @[decode.scala 393:{46,46}]
  wire  _GEN_2060 = 6'h1a == architecturalRegMap_6 ? 1'h0 : _GEN_1932; // @[decode.scala 393:{46,46}]
  wire  _GEN_2061 = 6'h1b == architecturalRegMap_6 ? 1'h0 : _GEN_1933; // @[decode.scala 393:{46,46}]
  wire  _GEN_2062 = 6'h1c == architecturalRegMap_6 ? 1'h0 : _GEN_1934; // @[decode.scala 393:{46,46}]
  wire  _GEN_2063 = 6'h1d == architecturalRegMap_6 ? 1'h0 : _GEN_1935; // @[decode.scala 393:{46,46}]
  wire  _GEN_2064 = 6'h1e == architecturalRegMap_6 ? 1'h0 : _GEN_1936; // @[decode.scala 393:{46,46}]
  wire  _GEN_2065 = 6'h1f == architecturalRegMap_6 ? 1'h0 : _GEN_1937; // @[decode.scala 393:{46,46}]
  wire  _GEN_2066 = 6'h20 == architecturalRegMap_6 ? 1'h0 : _GEN_1938; // @[decode.scala 393:{46,46}]
  wire  _GEN_2067 = 6'h21 == architecturalRegMap_6 ? 1'h0 : _GEN_1939; // @[decode.scala 393:{46,46}]
  wire  _GEN_2068 = 6'h22 == architecturalRegMap_6 ? 1'h0 : _GEN_1940; // @[decode.scala 393:{46,46}]
  wire  _GEN_2069 = 6'h23 == architecturalRegMap_6 ? 1'h0 : _GEN_1941; // @[decode.scala 393:{46,46}]
  wire  _GEN_2070 = 6'h24 == architecturalRegMap_6 ? 1'h0 : _GEN_1942; // @[decode.scala 393:{46,46}]
  wire  _GEN_2071 = 6'h25 == architecturalRegMap_6 ? 1'h0 : _GEN_1943; // @[decode.scala 393:{46,46}]
  wire  _GEN_2072 = 6'h26 == architecturalRegMap_6 ? 1'h0 : _GEN_1944; // @[decode.scala 393:{46,46}]
  wire  _GEN_2073 = 6'h27 == architecturalRegMap_6 ? 1'h0 : _GEN_1945; // @[decode.scala 393:{46,46}]
  wire  _GEN_2074 = 6'h28 == architecturalRegMap_6 ? 1'h0 : _GEN_1946; // @[decode.scala 393:{46,46}]
  wire  _GEN_2075 = 6'h29 == architecturalRegMap_6 ? 1'h0 : _GEN_1947; // @[decode.scala 393:{46,46}]
  wire  _GEN_2076 = 6'h2a == architecturalRegMap_6 ? 1'h0 : _GEN_1948; // @[decode.scala 393:{46,46}]
  wire  _GEN_2077 = 6'h2b == architecturalRegMap_6 ? 1'h0 : _GEN_1949; // @[decode.scala 393:{46,46}]
  wire  _GEN_2078 = 6'h2c == architecturalRegMap_6 ? 1'h0 : _GEN_1950; // @[decode.scala 393:{46,46}]
  wire  _GEN_2079 = 6'h2d == architecturalRegMap_6 ? 1'h0 : _GEN_1951; // @[decode.scala 393:{46,46}]
  wire  _GEN_2080 = 6'h2e == architecturalRegMap_6 ? 1'h0 : _GEN_1952; // @[decode.scala 393:{46,46}]
  wire  _GEN_2081 = 6'h2f == architecturalRegMap_6 ? 1'h0 : _GEN_1953; // @[decode.scala 393:{46,46}]
  wire  _GEN_2082 = 6'h30 == architecturalRegMap_6 ? 1'h0 : _GEN_1954; // @[decode.scala 393:{46,46}]
  wire  _GEN_2083 = 6'h31 == architecturalRegMap_6 ? 1'h0 : _GEN_1955; // @[decode.scala 393:{46,46}]
  wire  _GEN_2084 = 6'h32 == architecturalRegMap_6 ? 1'h0 : _GEN_1956; // @[decode.scala 393:{46,46}]
  wire  _GEN_2085 = 6'h33 == architecturalRegMap_6 ? 1'h0 : _GEN_1957; // @[decode.scala 393:{46,46}]
  wire  _GEN_2086 = 6'h34 == architecturalRegMap_6 ? 1'h0 : _GEN_1958; // @[decode.scala 393:{46,46}]
  wire  _GEN_2087 = 6'h35 == architecturalRegMap_6 ? 1'h0 : _GEN_1959; // @[decode.scala 393:{46,46}]
  wire  _GEN_2088 = 6'h36 == architecturalRegMap_6 ? 1'h0 : _GEN_1960; // @[decode.scala 393:{46,46}]
  wire  _GEN_2089 = 6'h37 == architecturalRegMap_6 ? 1'h0 : _GEN_1961; // @[decode.scala 393:{46,46}]
  wire  _GEN_2090 = 6'h38 == architecturalRegMap_6 ? 1'h0 : _GEN_1962; // @[decode.scala 393:{46,46}]
  wire  _GEN_2091 = 6'h39 == architecturalRegMap_6 ? 1'h0 : _GEN_1963; // @[decode.scala 393:{46,46}]
  wire  _GEN_2092 = 6'h3a == architecturalRegMap_6 ? 1'h0 : _GEN_1964; // @[decode.scala 393:{46,46}]
  wire  _GEN_2093 = 6'h3b == architecturalRegMap_6 ? 1'h0 : _GEN_1965; // @[decode.scala 393:{46,46}]
  wire  _GEN_2094 = 6'h3c == architecturalRegMap_6 ? 1'h0 : _GEN_1966; // @[decode.scala 393:{46,46}]
  wire  _GEN_2095 = 6'h3d == architecturalRegMap_6 ? 1'h0 : _GEN_1967; // @[decode.scala 393:{46,46}]
  wire  _GEN_2096 = 6'h3e == architecturalRegMap_6 ? 1'h0 : _GEN_1968; // @[decode.scala 393:{46,46}]
  wire  _GEN_2162 = 6'h0 == architecturalRegMap_7 ? 1'h0 : _GEN_2034; // @[decode.scala 393:{46,46}]
  wire  _GEN_2163 = 6'h1 == architecturalRegMap_7 ? 1'h0 : _GEN_2035; // @[decode.scala 393:{46,46}]
  wire  _GEN_2164 = 6'h2 == architecturalRegMap_7 ? 1'h0 : _GEN_2036; // @[decode.scala 393:{46,46}]
  wire  _GEN_2165 = 6'h3 == architecturalRegMap_7 ? 1'h0 : _GEN_2037; // @[decode.scala 393:{46,46}]
  wire  _GEN_2166 = 6'h4 == architecturalRegMap_7 ? 1'h0 : _GEN_2038; // @[decode.scala 393:{46,46}]
  wire  _GEN_2167 = 6'h5 == architecturalRegMap_7 ? 1'h0 : _GEN_2039; // @[decode.scala 393:{46,46}]
  wire  _GEN_2168 = 6'h6 == architecturalRegMap_7 ? 1'h0 : _GEN_2040; // @[decode.scala 393:{46,46}]
  wire  _GEN_2169 = 6'h7 == architecturalRegMap_7 ? 1'h0 : _GEN_2041; // @[decode.scala 393:{46,46}]
  wire  _GEN_2170 = 6'h8 == architecturalRegMap_7 ? 1'h0 : _GEN_2042; // @[decode.scala 393:{46,46}]
  wire  _GEN_2171 = 6'h9 == architecturalRegMap_7 ? 1'h0 : _GEN_2043; // @[decode.scala 393:{46,46}]
  wire  _GEN_2172 = 6'ha == architecturalRegMap_7 ? 1'h0 : _GEN_2044; // @[decode.scala 393:{46,46}]
  wire  _GEN_2173 = 6'hb == architecturalRegMap_7 ? 1'h0 : _GEN_2045; // @[decode.scala 393:{46,46}]
  wire  _GEN_2174 = 6'hc == architecturalRegMap_7 ? 1'h0 : _GEN_2046; // @[decode.scala 393:{46,46}]
  wire  _GEN_2175 = 6'hd == architecturalRegMap_7 ? 1'h0 : _GEN_2047; // @[decode.scala 393:{46,46}]
  wire  _GEN_2176 = 6'he == architecturalRegMap_7 ? 1'h0 : _GEN_2048; // @[decode.scala 393:{46,46}]
  wire  _GEN_2177 = 6'hf == architecturalRegMap_7 ? 1'h0 : _GEN_2049; // @[decode.scala 393:{46,46}]
  wire  _GEN_2178 = 6'h10 == architecturalRegMap_7 ? 1'h0 : _GEN_2050; // @[decode.scala 393:{46,46}]
  wire  _GEN_2179 = 6'h11 == architecturalRegMap_7 ? 1'h0 : _GEN_2051; // @[decode.scala 393:{46,46}]
  wire  _GEN_2180 = 6'h12 == architecturalRegMap_7 ? 1'h0 : _GEN_2052; // @[decode.scala 393:{46,46}]
  wire  _GEN_2181 = 6'h13 == architecturalRegMap_7 ? 1'h0 : _GEN_2053; // @[decode.scala 393:{46,46}]
  wire  _GEN_2182 = 6'h14 == architecturalRegMap_7 ? 1'h0 : _GEN_2054; // @[decode.scala 393:{46,46}]
  wire  _GEN_2183 = 6'h15 == architecturalRegMap_7 ? 1'h0 : _GEN_2055; // @[decode.scala 393:{46,46}]
  wire  _GEN_2184 = 6'h16 == architecturalRegMap_7 ? 1'h0 : _GEN_2056; // @[decode.scala 393:{46,46}]
  wire  _GEN_2185 = 6'h17 == architecturalRegMap_7 ? 1'h0 : _GEN_2057; // @[decode.scala 393:{46,46}]
  wire  _GEN_2186 = 6'h18 == architecturalRegMap_7 ? 1'h0 : _GEN_2058; // @[decode.scala 393:{46,46}]
  wire  _GEN_2187 = 6'h19 == architecturalRegMap_7 ? 1'h0 : _GEN_2059; // @[decode.scala 393:{46,46}]
  wire  _GEN_2188 = 6'h1a == architecturalRegMap_7 ? 1'h0 : _GEN_2060; // @[decode.scala 393:{46,46}]
  wire  _GEN_2189 = 6'h1b == architecturalRegMap_7 ? 1'h0 : _GEN_2061; // @[decode.scala 393:{46,46}]
  wire  _GEN_2190 = 6'h1c == architecturalRegMap_7 ? 1'h0 : _GEN_2062; // @[decode.scala 393:{46,46}]
  wire  _GEN_2191 = 6'h1d == architecturalRegMap_7 ? 1'h0 : _GEN_2063; // @[decode.scala 393:{46,46}]
  wire  _GEN_2192 = 6'h1e == architecturalRegMap_7 ? 1'h0 : _GEN_2064; // @[decode.scala 393:{46,46}]
  wire  _GEN_2193 = 6'h1f == architecturalRegMap_7 ? 1'h0 : _GEN_2065; // @[decode.scala 393:{46,46}]
  wire  _GEN_2194 = 6'h20 == architecturalRegMap_7 ? 1'h0 : _GEN_2066; // @[decode.scala 393:{46,46}]
  wire  _GEN_2195 = 6'h21 == architecturalRegMap_7 ? 1'h0 : _GEN_2067; // @[decode.scala 393:{46,46}]
  wire  _GEN_2196 = 6'h22 == architecturalRegMap_7 ? 1'h0 : _GEN_2068; // @[decode.scala 393:{46,46}]
  wire  _GEN_2197 = 6'h23 == architecturalRegMap_7 ? 1'h0 : _GEN_2069; // @[decode.scala 393:{46,46}]
  wire  _GEN_2198 = 6'h24 == architecturalRegMap_7 ? 1'h0 : _GEN_2070; // @[decode.scala 393:{46,46}]
  wire  _GEN_2199 = 6'h25 == architecturalRegMap_7 ? 1'h0 : _GEN_2071; // @[decode.scala 393:{46,46}]
  wire  _GEN_2200 = 6'h26 == architecturalRegMap_7 ? 1'h0 : _GEN_2072; // @[decode.scala 393:{46,46}]
  wire  _GEN_2201 = 6'h27 == architecturalRegMap_7 ? 1'h0 : _GEN_2073; // @[decode.scala 393:{46,46}]
  wire  _GEN_2202 = 6'h28 == architecturalRegMap_7 ? 1'h0 : _GEN_2074; // @[decode.scala 393:{46,46}]
  wire  _GEN_2203 = 6'h29 == architecturalRegMap_7 ? 1'h0 : _GEN_2075; // @[decode.scala 393:{46,46}]
  wire  _GEN_2204 = 6'h2a == architecturalRegMap_7 ? 1'h0 : _GEN_2076; // @[decode.scala 393:{46,46}]
  wire  _GEN_2205 = 6'h2b == architecturalRegMap_7 ? 1'h0 : _GEN_2077; // @[decode.scala 393:{46,46}]
  wire  _GEN_2206 = 6'h2c == architecturalRegMap_7 ? 1'h0 : _GEN_2078; // @[decode.scala 393:{46,46}]
  wire  _GEN_2207 = 6'h2d == architecturalRegMap_7 ? 1'h0 : _GEN_2079; // @[decode.scala 393:{46,46}]
  wire  _GEN_2208 = 6'h2e == architecturalRegMap_7 ? 1'h0 : _GEN_2080; // @[decode.scala 393:{46,46}]
  wire  _GEN_2209 = 6'h2f == architecturalRegMap_7 ? 1'h0 : _GEN_2081; // @[decode.scala 393:{46,46}]
  wire  _GEN_2210 = 6'h30 == architecturalRegMap_7 ? 1'h0 : _GEN_2082; // @[decode.scala 393:{46,46}]
  wire  _GEN_2211 = 6'h31 == architecturalRegMap_7 ? 1'h0 : _GEN_2083; // @[decode.scala 393:{46,46}]
  wire  _GEN_2212 = 6'h32 == architecturalRegMap_7 ? 1'h0 : _GEN_2084; // @[decode.scala 393:{46,46}]
  wire  _GEN_2213 = 6'h33 == architecturalRegMap_7 ? 1'h0 : _GEN_2085; // @[decode.scala 393:{46,46}]
  wire  _GEN_2214 = 6'h34 == architecturalRegMap_7 ? 1'h0 : _GEN_2086; // @[decode.scala 393:{46,46}]
  wire  _GEN_2215 = 6'h35 == architecturalRegMap_7 ? 1'h0 : _GEN_2087; // @[decode.scala 393:{46,46}]
  wire  _GEN_2216 = 6'h36 == architecturalRegMap_7 ? 1'h0 : _GEN_2088; // @[decode.scala 393:{46,46}]
  wire  _GEN_2217 = 6'h37 == architecturalRegMap_7 ? 1'h0 : _GEN_2089; // @[decode.scala 393:{46,46}]
  wire  _GEN_2218 = 6'h38 == architecturalRegMap_7 ? 1'h0 : _GEN_2090; // @[decode.scala 393:{46,46}]
  wire  _GEN_2219 = 6'h39 == architecturalRegMap_7 ? 1'h0 : _GEN_2091; // @[decode.scala 393:{46,46}]
  wire  _GEN_2220 = 6'h3a == architecturalRegMap_7 ? 1'h0 : _GEN_2092; // @[decode.scala 393:{46,46}]
  wire  _GEN_2221 = 6'h3b == architecturalRegMap_7 ? 1'h0 : _GEN_2093; // @[decode.scala 393:{46,46}]
  wire  _GEN_2222 = 6'h3c == architecturalRegMap_7 ? 1'h0 : _GEN_2094; // @[decode.scala 393:{46,46}]
  wire  _GEN_2223 = 6'h3d == architecturalRegMap_7 ? 1'h0 : _GEN_2095; // @[decode.scala 393:{46,46}]
  wire  _GEN_2224 = 6'h3e == architecturalRegMap_7 ? 1'h0 : _GEN_2096; // @[decode.scala 393:{46,46}]
  wire  _GEN_2290 = 6'h0 == architecturalRegMap_8 ? 1'h0 : _GEN_2162; // @[decode.scala 393:{46,46}]
  wire  _GEN_2291 = 6'h1 == architecturalRegMap_8 ? 1'h0 : _GEN_2163; // @[decode.scala 393:{46,46}]
  wire  _GEN_2292 = 6'h2 == architecturalRegMap_8 ? 1'h0 : _GEN_2164; // @[decode.scala 393:{46,46}]
  wire  _GEN_2293 = 6'h3 == architecturalRegMap_8 ? 1'h0 : _GEN_2165; // @[decode.scala 393:{46,46}]
  wire  _GEN_2294 = 6'h4 == architecturalRegMap_8 ? 1'h0 : _GEN_2166; // @[decode.scala 393:{46,46}]
  wire  _GEN_2295 = 6'h5 == architecturalRegMap_8 ? 1'h0 : _GEN_2167; // @[decode.scala 393:{46,46}]
  wire  _GEN_2296 = 6'h6 == architecturalRegMap_8 ? 1'h0 : _GEN_2168; // @[decode.scala 393:{46,46}]
  wire  _GEN_2297 = 6'h7 == architecturalRegMap_8 ? 1'h0 : _GEN_2169; // @[decode.scala 393:{46,46}]
  wire  _GEN_2298 = 6'h8 == architecturalRegMap_8 ? 1'h0 : _GEN_2170; // @[decode.scala 393:{46,46}]
  wire  _GEN_2299 = 6'h9 == architecturalRegMap_8 ? 1'h0 : _GEN_2171; // @[decode.scala 393:{46,46}]
  wire  _GEN_2300 = 6'ha == architecturalRegMap_8 ? 1'h0 : _GEN_2172; // @[decode.scala 393:{46,46}]
  wire  _GEN_2301 = 6'hb == architecturalRegMap_8 ? 1'h0 : _GEN_2173; // @[decode.scala 393:{46,46}]
  wire  _GEN_2302 = 6'hc == architecturalRegMap_8 ? 1'h0 : _GEN_2174; // @[decode.scala 393:{46,46}]
  wire  _GEN_2303 = 6'hd == architecturalRegMap_8 ? 1'h0 : _GEN_2175; // @[decode.scala 393:{46,46}]
  wire  _GEN_2304 = 6'he == architecturalRegMap_8 ? 1'h0 : _GEN_2176; // @[decode.scala 393:{46,46}]
  wire  _GEN_2305 = 6'hf == architecturalRegMap_8 ? 1'h0 : _GEN_2177; // @[decode.scala 393:{46,46}]
  wire  _GEN_2306 = 6'h10 == architecturalRegMap_8 ? 1'h0 : _GEN_2178; // @[decode.scala 393:{46,46}]
  wire  _GEN_2307 = 6'h11 == architecturalRegMap_8 ? 1'h0 : _GEN_2179; // @[decode.scala 393:{46,46}]
  wire  _GEN_2308 = 6'h12 == architecturalRegMap_8 ? 1'h0 : _GEN_2180; // @[decode.scala 393:{46,46}]
  wire  _GEN_2309 = 6'h13 == architecturalRegMap_8 ? 1'h0 : _GEN_2181; // @[decode.scala 393:{46,46}]
  wire  _GEN_2310 = 6'h14 == architecturalRegMap_8 ? 1'h0 : _GEN_2182; // @[decode.scala 393:{46,46}]
  wire  _GEN_2311 = 6'h15 == architecturalRegMap_8 ? 1'h0 : _GEN_2183; // @[decode.scala 393:{46,46}]
  wire  _GEN_2312 = 6'h16 == architecturalRegMap_8 ? 1'h0 : _GEN_2184; // @[decode.scala 393:{46,46}]
  wire  _GEN_2313 = 6'h17 == architecturalRegMap_8 ? 1'h0 : _GEN_2185; // @[decode.scala 393:{46,46}]
  wire  _GEN_2314 = 6'h18 == architecturalRegMap_8 ? 1'h0 : _GEN_2186; // @[decode.scala 393:{46,46}]
  wire  _GEN_2315 = 6'h19 == architecturalRegMap_8 ? 1'h0 : _GEN_2187; // @[decode.scala 393:{46,46}]
  wire  _GEN_2316 = 6'h1a == architecturalRegMap_8 ? 1'h0 : _GEN_2188; // @[decode.scala 393:{46,46}]
  wire  _GEN_2317 = 6'h1b == architecturalRegMap_8 ? 1'h0 : _GEN_2189; // @[decode.scala 393:{46,46}]
  wire  _GEN_2318 = 6'h1c == architecturalRegMap_8 ? 1'h0 : _GEN_2190; // @[decode.scala 393:{46,46}]
  wire  _GEN_2319 = 6'h1d == architecturalRegMap_8 ? 1'h0 : _GEN_2191; // @[decode.scala 393:{46,46}]
  wire  _GEN_2320 = 6'h1e == architecturalRegMap_8 ? 1'h0 : _GEN_2192; // @[decode.scala 393:{46,46}]
  wire  _GEN_2321 = 6'h1f == architecturalRegMap_8 ? 1'h0 : _GEN_2193; // @[decode.scala 393:{46,46}]
  wire  _GEN_2322 = 6'h20 == architecturalRegMap_8 ? 1'h0 : _GEN_2194; // @[decode.scala 393:{46,46}]
  wire  _GEN_2323 = 6'h21 == architecturalRegMap_8 ? 1'h0 : _GEN_2195; // @[decode.scala 393:{46,46}]
  wire  _GEN_2324 = 6'h22 == architecturalRegMap_8 ? 1'h0 : _GEN_2196; // @[decode.scala 393:{46,46}]
  wire  _GEN_2325 = 6'h23 == architecturalRegMap_8 ? 1'h0 : _GEN_2197; // @[decode.scala 393:{46,46}]
  wire  _GEN_2326 = 6'h24 == architecturalRegMap_8 ? 1'h0 : _GEN_2198; // @[decode.scala 393:{46,46}]
  wire  _GEN_2327 = 6'h25 == architecturalRegMap_8 ? 1'h0 : _GEN_2199; // @[decode.scala 393:{46,46}]
  wire  _GEN_2328 = 6'h26 == architecturalRegMap_8 ? 1'h0 : _GEN_2200; // @[decode.scala 393:{46,46}]
  wire  _GEN_2329 = 6'h27 == architecturalRegMap_8 ? 1'h0 : _GEN_2201; // @[decode.scala 393:{46,46}]
  wire  _GEN_2330 = 6'h28 == architecturalRegMap_8 ? 1'h0 : _GEN_2202; // @[decode.scala 393:{46,46}]
  wire  _GEN_2331 = 6'h29 == architecturalRegMap_8 ? 1'h0 : _GEN_2203; // @[decode.scala 393:{46,46}]
  wire  _GEN_2332 = 6'h2a == architecturalRegMap_8 ? 1'h0 : _GEN_2204; // @[decode.scala 393:{46,46}]
  wire  _GEN_2333 = 6'h2b == architecturalRegMap_8 ? 1'h0 : _GEN_2205; // @[decode.scala 393:{46,46}]
  wire  _GEN_2334 = 6'h2c == architecturalRegMap_8 ? 1'h0 : _GEN_2206; // @[decode.scala 393:{46,46}]
  wire  _GEN_2335 = 6'h2d == architecturalRegMap_8 ? 1'h0 : _GEN_2207; // @[decode.scala 393:{46,46}]
  wire  _GEN_2336 = 6'h2e == architecturalRegMap_8 ? 1'h0 : _GEN_2208; // @[decode.scala 393:{46,46}]
  wire  _GEN_2337 = 6'h2f == architecturalRegMap_8 ? 1'h0 : _GEN_2209; // @[decode.scala 393:{46,46}]
  wire  _GEN_2338 = 6'h30 == architecturalRegMap_8 ? 1'h0 : _GEN_2210; // @[decode.scala 393:{46,46}]
  wire  _GEN_2339 = 6'h31 == architecturalRegMap_8 ? 1'h0 : _GEN_2211; // @[decode.scala 393:{46,46}]
  wire  _GEN_2340 = 6'h32 == architecturalRegMap_8 ? 1'h0 : _GEN_2212; // @[decode.scala 393:{46,46}]
  wire  _GEN_2341 = 6'h33 == architecturalRegMap_8 ? 1'h0 : _GEN_2213; // @[decode.scala 393:{46,46}]
  wire  _GEN_2342 = 6'h34 == architecturalRegMap_8 ? 1'h0 : _GEN_2214; // @[decode.scala 393:{46,46}]
  wire  _GEN_2343 = 6'h35 == architecturalRegMap_8 ? 1'h0 : _GEN_2215; // @[decode.scala 393:{46,46}]
  wire  _GEN_2344 = 6'h36 == architecturalRegMap_8 ? 1'h0 : _GEN_2216; // @[decode.scala 393:{46,46}]
  wire  _GEN_2345 = 6'h37 == architecturalRegMap_8 ? 1'h0 : _GEN_2217; // @[decode.scala 393:{46,46}]
  wire  _GEN_2346 = 6'h38 == architecturalRegMap_8 ? 1'h0 : _GEN_2218; // @[decode.scala 393:{46,46}]
  wire  _GEN_2347 = 6'h39 == architecturalRegMap_8 ? 1'h0 : _GEN_2219; // @[decode.scala 393:{46,46}]
  wire  _GEN_2348 = 6'h3a == architecturalRegMap_8 ? 1'h0 : _GEN_2220; // @[decode.scala 393:{46,46}]
  wire  _GEN_2349 = 6'h3b == architecturalRegMap_8 ? 1'h0 : _GEN_2221; // @[decode.scala 393:{46,46}]
  wire  _GEN_2350 = 6'h3c == architecturalRegMap_8 ? 1'h0 : _GEN_2222; // @[decode.scala 393:{46,46}]
  wire  _GEN_2351 = 6'h3d == architecturalRegMap_8 ? 1'h0 : _GEN_2223; // @[decode.scala 393:{46,46}]
  wire  _GEN_2352 = 6'h3e == architecturalRegMap_8 ? 1'h0 : _GEN_2224; // @[decode.scala 393:{46,46}]
  wire  _GEN_2418 = 6'h0 == architecturalRegMap_9 ? 1'h0 : _GEN_2290; // @[decode.scala 393:{46,46}]
  wire  _GEN_2419 = 6'h1 == architecturalRegMap_9 ? 1'h0 : _GEN_2291; // @[decode.scala 393:{46,46}]
  wire  _GEN_2420 = 6'h2 == architecturalRegMap_9 ? 1'h0 : _GEN_2292; // @[decode.scala 393:{46,46}]
  wire  _GEN_2421 = 6'h3 == architecturalRegMap_9 ? 1'h0 : _GEN_2293; // @[decode.scala 393:{46,46}]
  wire  _GEN_2422 = 6'h4 == architecturalRegMap_9 ? 1'h0 : _GEN_2294; // @[decode.scala 393:{46,46}]
  wire  _GEN_2423 = 6'h5 == architecturalRegMap_9 ? 1'h0 : _GEN_2295; // @[decode.scala 393:{46,46}]
  wire  _GEN_2424 = 6'h6 == architecturalRegMap_9 ? 1'h0 : _GEN_2296; // @[decode.scala 393:{46,46}]
  wire  _GEN_2425 = 6'h7 == architecturalRegMap_9 ? 1'h0 : _GEN_2297; // @[decode.scala 393:{46,46}]
  wire  _GEN_2426 = 6'h8 == architecturalRegMap_9 ? 1'h0 : _GEN_2298; // @[decode.scala 393:{46,46}]
  wire  _GEN_2427 = 6'h9 == architecturalRegMap_9 ? 1'h0 : _GEN_2299; // @[decode.scala 393:{46,46}]
  wire  _GEN_2428 = 6'ha == architecturalRegMap_9 ? 1'h0 : _GEN_2300; // @[decode.scala 393:{46,46}]
  wire  _GEN_2429 = 6'hb == architecturalRegMap_9 ? 1'h0 : _GEN_2301; // @[decode.scala 393:{46,46}]
  wire  _GEN_2430 = 6'hc == architecturalRegMap_9 ? 1'h0 : _GEN_2302; // @[decode.scala 393:{46,46}]
  wire  _GEN_2431 = 6'hd == architecturalRegMap_9 ? 1'h0 : _GEN_2303; // @[decode.scala 393:{46,46}]
  wire  _GEN_2432 = 6'he == architecturalRegMap_9 ? 1'h0 : _GEN_2304; // @[decode.scala 393:{46,46}]
  wire  _GEN_2433 = 6'hf == architecturalRegMap_9 ? 1'h0 : _GEN_2305; // @[decode.scala 393:{46,46}]
  wire  _GEN_2434 = 6'h10 == architecturalRegMap_9 ? 1'h0 : _GEN_2306; // @[decode.scala 393:{46,46}]
  wire  _GEN_2435 = 6'h11 == architecturalRegMap_9 ? 1'h0 : _GEN_2307; // @[decode.scala 393:{46,46}]
  wire  _GEN_2436 = 6'h12 == architecturalRegMap_9 ? 1'h0 : _GEN_2308; // @[decode.scala 393:{46,46}]
  wire  _GEN_2437 = 6'h13 == architecturalRegMap_9 ? 1'h0 : _GEN_2309; // @[decode.scala 393:{46,46}]
  wire  _GEN_2438 = 6'h14 == architecturalRegMap_9 ? 1'h0 : _GEN_2310; // @[decode.scala 393:{46,46}]
  wire  _GEN_2439 = 6'h15 == architecturalRegMap_9 ? 1'h0 : _GEN_2311; // @[decode.scala 393:{46,46}]
  wire  _GEN_2440 = 6'h16 == architecturalRegMap_9 ? 1'h0 : _GEN_2312; // @[decode.scala 393:{46,46}]
  wire  _GEN_2441 = 6'h17 == architecturalRegMap_9 ? 1'h0 : _GEN_2313; // @[decode.scala 393:{46,46}]
  wire  _GEN_2442 = 6'h18 == architecturalRegMap_9 ? 1'h0 : _GEN_2314; // @[decode.scala 393:{46,46}]
  wire  _GEN_2443 = 6'h19 == architecturalRegMap_9 ? 1'h0 : _GEN_2315; // @[decode.scala 393:{46,46}]
  wire  _GEN_2444 = 6'h1a == architecturalRegMap_9 ? 1'h0 : _GEN_2316; // @[decode.scala 393:{46,46}]
  wire  _GEN_2445 = 6'h1b == architecturalRegMap_9 ? 1'h0 : _GEN_2317; // @[decode.scala 393:{46,46}]
  wire  _GEN_2446 = 6'h1c == architecturalRegMap_9 ? 1'h0 : _GEN_2318; // @[decode.scala 393:{46,46}]
  wire  _GEN_2447 = 6'h1d == architecturalRegMap_9 ? 1'h0 : _GEN_2319; // @[decode.scala 393:{46,46}]
  wire  _GEN_2448 = 6'h1e == architecturalRegMap_9 ? 1'h0 : _GEN_2320; // @[decode.scala 393:{46,46}]
  wire  _GEN_2449 = 6'h1f == architecturalRegMap_9 ? 1'h0 : _GEN_2321; // @[decode.scala 393:{46,46}]
  wire  _GEN_2450 = 6'h20 == architecturalRegMap_9 ? 1'h0 : _GEN_2322; // @[decode.scala 393:{46,46}]
  wire  _GEN_2451 = 6'h21 == architecturalRegMap_9 ? 1'h0 : _GEN_2323; // @[decode.scala 393:{46,46}]
  wire  _GEN_2452 = 6'h22 == architecturalRegMap_9 ? 1'h0 : _GEN_2324; // @[decode.scala 393:{46,46}]
  wire  _GEN_2453 = 6'h23 == architecturalRegMap_9 ? 1'h0 : _GEN_2325; // @[decode.scala 393:{46,46}]
  wire  _GEN_2454 = 6'h24 == architecturalRegMap_9 ? 1'h0 : _GEN_2326; // @[decode.scala 393:{46,46}]
  wire  _GEN_2455 = 6'h25 == architecturalRegMap_9 ? 1'h0 : _GEN_2327; // @[decode.scala 393:{46,46}]
  wire  _GEN_2456 = 6'h26 == architecturalRegMap_9 ? 1'h0 : _GEN_2328; // @[decode.scala 393:{46,46}]
  wire  _GEN_2457 = 6'h27 == architecturalRegMap_9 ? 1'h0 : _GEN_2329; // @[decode.scala 393:{46,46}]
  wire  _GEN_2458 = 6'h28 == architecturalRegMap_9 ? 1'h0 : _GEN_2330; // @[decode.scala 393:{46,46}]
  wire  _GEN_2459 = 6'h29 == architecturalRegMap_9 ? 1'h0 : _GEN_2331; // @[decode.scala 393:{46,46}]
  wire  _GEN_2460 = 6'h2a == architecturalRegMap_9 ? 1'h0 : _GEN_2332; // @[decode.scala 393:{46,46}]
  wire  _GEN_2461 = 6'h2b == architecturalRegMap_9 ? 1'h0 : _GEN_2333; // @[decode.scala 393:{46,46}]
  wire  _GEN_2462 = 6'h2c == architecturalRegMap_9 ? 1'h0 : _GEN_2334; // @[decode.scala 393:{46,46}]
  wire  _GEN_2463 = 6'h2d == architecturalRegMap_9 ? 1'h0 : _GEN_2335; // @[decode.scala 393:{46,46}]
  wire  _GEN_2464 = 6'h2e == architecturalRegMap_9 ? 1'h0 : _GEN_2336; // @[decode.scala 393:{46,46}]
  wire  _GEN_2465 = 6'h2f == architecturalRegMap_9 ? 1'h0 : _GEN_2337; // @[decode.scala 393:{46,46}]
  wire  _GEN_2466 = 6'h30 == architecturalRegMap_9 ? 1'h0 : _GEN_2338; // @[decode.scala 393:{46,46}]
  wire  _GEN_2467 = 6'h31 == architecturalRegMap_9 ? 1'h0 : _GEN_2339; // @[decode.scala 393:{46,46}]
  wire  _GEN_2468 = 6'h32 == architecturalRegMap_9 ? 1'h0 : _GEN_2340; // @[decode.scala 393:{46,46}]
  wire  _GEN_2469 = 6'h33 == architecturalRegMap_9 ? 1'h0 : _GEN_2341; // @[decode.scala 393:{46,46}]
  wire  _GEN_2470 = 6'h34 == architecturalRegMap_9 ? 1'h0 : _GEN_2342; // @[decode.scala 393:{46,46}]
  wire  _GEN_2471 = 6'h35 == architecturalRegMap_9 ? 1'h0 : _GEN_2343; // @[decode.scala 393:{46,46}]
  wire  _GEN_2472 = 6'h36 == architecturalRegMap_9 ? 1'h0 : _GEN_2344; // @[decode.scala 393:{46,46}]
  wire  _GEN_2473 = 6'h37 == architecturalRegMap_9 ? 1'h0 : _GEN_2345; // @[decode.scala 393:{46,46}]
  wire  _GEN_2474 = 6'h38 == architecturalRegMap_9 ? 1'h0 : _GEN_2346; // @[decode.scala 393:{46,46}]
  wire  _GEN_2475 = 6'h39 == architecturalRegMap_9 ? 1'h0 : _GEN_2347; // @[decode.scala 393:{46,46}]
  wire  _GEN_2476 = 6'h3a == architecturalRegMap_9 ? 1'h0 : _GEN_2348; // @[decode.scala 393:{46,46}]
  wire  _GEN_2477 = 6'h3b == architecturalRegMap_9 ? 1'h0 : _GEN_2349; // @[decode.scala 393:{46,46}]
  wire  _GEN_2478 = 6'h3c == architecturalRegMap_9 ? 1'h0 : _GEN_2350; // @[decode.scala 393:{46,46}]
  wire  _GEN_2479 = 6'h3d == architecturalRegMap_9 ? 1'h0 : _GEN_2351; // @[decode.scala 393:{46,46}]
  wire  _GEN_2480 = 6'h3e == architecturalRegMap_9 ? 1'h0 : _GEN_2352; // @[decode.scala 393:{46,46}]
  wire  _GEN_2546 = 6'h0 == architecturalRegMap_10 ? 1'h0 : _GEN_2418; // @[decode.scala 393:{46,46}]
  wire  _GEN_2547 = 6'h1 == architecturalRegMap_10 ? 1'h0 : _GEN_2419; // @[decode.scala 393:{46,46}]
  wire  _GEN_2548 = 6'h2 == architecturalRegMap_10 ? 1'h0 : _GEN_2420; // @[decode.scala 393:{46,46}]
  wire  _GEN_2549 = 6'h3 == architecturalRegMap_10 ? 1'h0 : _GEN_2421; // @[decode.scala 393:{46,46}]
  wire  _GEN_2550 = 6'h4 == architecturalRegMap_10 ? 1'h0 : _GEN_2422; // @[decode.scala 393:{46,46}]
  wire  _GEN_2551 = 6'h5 == architecturalRegMap_10 ? 1'h0 : _GEN_2423; // @[decode.scala 393:{46,46}]
  wire  _GEN_2552 = 6'h6 == architecturalRegMap_10 ? 1'h0 : _GEN_2424; // @[decode.scala 393:{46,46}]
  wire  _GEN_2553 = 6'h7 == architecturalRegMap_10 ? 1'h0 : _GEN_2425; // @[decode.scala 393:{46,46}]
  wire  _GEN_2554 = 6'h8 == architecturalRegMap_10 ? 1'h0 : _GEN_2426; // @[decode.scala 393:{46,46}]
  wire  _GEN_2555 = 6'h9 == architecturalRegMap_10 ? 1'h0 : _GEN_2427; // @[decode.scala 393:{46,46}]
  wire  _GEN_2556 = 6'ha == architecturalRegMap_10 ? 1'h0 : _GEN_2428; // @[decode.scala 393:{46,46}]
  wire  _GEN_2557 = 6'hb == architecturalRegMap_10 ? 1'h0 : _GEN_2429; // @[decode.scala 393:{46,46}]
  wire  _GEN_2558 = 6'hc == architecturalRegMap_10 ? 1'h0 : _GEN_2430; // @[decode.scala 393:{46,46}]
  wire  _GEN_2559 = 6'hd == architecturalRegMap_10 ? 1'h0 : _GEN_2431; // @[decode.scala 393:{46,46}]
  wire  _GEN_2560 = 6'he == architecturalRegMap_10 ? 1'h0 : _GEN_2432; // @[decode.scala 393:{46,46}]
  wire  _GEN_2561 = 6'hf == architecturalRegMap_10 ? 1'h0 : _GEN_2433; // @[decode.scala 393:{46,46}]
  wire  _GEN_2562 = 6'h10 == architecturalRegMap_10 ? 1'h0 : _GEN_2434; // @[decode.scala 393:{46,46}]
  wire  _GEN_2563 = 6'h11 == architecturalRegMap_10 ? 1'h0 : _GEN_2435; // @[decode.scala 393:{46,46}]
  wire  _GEN_2564 = 6'h12 == architecturalRegMap_10 ? 1'h0 : _GEN_2436; // @[decode.scala 393:{46,46}]
  wire  _GEN_2565 = 6'h13 == architecturalRegMap_10 ? 1'h0 : _GEN_2437; // @[decode.scala 393:{46,46}]
  wire  _GEN_2566 = 6'h14 == architecturalRegMap_10 ? 1'h0 : _GEN_2438; // @[decode.scala 393:{46,46}]
  wire  _GEN_2567 = 6'h15 == architecturalRegMap_10 ? 1'h0 : _GEN_2439; // @[decode.scala 393:{46,46}]
  wire  _GEN_2568 = 6'h16 == architecturalRegMap_10 ? 1'h0 : _GEN_2440; // @[decode.scala 393:{46,46}]
  wire  _GEN_2569 = 6'h17 == architecturalRegMap_10 ? 1'h0 : _GEN_2441; // @[decode.scala 393:{46,46}]
  wire  _GEN_2570 = 6'h18 == architecturalRegMap_10 ? 1'h0 : _GEN_2442; // @[decode.scala 393:{46,46}]
  wire  _GEN_2571 = 6'h19 == architecturalRegMap_10 ? 1'h0 : _GEN_2443; // @[decode.scala 393:{46,46}]
  wire  _GEN_2572 = 6'h1a == architecturalRegMap_10 ? 1'h0 : _GEN_2444; // @[decode.scala 393:{46,46}]
  wire  _GEN_2573 = 6'h1b == architecturalRegMap_10 ? 1'h0 : _GEN_2445; // @[decode.scala 393:{46,46}]
  wire  _GEN_2574 = 6'h1c == architecturalRegMap_10 ? 1'h0 : _GEN_2446; // @[decode.scala 393:{46,46}]
  wire  _GEN_2575 = 6'h1d == architecturalRegMap_10 ? 1'h0 : _GEN_2447; // @[decode.scala 393:{46,46}]
  wire  _GEN_2576 = 6'h1e == architecturalRegMap_10 ? 1'h0 : _GEN_2448; // @[decode.scala 393:{46,46}]
  wire  _GEN_2577 = 6'h1f == architecturalRegMap_10 ? 1'h0 : _GEN_2449; // @[decode.scala 393:{46,46}]
  wire  _GEN_2578 = 6'h20 == architecturalRegMap_10 ? 1'h0 : _GEN_2450; // @[decode.scala 393:{46,46}]
  wire  _GEN_2579 = 6'h21 == architecturalRegMap_10 ? 1'h0 : _GEN_2451; // @[decode.scala 393:{46,46}]
  wire  _GEN_2580 = 6'h22 == architecturalRegMap_10 ? 1'h0 : _GEN_2452; // @[decode.scala 393:{46,46}]
  wire  _GEN_2581 = 6'h23 == architecturalRegMap_10 ? 1'h0 : _GEN_2453; // @[decode.scala 393:{46,46}]
  wire  _GEN_2582 = 6'h24 == architecturalRegMap_10 ? 1'h0 : _GEN_2454; // @[decode.scala 393:{46,46}]
  wire  _GEN_2583 = 6'h25 == architecturalRegMap_10 ? 1'h0 : _GEN_2455; // @[decode.scala 393:{46,46}]
  wire  _GEN_2584 = 6'h26 == architecturalRegMap_10 ? 1'h0 : _GEN_2456; // @[decode.scala 393:{46,46}]
  wire  _GEN_2585 = 6'h27 == architecturalRegMap_10 ? 1'h0 : _GEN_2457; // @[decode.scala 393:{46,46}]
  wire  _GEN_2586 = 6'h28 == architecturalRegMap_10 ? 1'h0 : _GEN_2458; // @[decode.scala 393:{46,46}]
  wire  _GEN_2587 = 6'h29 == architecturalRegMap_10 ? 1'h0 : _GEN_2459; // @[decode.scala 393:{46,46}]
  wire  _GEN_2588 = 6'h2a == architecturalRegMap_10 ? 1'h0 : _GEN_2460; // @[decode.scala 393:{46,46}]
  wire  _GEN_2589 = 6'h2b == architecturalRegMap_10 ? 1'h0 : _GEN_2461; // @[decode.scala 393:{46,46}]
  wire  _GEN_2590 = 6'h2c == architecturalRegMap_10 ? 1'h0 : _GEN_2462; // @[decode.scala 393:{46,46}]
  wire  _GEN_2591 = 6'h2d == architecturalRegMap_10 ? 1'h0 : _GEN_2463; // @[decode.scala 393:{46,46}]
  wire  _GEN_2592 = 6'h2e == architecturalRegMap_10 ? 1'h0 : _GEN_2464; // @[decode.scala 393:{46,46}]
  wire  _GEN_2593 = 6'h2f == architecturalRegMap_10 ? 1'h0 : _GEN_2465; // @[decode.scala 393:{46,46}]
  wire  _GEN_2594 = 6'h30 == architecturalRegMap_10 ? 1'h0 : _GEN_2466; // @[decode.scala 393:{46,46}]
  wire  _GEN_2595 = 6'h31 == architecturalRegMap_10 ? 1'h0 : _GEN_2467; // @[decode.scala 393:{46,46}]
  wire  _GEN_2596 = 6'h32 == architecturalRegMap_10 ? 1'h0 : _GEN_2468; // @[decode.scala 393:{46,46}]
  wire  _GEN_2597 = 6'h33 == architecturalRegMap_10 ? 1'h0 : _GEN_2469; // @[decode.scala 393:{46,46}]
  wire  _GEN_2598 = 6'h34 == architecturalRegMap_10 ? 1'h0 : _GEN_2470; // @[decode.scala 393:{46,46}]
  wire  _GEN_2599 = 6'h35 == architecturalRegMap_10 ? 1'h0 : _GEN_2471; // @[decode.scala 393:{46,46}]
  wire  _GEN_2600 = 6'h36 == architecturalRegMap_10 ? 1'h0 : _GEN_2472; // @[decode.scala 393:{46,46}]
  wire  _GEN_2601 = 6'h37 == architecturalRegMap_10 ? 1'h0 : _GEN_2473; // @[decode.scala 393:{46,46}]
  wire  _GEN_2602 = 6'h38 == architecturalRegMap_10 ? 1'h0 : _GEN_2474; // @[decode.scala 393:{46,46}]
  wire  _GEN_2603 = 6'h39 == architecturalRegMap_10 ? 1'h0 : _GEN_2475; // @[decode.scala 393:{46,46}]
  wire  _GEN_2604 = 6'h3a == architecturalRegMap_10 ? 1'h0 : _GEN_2476; // @[decode.scala 393:{46,46}]
  wire  _GEN_2605 = 6'h3b == architecturalRegMap_10 ? 1'h0 : _GEN_2477; // @[decode.scala 393:{46,46}]
  wire  _GEN_2606 = 6'h3c == architecturalRegMap_10 ? 1'h0 : _GEN_2478; // @[decode.scala 393:{46,46}]
  wire  _GEN_2607 = 6'h3d == architecturalRegMap_10 ? 1'h0 : _GEN_2479; // @[decode.scala 393:{46,46}]
  wire  _GEN_2608 = 6'h3e == architecturalRegMap_10 ? 1'h0 : _GEN_2480; // @[decode.scala 393:{46,46}]
  wire  _GEN_2674 = 6'h0 == architecturalRegMap_11 ? 1'h0 : _GEN_2546; // @[decode.scala 393:{46,46}]
  wire  _GEN_2675 = 6'h1 == architecturalRegMap_11 ? 1'h0 : _GEN_2547; // @[decode.scala 393:{46,46}]
  wire  _GEN_2676 = 6'h2 == architecturalRegMap_11 ? 1'h0 : _GEN_2548; // @[decode.scala 393:{46,46}]
  wire  _GEN_2677 = 6'h3 == architecturalRegMap_11 ? 1'h0 : _GEN_2549; // @[decode.scala 393:{46,46}]
  wire  _GEN_2678 = 6'h4 == architecturalRegMap_11 ? 1'h0 : _GEN_2550; // @[decode.scala 393:{46,46}]
  wire  _GEN_2679 = 6'h5 == architecturalRegMap_11 ? 1'h0 : _GEN_2551; // @[decode.scala 393:{46,46}]
  wire  _GEN_2680 = 6'h6 == architecturalRegMap_11 ? 1'h0 : _GEN_2552; // @[decode.scala 393:{46,46}]
  wire  _GEN_2681 = 6'h7 == architecturalRegMap_11 ? 1'h0 : _GEN_2553; // @[decode.scala 393:{46,46}]
  wire  _GEN_2682 = 6'h8 == architecturalRegMap_11 ? 1'h0 : _GEN_2554; // @[decode.scala 393:{46,46}]
  wire  _GEN_2683 = 6'h9 == architecturalRegMap_11 ? 1'h0 : _GEN_2555; // @[decode.scala 393:{46,46}]
  wire  _GEN_2684 = 6'ha == architecturalRegMap_11 ? 1'h0 : _GEN_2556; // @[decode.scala 393:{46,46}]
  wire  _GEN_2685 = 6'hb == architecturalRegMap_11 ? 1'h0 : _GEN_2557; // @[decode.scala 393:{46,46}]
  wire  _GEN_2686 = 6'hc == architecturalRegMap_11 ? 1'h0 : _GEN_2558; // @[decode.scala 393:{46,46}]
  wire  _GEN_2687 = 6'hd == architecturalRegMap_11 ? 1'h0 : _GEN_2559; // @[decode.scala 393:{46,46}]
  wire  _GEN_2688 = 6'he == architecturalRegMap_11 ? 1'h0 : _GEN_2560; // @[decode.scala 393:{46,46}]
  wire  _GEN_2689 = 6'hf == architecturalRegMap_11 ? 1'h0 : _GEN_2561; // @[decode.scala 393:{46,46}]
  wire  _GEN_2690 = 6'h10 == architecturalRegMap_11 ? 1'h0 : _GEN_2562; // @[decode.scala 393:{46,46}]
  wire  _GEN_2691 = 6'h11 == architecturalRegMap_11 ? 1'h0 : _GEN_2563; // @[decode.scala 393:{46,46}]
  wire  _GEN_2692 = 6'h12 == architecturalRegMap_11 ? 1'h0 : _GEN_2564; // @[decode.scala 393:{46,46}]
  wire  _GEN_2693 = 6'h13 == architecturalRegMap_11 ? 1'h0 : _GEN_2565; // @[decode.scala 393:{46,46}]
  wire  _GEN_2694 = 6'h14 == architecturalRegMap_11 ? 1'h0 : _GEN_2566; // @[decode.scala 393:{46,46}]
  wire  _GEN_2695 = 6'h15 == architecturalRegMap_11 ? 1'h0 : _GEN_2567; // @[decode.scala 393:{46,46}]
  wire  _GEN_2696 = 6'h16 == architecturalRegMap_11 ? 1'h0 : _GEN_2568; // @[decode.scala 393:{46,46}]
  wire  _GEN_2697 = 6'h17 == architecturalRegMap_11 ? 1'h0 : _GEN_2569; // @[decode.scala 393:{46,46}]
  wire  _GEN_2698 = 6'h18 == architecturalRegMap_11 ? 1'h0 : _GEN_2570; // @[decode.scala 393:{46,46}]
  wire  _GEN_2699 = 6'h19 == architecturalRegMap_11 ? 1'h0 : _GEN_2571; // @[decode.scala 393:{46,46}]
  wire  _GEN_2700 = 6'h1a == architecturalRegMap_11 ? 1'h0 : _GEN_2572; // @[decode.scala 393:{46,46}]
  wire  _GEN_2701 = 6'h1b == architecturalRegMap_11 ? 1'h0 : _GEN_2573; // @[decode.scala 393:{46,46}]
  wire  _GEN_2702 = 6'h1c == architecturalRegMap_11 ? 1'h0 : _GEN_2574; // @[decode.scala 393:{46,46}]
  wire  _GEN_2703 = 6'h1d == architecturalRegMap_11 ? 1'h0 : _GEN_2575; // @[decode.scala 393:{46,46}]
  wire  _GEN_2704 = 6'h1e == architecturalRegMap_11 ? 1'h0 : _GEN_2576; // @[decode.scala 393:{46,46}]
  wire  _GEN_2705 = 6'h1f == architecturalRegMap_11 ? 1'h0 : _GEN_2577; // @[decode.scala 393:{46,46}]
  wire  _GEN_2706 = 6'h20 == architecturalRegMap_11 ? 1'h0 : _GEN_2578; // @[decode.scala 393:{46,46}]
  wire  _GEN_2707 = 6'h21 == architecturalRegMap_11 ? 1'h0 : _GEN_2579; // @[decode.scala 393:{46,46}]
  wire  _GEN_2708 = 6'h22 == architecturalRegMap_11 ? 1'h0 : _GEN_2580; // @[decode.scala 393:{46,46}]
  wire  _GEN_2709 = 6'h23 == architecturalRegMap_11 ? 1'h0 : _GEN_2581; // @[decode.scala 393:{46,46}]
  wire  _GEN_2710 = 6'h24 == architecturalRegMap_11 ? 1'h0 : _GEN_2582; // @[decode.scala 393:{46,46}]
  wire  _GEN_2711 = 6'h25 == architecturalRegMap_11 ? 1'h0 : _GEN_2583; // @[decode.scala 393:{46,46}]
  wire  _GEN_2712 = 6'h26 == architecturalRegMap_11 ? 1'h0 : _GEN_2584; // @[decode.scala 393:{46,46}]
  wire  _GEN_2713 = 6'h27 == architecturalRegMap_11 ? 1'h0 : _GEN_2585; // @[decode.scala 393:{46,46}]
  wire  _GEN_2714 = 6'h28 == architecturalRegMap_11 ? 1'h0 : _GEN_2586; // @[decode.scala 393:{46,46}]
  wire  _GEN_2715 = 6'h29 == architecturalRegMap_11 ? 1'h0 : _GEN_2587; // @[decode.scala 393:{46,46}]
  wire  _GEN_2716 = 6'h2a == architecturalRegMap_11 ? 1'h0 : _GEN_2588; // @[decode.scala 393:{46,46}]
  wire  _GEN_2717 = 6'h2b == architecturalRegMap_11 ? 1'h0 : _GEN_2589; // @[decode.scala 393:{46,46}]
  wire  _GEN_2718 = 6'h2c == architecturalRegMap_11 ? 1'h0 : _GEN_2590; // @[decode.scala 393:{46,46}]
  wire  _GEN_2719 = 6'h2d == architecturalRegMap_11 ? 1'h0 : _GEN_2591; // @[decode.scala 393:{46,46}]
  wire  _GEN_2720 = 6'h2e == architecturalRegMap_11 ? 1'h0 : _GEN_2592; // @[decode.scala 393:{46,46}]
  wire  _GEN_2721 = 6'h2f == architecturalRegMap_11 ? 1'h0 : _GEN_2593; // @[decode.scala 393:{46,46}]
  wire  _GEN_2722 = 6'h30 == architecturalRegMap_11 ? 1'h0 : _GEN_2594; // @[decode.scala 393:{46,46}]
  wire  _GEN_2723 = 6'h31 == architecturalRegMap_11 ? 1'h0 : _GEN_2595; // @[decode.scala 393:{46,46}]
  wire  _GEN_2724 = 6'h32 == architecturalRegMap_11 ? 1'h0 : _GEN_2596; // @[decode.scala 393:{46,46}]
  wire  _GEN_2725 = 6'h33 == architecturalRegMap_11 ? 1'h0 : _GEN_2597; // @[decode.scala 393:{46,46}]
  wire  _GEN_2726 = 6'h34 == architecturalRegMap_11 ? 1'h0 : _GEN_2598; // @[decode.scala 393:{46,46}]
  wire  _GEN_2727 = 6'h35 == architecturalRegMap_11 ? 1'h0 : _GEN_2599; // @[decode.scala 393:{46,46}]
  wire  _GEN_2728 = 6'h36 == architecturalRegMap_11 ? 1'h0 : _GEN_2600; // @[decode.scala 393:{46,46}]
  wire  _GEN_2729 = 6'h37 == architecturalRegMap_11 ? 1'h0 : _GEN_2601; // @[decode.scala 393:{46,46}]
  wire  _GEN_2730 = 6'h38 == architecturalRegMap_11 ? 1'h0 : _GEN_2602; // @[decode.scala 393:{46,46}]
  wire  _GEN_2731 = 6'h39 == architecturalRegMap_11 ? 1'h0 : _GEN_2603; // @[decode.scala 393:{46,46}]
  wire  _GEN_2732 = 6'h3a == architecturalRegMap_11 ? 1'h0 : _GEN_2604; // @[decode.scala 393:{46,46}]
  wire  _GEN_2733 = 6'h3b == architecturalRegMap_11 ? 1'h0 : _GEN_2605; // @[decode.scala 393:{46,46}]
  wire  _GEN_2734 = 6'h3c == architecturalRegMap_11 ? 1'h0 : _GEN_2606; // @[decode.scala 393:{46,46}]
  wire  _GEN_2735 = 6'h3d == architecturalRegMap_11 ? 1'h0 : _GEN_2607; // @[decode.scala 393:{46,46}]
  wire  _GEN_2736 = 6'h3e == architecturalRegMap_11 ? 1'h0 : _GEN_2608; // @[decode.scala 393:{46,46}]
  wire  _GEN_2802 = 6'h0 == architecturalRegMap_12 ? 1'h0 : _GEN_2674; // @[decode.scala 393:{46,46}]
  wire  _GEN_2803 = 6'h1 == architecturalRegMap_12 ? 1'h0 : _GEN_2675; // @[decode.scala 393:{46,46}]
  wire  _GEN_2804 = 6'h2 == architecturalRegMap_12 ? 1'h0 : _GEN_2676; // @[decode.scala 393:{46,46}]
  wire  _GEN_2805 = 6'h3 == architecturalRegMap_12 ? 1'h0 : _GEN_2677; // @[decode.scala 393:{46,46}]
  wire  _GEN_2806 = 6'h4 == architecturalRegMap_12 ? 1'h0 : _GEN_2678; // @[decode.scala 393:{46,46}]
  wire  _GEN_2807 = 6'h5 == architecturalRegMap_12 ? 1'h0 : _GEN_2679; // @[decode.scala 393:{46,46}]
  wire  _GEN_2808 = 6'h6 == architecturalRegMap_12 ? 1'h0 : _GEN_2680; // @[decode.scala 393:{46,46}]
  wire  _GEN_2809 = 6'h7 == architecturalRegMap_12 ? 1'h0 : _GEN_2681; // @[decode.scala 393:{46,46}]
  wire  _GEN_2810 = 6'h8 == architecturalRegMap_12 ? 1'h0 : _GEN_2682; // @[decode.scala 393:{46,46}]
  wire  _GEN_2811 = 6'h9 == architecturalRegMap_12 ? 1'h0 : _GEN_2683; // @[decode.scala 393:{46,46}]
  wire  _GEN_2812 = 6'ha == architecturalRegMap_12 ? 1'h0 : _GEN_2684; // @[decode.scala 393:{46,46}]
  wire  _GEN_2813 = 6'hb == architecturalRegMap_12 ? 1'h0 : _GEN_2685; // @[decode.scala 393:{46,46}]
  wire  _GEN_2814 = 6'hc == architecturalRegMap_12 ? 1'h0 : _GEN_2686; // @[decode.scala 393:{46,46}]
  wire  _GEN_2815 = 6'hd == architecturalRegMap_12 ? 1'h0 : _GEN_2687; // @[decode.scala 393:{46,46}]
  wire  _GEN_2816 = 6'he == architecturalRegMap_12 ? 1'h0 : _GEN_2688; // @[decode.scala 393:{46,46}]
  wire  _GEN_2817 = 6'hf == architecturalRegMap_12 ? 1'h0 : _GEN_2689; // @[decode.scala 393:{46,46}]
  wire  _GEN_2818 = 6'h10 == architecturalRegMap_12 ? 1'h0 : _GEN_2690; // @[decode.scala 393:{46,46}]
  wire  _GEN_2819 = 6'h11 == architecturalRegMap_12 ? 1'h0 : _GEN_2691; // @[decode.scala 393:{46,46}]
  wire  _GEN_2820 = 6'h12 == architecturalRegMap_12 ? 1'h0 : _GEN_2692; // @[decode.scala 393:{46,46}]
  wire  _GEN_2821 = 6'h13 == architecturalRegMap_12 ? 1'h0 : _GEN_2693; // @[decode.scala 393:{46,46}]
  wire  _GEN_2822 = 6'h14 == architecturalRegMap_12 ? 1'h0 : _GEN_2694; // @[decode.scala 393:{46,46}]
  wire  _GEN_2823 = 6'h15 == architecturalRegMap_12 ? 1'h0 : _GEN_2695; // @[decode.scala 393:{46,46}]
  wire  _GEN_2824 = 6'h16 == architecturalRegMap_12 ? 1'h0 : _GEN_2696; // @[decode.scala 393:{46,46}]
  wire  _GEN_2825 = 6'h17 == architecturalRegMap_12 ? 1'h0 : _GEN_2697; // @[decode.scala 393:{46,46}]
  wire  _GEN_2826 = 6'h18 == architecturalRegMap_12 ? 1'h0 : _GEN_2698; // @[decode.scala 393:{46,46}]
  wire  _GEN_2827 = 6'h19 == architecturalRegMap_12 ? 1'h0 : _GEN_2699; // @[decode.scala 393:{46,46}]
  wire  _GEN_2828 = 6'h1a == architecturalRegMap_12 ? 1'h0 : _GEN_2700; // @[decode.scala 393:{46,46}]
  wire  _GEN_2829 = 6'h1b == architecturalRegMap_12 ? 1'h0 : _GEN_2701; // @[decode.scala 393:{46,46}]
  wire  _GEN_2830 = 6'h1c == architecturalRegMap_12 ? 1'h0 : _GEN_2702; // @[decode.scala 393:{46,46}]
  wire  _GEN_2831 = 6'h1d == architecturalRegMap_12 ? 1'h0 : _GEN_2703; // @[decode.scala 393:{46,46}]
  wire  _GEN_2832 = 6'h1e == architecturalRegMap_12 ? 1'h0 : _GEN_2704; // @[decode.scala 393:{46,46}]
  wire  _GEN_2833 = 6'h1f == architecturalRegMap_12 ? 1'h0 : _GEN_2705; // @[decode.scala 393:{46,46}]
  wire  _GEN_2834 = 6'h20 == architecturalRegMap_12 ? 1'h0 : _GEN_2706; // @[decode.scala 393:{46,46}]
  wire  _GEN_2835 = 6'h21 == architecturalRegMap_12 ? 1'h0 : _GEN_2707; // @[decode.scala 393:{46,46}]
  wire  _GEN_2836 = 6'h22 == architecturalRegMap_12 ? 1'h0 : _GEN_2708; // @[decode.scala 393:{46,46}]
  wire  _GEN_2837 = 6'h23 == architecturalRegMap_12 ? 1'h0 : _GEN_2709; // @[decode.scala 393:{46,46}]
  wire  _GEN_2838 = 6'h24 == architecturalRegMap_12 ? 1'h0 : _GEN_2710; // @[decode.scala 393:{46,46}]
  wire  _GEN_2839 = 6'h25 == architecturalRegMap_12 ? 1'h0 : _GEN_2711; // @[decode.scala 393:{46,46}]
  wire  _GEN_2840 = 6'h26 == architecturalRegMap_12 ? 1'h0 : _GEN_2712; // @[decode.scala 393:{46,46}]
  wire  _GEN_2841 = 6'h27 == architecturalRegMap_12 ? 1'h0 : _GEN_2713; // @[decode.scala 393:{46,46}]
  wire  _GEN_2842 = 6'h28 == architecturalRegMap_12 ? 1'h0 : _GEN_2714; // @[decode.scala 393:{46,46}]
  wire  _GEN_2843 = 6'h29 == architecturalRegMap_12 ? 1'h0 : _GEN_2715; // @[decode.scala 393:{46,46}]
  wire  _GEN_2844 = 6'h2a == architecturalRegMap_12 ? 1'h0 : _GEN_2716; // @[decode.scala 393:{46,46}]
  wire  _GEN_2845 = 6'h2b == architecturalRegMap_12 ? 1'h0 : _GEN_2717; // @[decode.scala 393:{46,46}]
  wire  _GEN_2846 = 6'h2c == architecturalRegMap_12 ? 1'h0 : _GEN_2718; // @[decode.scala 393:{46,46}]
  wire  _GEN_2847 = 6'h2d == architecturalRegMap_12 ? 1'h0 : _GEN_2719; // @[decode.scala 393:{46,46}]
  wire  _GEN_2848 = 6'h2e == architecturalRegMap_12 ? 1'h0 : _GEN_2720; // @[decode.scala 393:{46,46}]
  wire  _GEN_2849 = 6'h2f == architecturalRegMap_12 ? 1'h0 : _GEN_2721; // @[decode.scala 393:{46,46}]
  wire  _GEN_2850 = 6'h30 == architecturalRegMap_12 ? 1'h0 : _GEN_2722; // @[decode.scala 393:{46,46}]
  wire  _GEN_2851 = 6'h31 == architecturalRegMap_12 ? 1'h0 : _GEN_2723; // @[decode.scala 393:{46,46}]
  wire  _GEN_2852 = 6'h32 == architecturalRegMap_12 ? 1'h0 : _GEN_2724; // @[decode.scala 393:{46,46}]
  wire  _GEN_2853 = 6'h33 == architecturalRegMap_12 ? 1'h0 : _GEN_2725; // @[decode.scala 393:{46,46}]
  wire  _GEN_2854 = 6'h34 == architecturalRegMap_12 ? 1'h0 : _GEN_2726; // @[decode.scala 393:{46,46}]
  wire  _GEN_2855 = 6'h35 == architecturalRegMap_12 ? 1'h0 : _GEN_2727; // @[decode.scala 393:{46,46}]
  wire  _GEN_2856 = 6'h36 == architecturalRegMap_12 ? 1'h0 : _GEN_2728; // @[decode.scala 393:{46,46}]
  wire  _GEN_2857 = 6'h37 == architecturalRegMap_12 ? 1'h0 : _GEN_2729; // @[decode.scala 393:{46,46}]
  wire  _GEN_2858 = 6'h38 == architecturalRegMap_12 ? 1'h0 : _GEN_2730; // @[decode.scala 393:{46,46}]
  wire  _GEN_2859 = 6'h39 == architecturalRegMap_12 ? 1'h0 : _GEN_2731; // @[decode.scala 393:{46,46}]
  wire  _GEN_2860 = 6'h3a == architecturalRegMap_12 ? 1'h0 : _GEN_2732; // @[decode.scala 393:{46,46}]
  wire  _GEN_2861 = 6'h3b == architecturalRegMap_12 ? 1'h0 : _GEN_2733; // @[decode.scala 393:{46,46}]
  wire  _GEN_2862 = 6'h3c == architecturalRegMap_12 ? 1'h0 : _GEN_2734; // @[decode.scala 393:{46,46}]
  wire  _GEN_2863 = 6'h3d == architecturalRegMap_12 ? 1'h0 : _GEN_2735; // @[decode.scala 393:{46,46}]
  wire  _GEN_2864 = 6'h3e == architecturalRegMap_12 ? 1'h0 : _GEN_2736; // @[decode.scala 393:{46,46}]
  wire  _GEN_2930 = 6'h0 == architecturalRegMap_13 ? 1'h0 : _GEN_2802; // @[decode.scala 393:{46,46}]
  wire  _GEN_2931 = 6'h1 == architecturalRegMap_13 ? 1'h0 : _GEN_2803; // @[decode.scala 393:{46,46}]
  wire  _GEN_2932 = 6'h2 == architecturalRegMap_13 ? 1'h0 : _GEN_2804; // @[decode.scala 393:{46,46}]
  wire  _GEN_2933 = 6'h3 == architecturalRegMap_13 ? 1'h0 : _GEN_2805; // @[decode.scala 393:{46,46}]
  wire  _GEN_2934 = 6'h4 == architecturalRegMap_13 ? 1'h0 : _GEN_2806; // @[decode.scala 393:{46,46}]
  wire  _GEN_2935 = 6'h5 == architecturalRegMap_13 ? 1'h0 : _GEN_2807; // @[decode.scala 393:{46,46}]
  wire  _GEN_2936 = 6'h6 == architecturalRegMap_13 ? 1'h0 : _GEN_2808; // @[decode.scala 393:{46,46}]
  wire  _GEN_2937 = 6'h7 == architecturalRegMap_13 ? 1'h0 : _GEN_2809; // @[decode.scala 393:{46,46}]
  wire  _GEN_2938 = 6'h8 == architecturalRegMap_13 ? 1'h0 : _GEN_2810; // @[decode.scala 393:{46,46}]
  wire  _GEN_2939 = 6'h9 == architecturalRegMap_13 ? 1'h0 : _GEN_2811; // @[decode.scala 393:{46,46}]
  wire  _GEN_2940 = 6'ha == architecturalRegMap_13 ? 1'h0 : _GEN_2812; // @[decode.scala 393:{46,46}]
  wire  _GEN_2941 = 6'hb == architecturalRegMap_13 ? 1'h0 : _GEN_2813; // @[decode.scala 393:{46,46}]
  wire  _GEN_2942 = 6'hc == architecturalRegMap_13 ? 1'h0 : _GEN_2814; // @[decode.scala 393:{46,46}]
  wire  _GEN_2943 = 6'hd == architecturalRegMap_13 ? 1'h0 : _GEN_2815; // @[decode.scala 393:{46,46}]
  wire  _GEN_2944 = 6'he == architecturalRegMap_13 ? 1'h0 : _GEN_2816; // @[decode.scala 393:{46,46}]
  wire  _GEN_2945 = 6'hf == architecturalRegMap_13 ? 1'h0 : _GEN_2817; // @[decode.scala 393:{46,46}]
  wire  _GEN_2946 = 6'h10 == architecturalRegMap_13 ? 1'h0 : _GEN_2818; // @[decode.scala 393:{46,46}]
  wire  _GEN_2947 = 6'h11 == architecturalRegMap_13 ? 1'h0 : _GEN_2819; // @[decode.scala 393:{46,46}]
  wire  _GEN_2948 = 6'h12 == architecturalRegMap_13 ? 1'h0 : _GEN_2820; // @[decode.scala 393:{46,46}]
  wire  _GEN_2949 = 6'h13 == architecturalRegMap_13 ? 1'h0 : _GEN_2821; // @[decode.scala 393:{46,46}]
  wire  _GEN_2950 = 6'h14 == architecturalRegMap_13 ? 1'h0 : _GEN_2822; // @[decode.scala 393:{46,46}]
  wire  _GEN_2951 = 6'h15 == architecturalRegMap_13 ? 1'h0 : _GEN_2823; // @[decode.scala 393:{46,46}]
  wire  _GEN_2952 = 6'h16 == architecturalRegMap_13 ? 1'h0 : _GEN_2824; // @[decode.scala 393:{46,46}]
  wire  _GEN_2953 = 6'h17 == architecturalRegMap_13 ? 1'h0 : _GEN_2825; // @[decode.scala 393:{46,46}]
  wire  _GEN_2954 = 6'h18 == architecturalRegMap_13 ? 1'h0 : _GEN_2826; // @[decode.scala 393:{46,46}]
  wire  _GEN_2955 = 6'h19 == architecturalRegMap_13 ? 1'h0 : _GEN_2827; // @[decode.scala 393:{46,46}]
  wire  _GEN_2956 = 6'h1a == architecturalRegMap_13 ? 1'h0 : _GEN_2828; // @[decode.scala 393:{46,46}]
  wire  _GEN_2957 = 6'h1b == architecturalRegMap_13 ? 1'h0 : _GEN_2829; // @[decode.scala 393:{46,46}]
  wire  _GEN_2958 = 6'h1c == architecturalRegMap_13 ? 1'h0 : _GEN_2830; // @[decode.scala 393:{46,46}]
  wire  _GEN_2959 = 6'h1d == architecturalRegMap_13 ? 1'h0 : _GEN_2831; // @[decode.scala 393:{46,46}]
  wire  _GEN_2960 = 6'h1e == architecturalRegMap_13 ? 1'h0 : _GEN_2832; // @[decode.scala 393:{46,46}]
  wire  _GEN_2961 = 6'h1f == architecturalRegMap_13 ? 1'h0 : _GEN_2833; // @[decode.scala 393:{46,46}]
  wire  _GEN_2962 = 6'h20 == architecturalRegMap_13 ? 1'h0 : _GEN_2834; // @[decode.scala 393:{46,46}]
  wire  _GEN_2963 = 6'h21 == architecturalRegMap_13 ? 1'h0 : _GEN_2835; // @[decode.scala 393:{46,46}]
  wire  _GEN_2964 = 6'h22 == architecturalRegMap_13 ? 1'h0 : _GEN_2836; // @[decode.scala 393:{46,46}]
  wire  _GEN_2965 = 6'h23 == architecturalRegMap_13 ? 1'h0 : _GEN_2837; // @[decode.scala 393:{46,46}]
  wire  _GEN_2966 = 6'h24 == architecturalRegMap_13 ? 1'h0 : _GEN_2838; // @[decode.scala 393:{46,46}]
  wire  _GEN_2967 = 6'h25 == architecturalRegMap_13 ? 1'h0 : _GEN_2839; // @[decode.scala 393:{46,46}]
  wire  _GEN_2968 = 6'h26 == architecturalRegMap_13 ? 1'h0 : _GEN_2840; // @[decode.scala 393:{46,46}]
  wire  _GEN_2969 = 6'h27 == architecturalRegMap_13 ? 1'h0 : _GEN_2841; // @[decode.scala 393:{46,46}]
  wire  _GEN_2970 = 6'h28 == architecturalRegMap_13 ? 1'h0 : _GEN_2842; // @[decode.scala 393:{46,46}]
  wire  _GEN_2971 = 6'h29 == architecturalRegMap_13 ? 1'h0 : _GEN_2843; // @[decode.scala 393:{46,46}]
  wire  _GEN_2972 = 6'h2a == architecturalRegMap_13 ? 1'h0 : _GEN_2844; // @[decode.scala 393:{46,46}]
  wire  _GEN_2973 = 6'h2b == architecturalRegMap_13 ? 1'h0 : _GEN_2845; // @[decode.scala 393:{46,46}]
  wire  _GEN_2974 = 6'h2c == architecturalRegMap_13 ? 1'h0 : _GEN_2846; // @[decode.scala 393:{46,46}]
  wire  _GEN_2975 = 6'h2d == architecturalRegMap_13 ? 1'h0 : _GEN_2847; // @[decode.scala 393:{46,46}]
  wire  _GEN_2976 = 6'h2e == architecturalRegMap_13 ? 1'h0 : _GEN_2848; // @[decode.scala 393:{46,46}]
  wire  _GEN_2977 = 6'h2f == architecturalRegMap_13 ? 1'h0 : _GEN_2849; // @[decode.scala 393:{46,46}]
  wire  _GEN_2978 = 6'h30 == architecturalRegMap_13 ? 1'h0 : _GEN_2850; // @[decode.scala 393:{46,46}]
  wire  _GEN_2979 = 6'h31 == architecturalRegMap_13 ? 1'h0 : _GEN_2851; // @[decode.scala 393:{46,46}]
  wire  _GEN_2980 = 6'h32 == architecturalRegMap_13 ? 1'h0 : _GEN_2852; // @[decode.scala 393:{46,46}]
  wire  _GEN_2981 = 6'h33 == architecturalRegMap_13 ? 1'h0 : _GEN_2853; // @[decode.scala 393:{46,46}]
  wire  _GEN_2982 = 6'h34 == architecturalRegMap_13 ? 1'h0 : _GEN_2854; // @[decode.scala 393:{46,46}]
  wire  _GEN_2983 = 6'h35 == architecturalRegMap_13 ? 1'h0 : _GEN_2855; // @[decode.scala 393:{46,46}]
  wire  _GEN_2984 = 6'h36 == architecturalRegMap_13 ? 1'h0 : _GEN_2856; // @[decode.scala 393:{46,46}]
  wire  _GEN_2985 = 6'h37 == architecturalRegMap_13 ? 1'h0 : _GEN_2857; // @[decode.scala 393:{46,46}]
  wire  _GEN_2986 = 6'h38 == architecturalRegMap_13 ? 1'h0 : _GEN_2858; // @[decode.scala 393:{46,46}]
  wire  _GEN_2987 = 6'h39 == architecturalRegMap_13 ? 1'h0 : _GEN_2859; // @[decode.scala 393:{46,46}]
  wire  _GEN_2988 = 6'h3a == architecturalRegMap_13 ? 1'h0 : _GEN_2860; // @[decode.scala 393:{46,46}]
  wire  _GEN_2989 = 6'h3b == architecturalRegMap_13 ? 1'h0 : _GEN_2861; // @[decode.scala 393:{46,46}]
  wire  _GEN_2990 = 6'h3c == architecturalRegMap_13 ? 1'h0 : _GEN_2862; // @[decode.scala 393:{46,46}]
  wire  _GEN_2991 = 6'h3d == architecturalRegMap_13 ? 1'h0 : _GEN_2863; // @[decode.scala 393:{46,46}]
  wire  _GEN_2992 = 6'h3e == architecturalRegMap_13 ? 1'h0 : _GEN_2864; // @[decode.scala 393:{46,46}]
  wire  _GEN_3058 = 6'h0 == architecturalRegMap_14 ? 1'h0 : _GEN_2930; // @[decode.scala 393:{46,46}]
  wire  _GEN_3059 = 6'h1 == architecturalRegMap_14 ? 1'h0 : _GEN_2931; // @[decode.scala 393:{46,46}]
  wire  _GEN_3060 = 6'h2 == architecturalRegMap_14 ? 1'h0 : _GEN_2932; // @[decode.scala 393:{46,46}]
  wire  _GEN_3061 = 6'h3 == architecturalRegMap_14 ? 1'h0 : _GEN_2933; // @[decode.scala 393:{46,46}]
  wire  _GEN_3062 = 6'h4 == architecturalRegMap_14 ? 1'h0 : _GEN_2934; // @[decode.scala 393:{46,46}]
  wire  _GEN_3063 = 6'h5 == architecturalRegMap_14 ? 1'h0 : _GEN_2935; // @[decode.scala 393:{46,46}]
  wire  _GEN_3064 = 6'h6 == architecturalRegMap_14 ? 1'h0 : _GEN_2936; // @[decode.scala 393:{46,46}]
  wire  _GEN_3065 = 6'h7 == architecturalRegMap_14 ? 1'h0 : _GEN_2937; // @[decode.scala 393:{46,46}]
  wire  _GEN_3066 = 6'h8 == architecturalRegMap_14 ? 1'h0 : _GEN_2938; // @[decode.scala 393:{46,46}]
  wire  _GEN_3067 = 6'h9 == architecturalRegMap_14 ? 1'h0 : _GEN_2939; // @[decode.scala 393:{46,46}]
  wire  _GEN_3068 = 6'ha == architecturalRegMap_14 ? 1'h0 : _GEN_2940; // @[decode.scala 393:{46,46}]
  wire  _GEN_3069 = 6'hb == architecturalRegMap_14 ? 1'h0 : _GEN_2941; // @[decode.scala 393:{46,46}]
  wire  _GEN_3070 = 6'hc == architecturalRegMap_14 ? 1'h0 : _GEN_2942; // @[decode.scala 393:{46,46}]
  wire  _GEN_3071 = 6'hd == architecturalRegMap_14 ? 1'h0 : _GEN_2943; // @[decode.scala 393:{46,46}]
  wire  _GEN_3072 = 6'he == architecturalRegMap_14 ? 1'h0 : _GEN_2944; // @[decode.scala 393:{46,46}]
  wire  _GEN_3073 = 6'hf == architecturalRegMap_14 ? 1'h0 : _GEN_2945; // @[decode.scala 393:{46,46}]
  wire  _GEN_3074 = 6'h10 == architecturalRegMap_14 ? 1'h0 : _GEN_2946; // @[decode.scala 393:{46,46}]
  wire  _GEN_3075 = 6'h11 == architecturalRegMap_14 ? 1'h0 : _GEN_2947; // @[decode.scala 393:{46,46}]
  wire  _GEN_3076 = 6'h12 == architecturalRegMap_14 ? 1'h0 : _GEN_2948; // @[decode.scala 393:{46,46}]
  wire  _GEN_3077 = 6'h13 == architecturalRegMap_14 ? 1'h0 : _GEN_2949; // @[decode.scala 393:{46,46}]
  wire  _GEN_3078 = 6'h14 == architecturalRegMap_14 ? 1'h0 : _GEN_2950; // @[decode.scala 393:{46,46}]
  wire  _GEN_3079 = 6'h15 == architecturalRegMap_14 ? 1'h0 : _GEN_2951; // @[decode.scala 393:{46,46}]
  wire  _GEN_3080 = 6'h16 == architecturalRegMap_14 ? 1'h0 : _GEN_2952; // @[decode.scala 393:{46,46}]
  wire  _GEN_3081 = 6'h17 == architecturalRegMap_14 ? 1'h0 : _GEN_2953; // @[decode.scala 393:{46,46}]
  wire  _GEN_3082 = 6'h18 == architecturalRegMap_14 ? 1'h0 : _GEN_2954; // @[decode.scala 393:{46,46}]
  wire  _GEN_3083 = 6'h19 == architecturalRegMap_14 ? 1'h0 : _GEN_2955; // @[decode.scala 393:{46,46}]
  wire  _GEN_3084 = 6'h1a == architecturalRegMap_14 ? 1'h0 : _GEN_2956; // @[decode.scala 393:{46,46}]
  wire  _GEN_3085 = 6'h1b == architecturalRegMap_14 ? 1'h0 : _GEN_2957; // @[decode.scala 393:{46,46}]
  wire  _GEN_3086 = 6'h1c == architecturalRegMap_14 ? 1'h0 : _GEN_2958; // @[decode.scala 393:{46,46}]
  wire  _GEN_3087 = 6'h1d == architecturalRegMap_14 ? 1'h0 : _GEN_2959; // @[decode.scala 393:{46,46}]
  wire  _GEN_3088 = 6'h1e == architecturalRegMap_14 ? 1'h0 : _GEN_2960; // @[decode.scala 393:{46,46}]
  wire  _GEN_3089 = 6'h1f == architecturalRegMap_14 ? 1'h0 : _GEN_2961; // @[decode.scala 393:{46,46}]
  wire  _GEN_3090 = 6'h20 == architecturalRegMap_14 ? 1'h0 : _GEN_2962; // @[decode.scala 393:{46,46}]
  wire  _GEN_3091 = 6'h21 == architecturalRegMap_14 ? 1'h0 : _GEN_2963; // @[decode.scala 393:{46,46}]
  wire  _GEN_3092 = 6'h22 == architecturalRegMap_14 ? 1'h0 : _GEN_2964; // @[decode.scala 393:{46,46}]
  wire  _GEN_3093 = 6'h23 == architecturalRegMap_14 ? 1'h0 : _GEN_2965; // @[decode.scala 393:{46,46}]
  wire  _GEN_3094 = 6'h24 == architecturalRegMap_14 ? 1'h0 : _GEN_2966; // @[decode.scala 393:{46,46}]
  wire  _GEN_3095 = 6'h25 == architecturalRegMap_14 ? 1'h0 : _GEN_2967; // @[decode.scala 393:{46,46}]
  wire  _GEN_3096 = 6'h26 == architecturalRegMap_14 ? 1'h0 : _GEN_2968; // @[decode.scala 393:{46,46}]
  wire  _GEN_3097 = 6'h27 == architecturalRegMap_14 ? 1'h0 : _GEN_2969; // @[decode.scala 393:{46,46}]
  wire  _GEN_3098 = 6'h28 == architecturalRegMap_14 ? 1'h0 : _GEN_2970; // @[decode.scala 393:{46,46}]
  wire  _GEN_3099 = 6'h29 == architecturalRegMap_14 ? 1'h0 : _GEN_2971; // @[decode.scala 393:{46,46}]
  wire  _GEN_3100 = 6'h2a == architecturalRegMap_14 ? 1'h0 : _GEN_2972; // @[decode.scala 393:{46,46}]
  wire  _GEN_3101 = 6'h2b == architecturalRegMap_14 ? 1'h0 : _GEN_2973; // @[decode.scala 393:{46,46}]
  wire  _GEN_3102 = 6'h2c == architecturalRegMap_14 ? 1'h0 : _GEN_2974; // @[decode.scala 393:{46,46}]
  wire  _GEN_3103 = 6'h2d == architecturalRegMap_14 ? 1'h0 : _GEN_2975; // @[decode.scala 393:{46,46}]
  wire  _GEN_3104 = 6'h2e == architecturalRegMap_14 ? 1'h0 : _GEN_2976; // @[decode.scala 393:{46,46}]
  wire  _GEN_3105 = 6'h2f == architecturalRegMap_14 ? 1'h0 : _GEN_2977; // @[decode.scala 393:{46,46}]
  wire  _GEN_3106 = 6'h30 == architecturalRegMap_14 ? 1'h0 : _GEN_2978; // @[decode.scala 393:{46,46}]
  wire  _GEN_3107 = 6'h31 == architecturalRegMap_14 ? 1'h0 : _GEN_2979; // @[decode.scala 393:{46,46}]
  wire  _GEN_3108 = 6'h32 == architecturalRegMap_14 ? 1'h0 : _GEN_2980; // @[decode.scala 393:{46,46}]
  wire  _GEN_3109 = 6'h33 == architecturalRegMap_14 ? 1'h0 : _GEN_2981; // @[decode.scala 393:{46,46}]
  wire  _GEN_3110 = 6'h34 == architecturalRegMap_14 ? 1'h0 : _GEN_2982; // @[decode.scala 393:{46,46}]
  wire  _GEN_3111 = 6'h35 == architecturalRegMap_14 ? 1'h0 : _GEN_2983; // @[decode.scala 393:{46,46}]
  wire  _GEN_3112 = 6'h36 == architecturalRegMap_14 ? 1'h0 : _GEN_2984; // @[decode.scala 393:{46,46}]
  wire  _GEN_3113 = 6'h37 == architecturalRegMap_14 ? 1'h0 : _GEN_2985; // @[decode.scala 393:{46,46}]
  wire  _GEN_3114 = 6'h38 == architecturalRegMap_14 ? 1'h0 : _GEN_2986; // @[decode.scala 393:{46,46}]
  wire  _GEN_3115 = 6'h39 == architecturalRegMap_14 ? 1'h0 : _GEN_2987; // @[decode.scala 393:{46,46}]
  wire  _GEN_3116 = 6'h3a == architecturalRegMap_14 ? 1'h0 : _GEN_2988; // @[decode.scala 393:{46,46}]
  wire  _GEN_3117 = 6'h3b == architecturalRegMap_14 ? 1'h0 : _GEN_2989; // @[decode.scala 393:{46,46}]
  wire  _GEN_3118 = 6'h3c == architecturalRegMap_14 ? 1'h0 : _GEN_2990; // @[decode.scala 393:{46,46}]
  wire  _GEN_3119 = 6'h3d == architecturalRegMap_14 ? 1'h0 : _GEN_2991; // @[decode.scala 393:{46,46}]
  wire  _GEN_3120 = 6'h3e == architecturalRegMap_14 ? 1'h0 : _GEN_2992; // @[decode.scala 393:{46,46}]
  wire  _GEN_3122 = 6'h0 == architecturalRegMap_15 | (6'h0 == architecturalRegMap_14 | (6'h0 == architecturalRegMap_13
     | (6'h0 == architecturalRegMap_12 | (6'h0 == architecturalRegMap_11 | (6'h0 == architecturalRegMap_10 | (6'h0 ==
    architecturalRegMap_9 | (6'h0 == architecturalRegMap_8 | (6'h0 == architecturalRegMap_7 | (6'h0 ==
    architecturalRegMap_6 | (6'h0 == architecturalRegMap_5 | (6'h0 == architecturalRegMap_4 | (6'h0 ==
    architecturalRegMap_3 | (6'h0 == architecturalRegMap_2 | (6'h0 == architecturalRegMap_1 | _GEN_1202)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3123 = 6'h1 == architecturalRegMap_15 | (6'h1 == architecturalRegMap_14 | (6'h1 == architecturalRegMap_13
     | (6'h1 == architecturalRegMap_12 | (6'h1 == architecturalRegMap_11 | (6'h1 == architecturalRegMap_10 | (6'h1 ==
    architecturalRegMap_9 | (6'h1 == architecturalRegMap_8 | (6'h1 == architecturalRegMap_7 | (6'h1 ==
    architecturalRegMap_6 | (6'h1 == architecturalRegMap_5 | (6'h1 == architecturalRegMap_4 | (6'h1 ==
    architecturalRegMap_3 | (6'h1 == architecturalRegMap_2 | (6'h1 == architecturalRegMap_1 | _GEN_1203)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3124 = 6'h2 == architecturalRegMap_15 | (6'h2 == architecturalRegMap_14 | (6'h2 == architecturalRegMap_13
     | (6'h2 == architecturalRegMap_12 | (6'h2 == architecturalRegMap_11 | (6'h2 == architecturalRegMap_10 | (6'h2 ==
    architecturalRegMap_9 | (6'h2 == architecturalRegMap_8 | (6'h2 == architecturalRegMap_7 | (6'h2 ==
    architecturalRegMap_6 | (6'h2 == architecturalRegMap_5 | (6'h2 == architecturalRegMap_4 | (6'h2 ==
    architecturalRegMap_3 | (6'h2 == architecturalRegMap_2 | (6'h2 == architecturalRegMap_1 | _GEN_1204)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3125 = 6'h3 == architecturalRegMap_15 | (6'h3 == architecturalRegMap_14 | (6'h3 == architecturalRegMap_13
     | (6'h3 == architecturalRegMap_12 | (6'h3 == architecturalRegMap_11 | (6'h3 == architecturalRegMap_10 | (6'h3 ==
    architecturalRegMap_9 | (6'h3 == architecturalRegMap_8 | (6'h3 == architecturalRegMap_7 | (6'h3 ==
    architecturalRegMap_6 | (6'h3 == architecturalRegMap_5 | (6'h3 == architecturalRegMap_4 | (6'h3 ==
    architecturalRegMap_3 | (6'h3 == architecturalRegMap_2 | (6'h3 == architecturalRegMap_1 | _GEN_1205)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3126 = 6'h4 == architecturalRegMap_15 | (6'h4 == architecturalRegMap_14 | (6'h4 == architecturalRegMap_13
     | (6'h4 == architecturalRegMap_12 | (6'h4 == architecturalRegMap_11 | (6'h4 == architecturalRegMap_10 | (6'h4 ==
    architecturalRegMap_9 | (6'h4 == architecturalRegMap_8 | (6'h4 == architecturalRegMap_7 | (6'h4 ==
    architecturalRegMap_6 | (6'h4 == architecturalRegMap_5 | (6'h4 == architecturalRegMap_4 | (6'h4 ==
    architecturalRegMap_3 | (6'h4 == architecturalRegMap_2 | (6'h4 == architecturalRegMap_1 | _GEN_1206)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3127 = 6'h5 == architecturalRegMap_15 | (6'h5 == architecturalRegMap_14 | (6'h5 == architecturalRegMap_13
     | (6'h5 == architecturalRegMap_12 | (6'h5 == architecturalRegMap_11 | (6'h5 == architecturalRegMap_10 | (6'h5 ==
    architecturalRegMap_9 | (6'h5 == architecturalRegMap_8 | (6'h5 == architecturalRegMap_7 | (6'h5 ==
    architecturalRegMap_6 | (6'h5 == architecturalRegMap_5 | (6'h5 == architecturalRegMap_4 | (6'h5 ==
    architecturalRegMap_3 | (6'h5 == architecturalRegMap_2 | (6'h5 == architecturalRegMap_1 | _GEN_1207)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3128 = 6'h6 == architecturalRegMap_15 | (6'h6 == architecturalRegMap_14 | (6'h6 == architecturalRegMap_13
     | (6'h6 == architecturalRegMap_12 | (6'h6 == architecturalRegMap_11 | (6'h6 == architecturalRegMap_10 | (6'h6 ==
    architecturalRegMap_9 | (6'h6 == architecturalRegMap_8 | (6'h6 == architecturalRegMap_7 | (6'h6 ==
    architecturalRegMap_6 | (6'h6 == architecturalRegMap_5 | (6'h6 == architecturalRegMap_4 | (6'h6 ==
    architecturalRegMap_3 | (6'h6 == architecturalRegMap_2 | (6'h6 == architecturalRegMap_1 | _GEN_1208)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3129 = 6'h7 == architecturalRegMap_15 | (6'h7 == architecturalRegMap_14 | (6'h7 == architecturalRegMap_13
     | (6'h7 == architecturalRegMap_12 | (6'h7 == architecturalRegMap_11 | (6'h7 == architecturalRegMap_10 | (6'h7 ==
    architecturalRegMap_9 | (6'h7 == architecturalRegMap_8 | (6'h7 == architecturalRegMap_7 | (6'h7 ==
    architecturalRegMap_6 | (6'h7 == architecturalRegMap_5 | (6'h7 == architecturalRegMap_4 | (6'h7 ==
    architecturalRegMap_3 | (6'h7 == architecturalRegMap_2 | (6'h7 == architecturalRegMap_1 | _GEN_1209)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3130 = 6'h8 == architecturalRegMap_15 | (6'h8 == architecturalRegMap_14 | (6'h8 == architecturalRegMap_13
     | (6'h8 == architecturalRegMap_12 | (6'h8 == architecturalRegMap_11 | (6'h8 == architecturalRegMap_10 | (6'h8 ==
    architecturalRegMap_9 | (6'h8 == architecturalRegMap_8 | (6'h8 == architecturalRegMap_7 | (6'h8 ==
    architecturalRegMap_6 | (6'h8 == architecturalRegMap_5 | (6'h8 == architecturalRegMap_4 | (6'h8 ==
    architecturalRegMap_3 | (6'h8 == architecturalRegMap_2 | (6'h8 == architecturalRegMap_1 | _GEN_1210)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3131 = 6'h9 == architecturalRegMap_15 | (6'h9 == architecturalRegMap_14 | (6'h9 == architecturalRegMap_13
     | (6'h9 == architecturalRegMap_12 | (6'h9 == architecturalRegMap_11 | (6'h9 == architecturalRegMap_10 | (6'h9 ==
    architecturalRegMap_9 | (6'h9 == architecturalRegMap_8 | (6'h9 == architecturalRegMap_7 | (6'h9 ==
    architecturalRegMap_6 | (6'h9 == architecturalRegMap_5 | (6'h9 == architecturalRegMap_4 | (6'h9 ==
    architecturalRegMap_3 | (6'h9 == architecturalRegMap_2 | (6'h9 == architecturalRegMap_1 | _GEN_1211)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3132 = 6'ha == architecturalRegMap_15 | (6'ha == architecturalRegMap_14 | (6'ha == architecturalRegMap_13
     | (6'ha == architecturalRegMap_12 | (6'ha == architecturalRegMap_11 | (6'ha == architecturalRegMap_10 | (6'ha ==
    architecturalRegMap_9 | (6'ha == architecturalRegMap_8 | (6'ha == architecturalRegMap_7 | (6'ha ==
    architecturalRegMap_6 | (6'ha == architecturalRegMap_5 | (6'ha == architecturalRegMap_4 | (6'ha ==
    architecturalRegMap_3 | (6'ha == architecturalRegMap_2 | (6'ha == architecturalRegMap_1 | _GEN_1212)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3133 = 6'hb == architecturalRegMap_15 | (6'hb == architecturalRegMap_14 | (6'hb == architecturalRegMap_13
     | (6'hb == architecturalRegMap_12 | (6'hb == architecturalRegMap_11 | (6'hb == architecturalRegMap_10 | (6'hb ==
    architecturalRegMap_9 | (6'hb == architecturalRegMap_8 | (6'hb == architecturalRegMap_7 | (6'hb ==
    architecturalRegMap_6 | (6'hb == architecturalRegMap_5 | (6'hb == architecturalRegMap_4 | (6'hb ==
    architecturalRegMap_3 | (6'hb == architecturalRegMap_2 | (6'hb == architecturalRegMap_1 | _GEN_1213)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3134 = 6'hc == architecturalRegMap_15 | (6'hc == architecturalRegMap_14 | (6'hc == architecturalRegMap_13
     | (6'hc == architecturalRegMap_12 | (6'hc == architecturalRegMap_11 | (6'hc == architecturalRegMap_10 | (6'hc ==
    architecturalRegMap_9 | (6'hc == architecturalRegMap_8 | (6'hc == architecturalRegMap_7 | (6'hc ==
    architecturalRegMap_6 | (6'hc == architecturalRegMap_5 | (6'hc == architecturalRegMap_4 | (6'hc ==
    architecturalRegMap_3 | (6'hc == architecturalRegMap_2 | (6'hc == architecturalRegMap_1 | _GEN_1214)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3135 = 6'hd == architecturalRegMap_15 | (6'hd == architecturalRegMap_14 | (6'hd == architecturalRegMap_13
     | (6'hd == architecturalRegMap_12 | (6'hd == architecturalRegMap_11 | (6'hd == architecturalRegMap_10 | (6'hd ==
    architecturalRegMap_9 | (6'hd == architecturalRegMap_8 | (6'hd == architecturalRegMap_7 | (6'hd ==
    architecturalRegMap_6 | (6'hd == architecturalRegMap_5 | (6'hd == architecturalRegMap_4 | (6'hd ==
    architecturalRegMap_3 | (6'hd == architecturalRegMap_2 | (6'hd == architecturalRegMap_1 | _GEN_1215)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3136 = 6'he == architecturalRegMap_15 | (6'he == architecturalRegMap_14 | (6'he == architecturalRegMap_13
     | (6'he == architecturalRegMap_12 | (6'he == architecturalRegMap_11 | (6'he == architecturalRegMap_10 | (6'he ==
    architecturalRegMap_9 | (6'he == architecturalRegMap_8 | (6'he == architecturalRegMap_7 | (6'he ==
    architecturalRegMap_6 | (6'he == architecturalRegMap_5 | (6'he == architecturalRegMap_4 | (6'he ==
    architecturalRegMap_3 | (6'he == architecturalRegMap_2 | (6'he == architecturalRegMap_1 | _GEN_1216)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3137 = 6'hf == architecturalRegMap_15 | (6'hf == architecturalRegMap_14 | (6'hf == architecturalRegMap_13
     | (6'hf == architecturalRegMap_12 | (6'hf == architecturalRegMap_11 | (6'hf == architecturalRegMap_10 | (6'hf ==
    architecturalRegMap_9 | (6'hf == architecturalRegMap_8 | (6'hf == architecturalRegMap_7 | (6'hf ==
    architecturalRegMap_6 | (6'hf == architecturalRegMap_5 | (6'hf == architecturalRegMap_4 | (6'hf ==
    architecturalRegMap_3 | (6'hf == architecturalRegMap_2 | (6'hf == architecturalRegMap_1 | _GEN_1217)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3138 = 6'h10 == architecturalRegMap_15 | (6'h10 == architecturalRegMap_14 | (6'h10 ==
    architecturalRegMap_13 | (6'h10 == architecturalRegMap_12 | (6'h10 == architecturalRegMap_11 | (6'h10 ==
    architecturalRegMap_10 | (6'h10 == architecturalRegMap_9 | (6'h10 == architecturalRegMap_8 | (6'h10 ==
    architecturalRegMap_7 | (6'h10 == architecturalRegMap_6 | (6'h10 == architecturalRegMap_5 | (6'h10 ==
    architecturalRegMap_4 | (6'h10 == architecturalRegMap_3 | (6'h10 == architecturalRegMap_2 | (6'h10 ==
    architecturalRegMap_1 | _GEN_1218)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3139 = 6'h11 == architecturalRegMap_15 | (6'h11 == architecturalRegMap_14 | (6'h11 ==
    architecturalRegMap_13 | (6'h11 == architecturalRegMap_12 | (6'h11 == architecturalRegMap_11 | (6'h11 ==
    architecturalRegMap_10 | (6'h11 == architecturalRegMap_9 | (6'h11 == architecturalRegMap_8 | (6'h11 ==
    architecturalRegMap_7 | (6'h11 == architecturalRegMap_6 | (6'h11 == architecturalRegMap_5 | (6'h11 ==
    architecturalRegMap_4 | (6'h11 == architecturalRegMap_3 | (6'h11 == architecturalRegMap_2 | (6'h11 ==
    architecturalRegMap_1 | _GEN_1219)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3140 = 6'h12 == architecturalRegMap_15 | (6'h12 == architecturalRegMap_14 | (6'h12 ==
    architecturalRegMap_13 | (6'h12 == architecturalRegMap_12 | (6'h12 == architecturalRegMap_11 | (6'h12 ==
    architecturalRegMap_10 | (6'h12 == architecturalRegMap_9 | (6'h12 == architecturalRegMap_8 | (6'h12 ==
    architecturalRegMap_7 | (6'h12 == architecturalRegMap_6 | (6'h12 == architecturalRegMap_5 | (6'h12 ==
    architecturalRegMap_4 | (6'h12 == architecturalRegMap_3 | (6'h12 == architecturalRegMap_2 | (6'h12 ==
    architecturalRegMap_1 | _GEN_1220)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3141 = 6'h13 == architecturalRegMap_15 | (6'h13 == architecturalRegMap_14 | (6'h13 ==
    architecturalRegMap_13 | (6'h13 == architecturalRegMap_12 | (6'h13 == architecturalRegMap_11 | (6'h13 ==
    architecturalRegMap_10 | (6'h13 == architecturalRegMap_9 | (6'h13 == architecturalRegMap_8 | (6'h13 ==
    architecturalRegMap_7 | (6'h13 == architecturalRegMap_6 | (6'h13 == architecturalRegMap_5 | (6'h13 ==
    architecturalRegMap_4 | (6'h13 == architecturalRegMap_3 | (6'h13 == architecturalRegMap_2 | (6'h13 ==
    architecturalRegMap_1 | _GEN_1221)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3142 = 6'h14 == architecturalRegMap_15 | (6'h14 == architecturalRegMap_14 | (6'h14 ==
    architecturalRegMap_13 | (6'h14 == architecturalRegMap_12 | (6'h14 == architecturalRegMap_11 | (6'h14 ==
    architecturalRegMap_10 | (6'h14 == architecturalRegMap_9 | (6'h14 == architecturalRegMap_8 | (6'h14 ==
    architecturalRegMap_7 | (6'h14 == architecturalRegMap_6 | (6'h14 == architecturalRegMap_5 | (6'h14 ==
    architecturalRegMap_4 | (6'h14 == architecturalRegMap_3 | (6'h14 == architecturalRegMap_2 | (6'h14 ==
    architecturalRegMap_1 | _GEN_1222)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3143 = 6'h15 == architecturalRegMap_15 | (6'h15 == architecturalRegMap_14 | (6'h15 ==
    architecturalRegMap_13 | (6'h15 == architecturalRegMap_12 | (6'h15 == architecturalRegMap_11 | (6'h15 ==
    architecturalRegMap_10 | (6'h15 == architecturalRegMap_9 | (6'h15 == architecturalRegMap_8 | (6'h15 ==
    architecturalRegMap_7 | (6'h15 == architecturalRegMap_6 | (6'h15 == architecturalRegMap_5 | (6'h15 ==
    architecturalRegMap_4 | (6'h15 == architecturalRegMap_3 | (6'h15 == architecturalRegMap_2 | (6'h15 ==
    architecturalRegMap_1 | _GEN_1223)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3144 = 6'h16 == architecturalRegMap_15 | (6'h16 == architecturalRegMap_14 | (6'h16 ==
    architecturalRegMap_13 | (6'h16 == architecturalRegMap_12 | (6'h16 == architecturalRegMap_11 | (6'h16 ==
    architecturalRegMap_10 | (6'h16 == architecturalRegMap_9 | (6'h16 == architecturalRegMap_8 | (6'h16 ==
    architecturalRegMap_7 | (6'h16 == architecturalRegMap_6 | (6'h16 == architecturalRegMap_5 | (6'h16 ==
    architecturalRegMap_4 | (6'h16 == architecturalRegMap_3 | (6'h16 == architecturalRegMap_2 | (6'h16 ==
    architecturalRegMap_1 | _GEN_1224)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3145 = 6'h17 == architecturalRegMap_15 | (6'h17 == architecturalRegMap_14 | (6'h17 ==
    architecturalRegMap_13 | (6'h17 == architecturalRegMap_12 | (6'h17 == architecturalRegMap_11 | (6'h17 ==
    architecturalRegMap_10 | (6'h17 == architecturalRegMap_9 | (6'h17 == architecturalRegMap_8 | (6'h17 ==
    architecturalRegMap_7 | (6'h17 == architecturalRegMap_6 | (6'h17 == architecturalRegMap_5 | (6'h17 ==
    architecturalRegMap_4 | (6'h17 == architecturalRegMap_3 | (6'h17 == architecturalRegMap_2 | (6'h17 ==
    architecturalRegMap_1 | _GEN_1225)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3146 = 6'h18 == architecturalRegMap_15 | (6'h18 == architecturalRegMap_14 | (6'h18 ==
    architecturalRegMap_13 | (6'h18 == architecturalRegMap_12 | (6'h18 == architecturalRegMap_11 | (6'h18 ==
    architecturalRegMap_10 | (6'h18 == architecturalRegMap_9 | (6'h18 == architecturalRegMap_8 | (6'h18 ==
    architecturalRegMap_7 | (6'h18 == architecturalRegMap_6 | (6'h18 == architecturalRegMap_5 | (6'h18 ==
    architecturalRegMap_4 | (6'h18 == architecturalRegMap_3 | (6'h18 == architecturalRegMap_2 | (6'h18 ==
    architecturalRegMap_1 | _GEN_1226)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3147 = 6'h19 == architecturalRegMap_15 | (6'h19 == architecturalRegMap_14 | (6'h19 ==
    architecturalRegMap_13 | (6'h19 == architecturalRegMap_12 | (6'h19 == architecturalRegMap_11 | (6'h19 ==
    architecturalRegMap_10 | (6'h19 == architecturalRegMap_9 | (6'h19 == architecturalRegMap_8 | (6'h19 ==
    architecturalRegMap_7 | (6'h19 == architecturalRegMap_6 | (6'h19 == architecturalRegMap_5 | (6'h19 ==
    architecturalRegMap_4 | (6'h19 == architecturalRegMap_3 | (6'h19 == architecturalRegMap_2 | (6'h19 ==
    architecturalRegMap_1 | _GEN_1227)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3148 = 6'h1a == architecturalRegMap_15 | (6'h1a == architecturalRegMap_14 | (6'h1a ==
    architecturalRegMap_13 | (6'h1a == architecturalRegMap_12 | (6'h1a == architecturalRegMap_11 | (6'h1a ==
    architecturalRegMap_10 | (6'h1a == architecturalRegMap_9 | (6'h1a == architecturalRegMap_8 | (6'h1a ==
    architecturalRegMap_7 | (6'h1a == architecturalRegMap_6 | (6'h1a == architecturalRegMap_5 | (6'h1a ==
    architecturalRegMap_4 | (6'h1a == architecturalRegMap_3 | (6'h1a == architecturalRegMap_2 | (6'h1a ==
    architecturalRegMap_1 | _GEN_1228)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3149 = 6'h1b == architecturalRegMap_15 | (6'h1b == architecturalRegMap_14 | (6'h1b ==
    architecturalRegMap_13 | (6'h1b == architecturalRegMap_12 | (6'h1b == architecturalRegMap_11 | (6'h1b ==
    architecturalRegMap_10 | (6'h1b == architecturalRegMap_9 | (6'h1b == architecturalRegMap_8 | (6'h1b ==
    architecturalRegMap_7 | (6'h1b == architecturalRegMap_6 | (6'h1b == architecturalRegMap_5 | (6'h1b ==
    architecturalRegMap_4 | (6'h1b == architecturalRegMap_3 | (6'h1b == architecturalRegMap_2 | (6'h1b ==
    architecturalRegMap_1 | _GEN_1229)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3150 = 6'h1c == architecturalRegMap_15 | (6'h1c == architecturalRegMap_14 | (6'h1c ==
    architecturalRegMap_13 | (6'h1c == architecturalRegMap_12 | (6'h1c == architecturalRegMap_11 | (6'h1c ==
    architecturalRegMap_10 | (6'h1c == architecturalRegMap_9 | (6'h1c == architecturalRegMap_8 | (6'h1c ==
    architecturalRegMap_7 | (6'h1c == architecturalRegMap_6 | (6'h1c == architecturalRegMap_5 | (6'h1c ==
    architecturalRegMap_4 | (6'h1c == architecturalRegMap_3 | (6'h1c == architecturalRegMap_2 | (6'h1c ==
    architecturalRegMap_1 | _GEN_1230)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3151 = 6'h1d == architecturalRegMap_15 | (6'h1d == architecturalRegMap_14 | (6'h1d ==
    architecturalRegMap_13 | (6'h1d == architecturalRegMap_12 | (6'h1d == architecturalRegMap_11 | (6'h1d ==
    architecturalRegMap_10 | (6'h1d == architecturalRegMap_9 | (6'h1d == architecturalRegMap_8 | (6'h1d ==
    architecturalRegMap_7 | (6'h1d == architecturalRegMap_6 | (6'h1d == architecturalRegMap_5 | (6'h1d ==
    architecturalRegMap_4 | (6'h1d == architecturalRegMap_3 | (6'h1d == architecturalRegMap_2 | (6'h1d ==
    architecturalRegMap_1 | _GEN_1231)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3152 = 6'h1e == architecturalRegMap_15 | (6'h1e == architecturalRegMap_14 | (6'h1e ==
    architecturalRegMap_13 | (6'h1e == architecturalRegMap_12 | (6'h1e == architecturalRegMap_11 | (6'h1e ==
    architecturalRegMap_10 | (6'h1e == architecturalRegMap_9 | (6'h1e == architecturalRegMap_8 | (6'h1e ==
    architecturalRegMap_7 | (6'h1e == architecturalRegMap_6 | (6'h1e == architecturalRegMap_5 | (6'h1e ==
    architecturalRegMap_4 | (6'h1e == architecturalRegMap_3 | (6'h1e == architecturalRegMap_2 | (6'h1e ==
    architecturalRegMap_1 | _GEN_1232)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3153 = 6'h1f == architecturalRegMap_15 | (6'h1f == architecturalRegMap_14 | (6'h1f ==
    architecturalRegMap_13 | (6'h1f == architecturalRegMap_12 | (6'h1f == architecturalRegMap_11 | (6'h1f ==
    architecturalRegMap_10 | (6'h1f == architecturalRegMap_9 | (6'h1f == architecturalRegMap_8 | (6'h1f ==
    architecturalRegMap_7 | (6'h1f == architecturalRegMap_6 | (6'h1f == architecturalRegMap_5 | (6'h1f ==
    architecturalRegMap_4 | (6'h1f == architecturalRegMap_3 | (6'h1f == architecturalRegMap_2 | (6'h1f ==
    architecturalRegMap_1 | _GEN_1233)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3154 = 6'h20 == architecturalRegMap_15 | (6'h20 == architecturalRegMap_14 | (6'h20 ==
    architecturalRegMap_13 | (6'h20 == architecturalRegMap_12 | (6'h20 == architecturalRegMap_11 | (6'h20 ==
    architecturalRegMap_10 | (6'h20 == architecturalRegMap_9 | (6'h20 == architecturalRegMap_8 | (6'h20 ==
    architecturalRegMap_7 | (6'h20 == architecturalRegMap_6 | (6'h20 == architecturalRegMap_5 | (6'h20 ==
    architecturalRegMap_4 | (6'h20 == architecturalRegMap_3 | (6'h20 == architecturalRegMap_2 | (6'h20 ==
    architecturalRegMap_1 | _GEN_1234)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3155 = 6'h21 == architecturalRegMap_15 | (6'h21 == architecturalRegMap_14 | (6'h21 ==
    architecturalRegMap_13 | (6'h21 == architecturalRegMap_12 | (6'h21 == architecturalRegMap_11 | (6'h21 ==
    architecturalRegMap_10 | (6'h21 == architecturalRegMap_9 | (6'h21 == architecturalRegMap_8 | (6'h21 ==
    architecturalRegMap_7 | (6'h21 == architecturalRegMap_6 | (6'h21 == architecturalRegMap_5 | (6'h21 ==
    architecturalRegMap_4 | (6'h21 == architecturalRegMap_3 | (6'h21 == architecturalRegMap_2 | (6'h21 ==
    architecturalRegMap_1 | _GEN_1235)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3156 = 6'h22 == architecturalRegMap_15 | (6'h22 == architecturalRegMap_14 | (6'h22 ==
    architecturalRegMap_13 | (6'h22 == architecturalRegMap_12 | (6'h22 == architecturalRegMap_11 | (6'h22 ==
    architecturalRegMap_10 | (6'h22 == architecturalRegMap_9 | (6'h22 == architecturalRegMap_8 | (6'h22 ==
    architecturalRegMap_7 | (6'h22 == architecturalRegMap_6 | (6'h22 == architecturalRegMap_5 | (6'h22 ==
    architecturalRegMap_4 | (6'h22 == architecturalRegMap_3 | (6'h22 == architecturalRegMap_2 | (6'h22 ==
    architecturalRegMap_1 | _GEN_1236)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3157 = 6'h23 == architecturalRegMap_15 | (6'h23 == architecturalRegMap_14 | (6'h23 ==
    architecturalRegMap_13 | (6'h23 == architecturalRegMap_12 | (6'h23 == architecturalRegMap_11 | (6'h23 ==
    architecturalRegMap_10 | (6'h23 == architecturalRegMap_9 | (6'h23 == architecturalRegMap_8 | (6'h23 ==
    architecturalRegMap_7 | (6'h23 == architecturalRegMap_6 | (6'h23 == architecturalRegMap_5 | (6'h23 ==
    architecturalRegMap_4 | (6'h23 == architecturalRegMap_3 | (6'h23 == architecturalRegMap_2 | (6'h23 ==
    architecturalRegMap_1 | _GEN_1237)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3158 = 6'h24 == architecturalRegMap_15 | (6'h24 == architecturalRegMap_14 | (6'h24 ==
    architecturalRegMap_13 | (6'h24 == architecturalRegMap_12 | (6'h24 == architecturalRegMap_11 | (6'h24 ==
    architecturalRegMap_10 | (6'h24 == architecturalRegMap_9 | (6'h24 == architecturalRegMap_8 | (6'h24 ==
    architecturalRegMap_7 | (6'h24 == architecturalRegMap_6 | (6'h24 == architecturalRegMap_5 | (6'h24 ==
    architecturalRegMap_4 | (6'h24 == architecturalRegMap_3 | (6'h24 == architecturalRegMap_2 | (6'h24 ==
    architecturalRegMap_1 | _GEN_1238)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3159 = 6'h25 == architecturalRegMap_15 | (6'h25 == architecturalRegMap_14 | (6'h25 ==
    architecturalRegMap_13 | (6'h25 == architecturalRegMap_12 | (6'h25 == architecturalRegMap_11 | (6'h25 ==
    architecturalRegMap_10 | (6'h25 == architecturalRegMap_9 | (6'h25 == architecturalRegMap_8 | (6'h25 ==
    architecturalRegMap_7 | (6'h25 == architecturalRegMap_6 | (6'h25 == architecturalRegMap_5 | (6'h25 ==
    architecturalRegMap_4 | (6'h25 == architecturalRegMap_3 | (6'h25 == architecturalRegMap_2 | (6'h25 ==
    architecturalRegMap_1 | _GEN_1239)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3160 = 6'h26 == architecturalRegMap_15 | (6'h26 == architecturalRegMap_14 | (6'h26 ==
    architecturalRegMap_13 | (6'h26 == architecturalRegMap_12 | (6'h26 == architecturalRegMap_11 | (6'h26 ==
    architecturalRegMap_10 | (6'h26 == architecturalRegMap_9 | (6'h26 == architecturalRegMap_8 | (6'h26 ==
    architecturalRegMap_7 | (6'h26 == architecturalRegMap_6 | (6'h26 == architecturalRegMap_5 | (6'h26 ==
    architecturalRegMap_4 | (6'h26 == architecturalRegMap_3 | (6'h26 == architecturalRegMap_2 | (6'h26 ==
    architecturalRegMap_1 | _GEN_1240)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3161 = 6'h27 == architecturalRegMap_15 | (6'h27 == architecturalRegMap_14 | (6'h27 ==
    architecturalRegMap_13 | (6'h27 == architecturalRegMap_12 | (6'h27 == architecturalRegMap_11 | (6'h27 ==
    architecturalRegMap_10 | (6'h27 == architecturalRegMap_9 | (6'h27 == architecturalRegMap_8 | (6'h27 ==
    architecturalRegMap_7 | (6'h27 == architecturalRegMap_6 | (6'h27 == architecturalRegMap_5 | (6'h27 ==
    architecturalRegMap_4 | (6'h27 == architecturalRegMap_3 | (6'h27 == architecturalRegMap_2 | (6'h27 ==
    architecturalRegMap_1 | _GEN_1241)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3162 = 6'h28 == architecturalRegMap_15 | (6'h28 == architecturalRegMap_14 | (6'h28 ==
    architecturalRegMap_13 | (6'h28 == architecturalRegMap_12 | (6'h28 == architecturalRegMap_11 | (6'h28 ==
    architecturalRegMap_10 | (6'h28 == architecturalRegMap_9 | (6'h28 == architecturalRegMap_8 | (6'h28 ==
    architecturalRegMap_7 | (6'h28 == architecturalRegMap_6 | (6'h28 == architecturalRegMap_5 | (6'h28 ==
    architecturalRegMap_4 | (6'h28 == architecturalRegMap_3 | (6'h28 == architecturalRegMap_2 | (6'h28 ==
    architecturalRegMap_1 | _GEN_1242)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3163 = 6'h29 == architecturalRegMap_15 | (6'h29 == architecturalRegMap_14 | (6'h29 ==
    architecturalRegMap_13 | (6'h29 == architecturalRegMap_12 | (6'h29 == architecturalRegMap_11 | (6'h29 ==
    architecturalRegMap_10 | (6'h29 == architecturalRegMap_9 | (6'h29 == architecturalRegMap_8 | (6'h29 ==
    architecturalRegMap_7 | (6'h29 == architecturalRegMap_6 | (6'h29 == architecturalRegMap_5 | (6'h29 ==
    architecturalRegMap_4 | (6'h29 == architecturalRegMap_3 | (6'h29 == architecturalRegMap_2 | (6'h29 ==
    architecturalRegMap_1 | _GEN_1243)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3164 = 6'h2a == architecturalRegMap_15 | (6'h2a == architecturalRegMap_14 | (6'h2a ==
    architecturalRegMap_13 | (6'h2a == architecturalRegMap_12 | (6'h2a == architecturalRegMap_11 | (6'h2a ==
    architecturalRegMap_10 | (6'h2a == architecturalRegMap_9 | (6'h2a == architecturalRegMap_8 | (6'h2a ==
    architecturalRegMap_7 | (6'h2a == architecturalRegMap_6 | (6'h2a == architecturalRegMap_5 | (6'h2a ==
    architecturalRegMap_4 | (6'h2a == architecturalRegMap_3 | (6'h2a == architecturalRegMap_2 | (6'h2a ==
    architecturalRegMap_1 | _GEN_1244)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3165 = 6'h2b == architecturalRegMap_15 | (6'h2b == architecturalRegMap_14 | (6'h2b ==
    architecturalRegMap_13 | (6'h2b == architecturalRegMap_12 | (6'h2b == architecturalRegMap_11 | (6'h2b ==
    architecturalRegMap_10 | (6'h2b == architecturalRegMap_9 | (6'h2b == architecturalRegMap_8 | (6'h2b ==
    architecturalRegMap_7 | (6'h2b == architecturalRegMap_6 | (6'h2b == architecturalRegMap_5 | (6'h2b ==
    architecturalRegMap_4 | (6'h2b == architecturalRegMap_3 | (6'h2b == architecturalRegMap_2 | (6'h2b ==
    architecturalRegMap_1 | _GEN_1245)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3166 = 6'h2c == architecturalRegMap_15 | (6'h2c == architecturalRegMap_14 | (6'h2c ==
    architecturalRegMap_13 | (6'h2c == architecturalRegMap_12 | (6'h2c == architecturalRegMap_11 | (6'h2c ==
    architecturalRegMap_10 | (6'h2c == architecturalRegMap_9 | (6'h2c == architecturalRegMap_8 | (6'h2c ==
    architecturalRegMap_7 | (6'h2c == architecturalRegMap_6 | (6'h2c == architecturalRegMap_5 | (6'h2c ==
    architecturalRegMap_4 | (6'h2c == architecturalRegMap_3 | (6'h2c == architecturalRegMap_2 | (6'h2c ==
    architecturalRegMap_1 | _GEN_1246)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3167 = 6'h2d == architecturalRegMap_15 | (6'h2d == architecturalRegMap_14 | (6'h2d ==
    architecturalRegMap_13 | (6'h2d == architecturalRegMap_12 | (6'h2d == architecturalRegMap_11 | (6'h2d ==
    architecturalRegMap_10 | (6'h2d == architecturalRegMap_9 | (6'h2d == architecturalRegMap_8 | (6'h2d ==
    architecturalRegMap_7 | (6'h2d == architecturalRegMap_6 | (6'h2d == architecturalRegMap_5 | (6'h2d ==
    architecturalRegMap_4 | (6'h2d == architecturalRegMap_3 | (6'h2d == architecturalRegMap_2 | (6'h2d ==
    architecturalRegMap_1 | _GEN_1247)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3168 = 6'h2e == architecturalRegMap_15 | (6'h2e == architecturalRegMap_14 | (6'h2e ==
    architecturalRegMap_13 | (6'h2e == architecturalRegMap_12 | (6'h2e == architecturalRegMap_11 | (6'h2e ==
    architecturalRegMap_10 | (6'h2e == architecturalRegMap_9 | (6'h2e == architecturalRegMap_8 | (6'h2e ==
    architecturalRegMap_7 | (6'h2e == architecturalRegMap_6 | (6'h2e == architecturalRegMap_5 | (6'h2e ==
    architecturalRegMap_4 | (6'h2e == architecturalRegMap_3 | (6'h2e == architecturalRegMap_2 | (6'h2e ==
    architecturalRegMap_1 | _GEN_1248)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3169 = 6'h2f == architecturalRegMap_15 | (6'h2f == architecturalRegMap_14 | (6'h2f ==
    architecturalRegMap_13 | (6'h2f == architecturalRegMap_12 | (6'h2f == architecturalRegMap_11 | (6'h2f ==
    architecturalRegMap_10 | (6'h2f == architecturalRegMap_9 | (6'h2f == architecturalRegMap_8 | (6'h2f ==
    architecturalRegMap_7 | (6'h2f == architecturalRegMap_6 | (6'h2f == architecturalRegMap_5 | (6'h2f ==
    architecturalRegMap_4 | (6'h2f == architecturalRegMap_3 | (6'h2f == architecturalRegMap_2 | (6'h2f ==
    architecturalRegMap_1 | _GEN_1249)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3170 = 6'h30 == architecturalRegMap_15 | (6'h30 == architecturalRegMap_14 | (6'h30 ==
    architecturalRegMap_13 | (6'h30 == architecturalRegMap_12 | (6'h30 == architecturalRegMap_11 | (6'h30 ==
    architecturalRegMap_10 | (6'h30 == architecturalRegMap_9 | (6'h30 == architecturalRegMap_8 | (6'h30 ==
    architecturalRegMap_7 | (6'h30 == architecturalRegMap_6 | (6'h30 == architecturalRegMap_5 | (6'h30 ==
    architecturalRegMap_4 | (6'h30 == architecturalRegMap_3 | (6'h30 == architecturalRegMap_2 | (6'h30 ==
    architecturalRegMap_1 | _GEN_1250)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3171 = 6'h31 == architecturalRegMap_15 | (6'h31 == architecturalRegMap_14 | (6'h31 ==
    architecturalRegMap_13 | (6'h31 == architecturalRegMap_12 | (6'h31 == architecturalRegMap_11 | (6'h31 ==
    architecturalRegMap_10 | (6'h31 == architecturalRegMap_9 | (6'h31 == architecturalRegMap_8 | (6'h31 ==
    architecturalRegMap_7 | (6'h31 == architecturalRegMap_6 | (6'h31 == architecturalRegMap_5 | (6'h31 ==
    architecturalRegMap_4 | (6'h31 == architecturalRegMap_3 | (6'h31 == architecturalRegMap_2 | (6'h31 ==
    architecturalRegMap_1 | _GEN_1251)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3172 = 6'h32 == architecturalRegMap_15 | (6'h32 == architecturalRegMap_14 | (6'h32 ==
    architecturalRegMap_13 | (6'h32 == architecturalRegMap_12 | (6'h32 == architecturalRegMap_11 | (6'h32 ==
    architecturalRegMap_10 | (6'h32 == architecturalRegMap_9 | (6'h32 == architecturalRegMap_8 | (6'h32 ==
    architecturalRegMap_7 | (6'h32 == architecturalRegMap_6 | (6'h32 == architecturalRegMap_5 | (6'h32 ==
    architecturalRegMap_4 | (6'h32 == architecturalRegMap_3 | (6'h32 == architecturalRegMap_2 | (6'h32 ==
    architecturalRegMap_1 | _GEN_1252)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3173 = 6'h33 == architecturalRegMap_15 | (6'h33 == architecturalRegMap_14 | (6'h33 ==
    architecturalRegMap_13 | (6'h33 == architecturalRegMap_12 | (6'h33 == architecturalRegMap_11 | (6'h33 ==
    architecturalRegMap_10 | (6'h33 == architecturalRegMap_9 | (6'h33 == architecturalRegMap_8 | (6'h33 ==
    architecturalRegMap_7 | (6'h33 == architecturalRegMap_6 | (6'h33 == architecturalRegMap_5 | (6'h33 ==
    architecturalRegMap_4 | (6'h33 == architecturalRegMap_3 | (6'h33 == architecturalRegMap_2 | (6'h33 ==
    architecturalRegMap_1 | _GEN_1253)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3174 = 6'h34 == architecturalRegMap_15 | (6'h34 == architecturalRegMap_14 | (6'h34 ==
    architecturalRegMap_13 | (6'h34 == architecturalRegMap_12 | (6'h34 == architecturalRegMap_11 | (6'h34 ==
    architecturalRegMap_10 | (6'h34 == architecturalRegMap_9 | (6'h34 == architecturalRegMap_8 | (6'h34 ==
    architecturalRegMap_7 | (6'h34 == architecturalRegMap_6 | (6'h34 == architecturalRegMap_5 | (6'h34 ==
    architecturalRegMap_4 | (6'h34 == architecturalRegMap_3 | (6'h34 == architecturalRegMap_2 | (6'h34 ==
    architecturalRegMap_1 | _GEN_1254)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3175 = 6'h35 == architecturalRegMap_15 | (6'h35 == architecturalRegMap_14 | (6'h35 ==
    architecturalRegMap_13 | (6'h35 == architecturalRegMap_12 | (6'h35 == architecturalRegMap_11 | (6'h35 ==
    architecturalRegMap_10 | (6'h35 == architecturalRegMap_9 | (6'h35 == architecturalRegMap_8 | (6'h35 ==
    architecturalRegMap_7 | (6'h35 == architecturalRegMap_6 | (6'h35 == architecturalRegMap_5 | (6'h35 ==
    architecturalRegMap_4 | (6'h35 == architecturalRegMap_3 | (6'h35 == architecturalRegMap_2 | (6'h35 ==
    architecturalRegMap_1 | _GEN_1255)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3176 = 6'h36 == architecturalRegMap_15 | (6'h36 == architecturalRegMap_14 | (6'h36 ==
    architecturalRegMap_13 | (6'h36 == architecturalRegMap_12 | (6'h36 == architecturalRegMap_11 | (6'h36 ==
    architecturalRegMap_10 | (6'h36 == architecturalRegMap_9 | (6'h36 == architecturalRegMap_8 | (6'h36 ==
    architecturalRegMap_7 | (6'h36 == architecturalRegMap_6 | (6'h36 == architecturalRegMap_5 | (6'h36 ==
    architecturalRegMap_4 | (6'h36 == architecturalRegMap_3 | (6'h36 == architecturalRegMap_2 | (6'h36 ==
    architecturalRegMap_1 | _GEN_1256)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3177 = 6'h37 == architecturalRegMap_15 | (6'h37 == architecturalRegMap_14 | (6'h37 ==
    architecturalRegMap_13 | (6'h37 == architecturalRegMap_12 | (6'h37 == architecturalRegMap_11 | (6'h37 ==
    architecturalRegMap_10 | (6'h37 == architecturalRegMap_9 | (6'h37 == architecturalRegMap_8 | (6'h37 ==
    architecturalRegMap_7 | (6'h37 == architecturalRegMap_6 | (6'h37 == architecturalRegMap_5 | (6'h37 ==
    architecturalRegMap_4 | (6'h37 == architecturalRegMap_3 | (6'h37 == architecturalRegMap_2 | (6'h37 ==
    architecturalRegMap_1 | _GEN_1257)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3178 = 6'h38 == architecturalRegMap_15 | (6'h38 == architecturalRegMap_14 | (6'h38 ==
    architecturalRegMap_13 | (6'h38 == architecturalRegMap_12 | (6'h38 == architecturalRegMap_11 | (6'h38 ==
    architecturalRegMap_10 | (6'h38 == architecturalRegMap_9 | (6'h38 == architecturalRegMap_8 | (6'h38 ==
    architecturalRegMap_7 | (6'h38 == architecturalRegMap_6 | (6'h38 == architecturalRegMap_5 | (6'h38 ==
    architecturalRegMap_4 | (6'h38 == architecturalRegMap_3 | (6'h38 == architecturalRegMap_2 | (6'h38 ==
    architecturalRegMap_1 | _GEN_1258)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3179 = 6'h39 == architecturalRegMap_15 | (6'h39 == architecturalRegMap_14 | (6'h39 ==
    architecturalRegMap_13 | (6'h39 == architecturalRegMap_12 | (6'h39 == architecturalRegMap_11 | (6'h39 ==
    architecturalRegMap_10 | (6'h39 == architecturalRegMap_9 | (6'h39 == architecturalRegMap_8 | (6'h39 ==
    architecturalRegMap_7 | (6'h39 == architecturalRegMap_6 | (6'h39 == architecturalRegMap_5 | (6'h39 ==
    architecturalRegMap_4 | (6'h39 == architecturalRegMap_3 | (6'h39 == architecturalRegMap_2 | (6'h39 ==
    architecturalRegMap_1 | _GEN_1259)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3180 = 6'h3a == architecturalRegMap_15 | (6'h3a == architecturalRegMap_14 | (6'h3a ==
    architecturalRegMap_13 | (6'h3a == architecturalRegMap_12 | (6'h3a == architecturalRegMap_11 | (6'h3a ==
    architecturalRegMap_10 | (6'h3a == architecturalRegMap_9 | (6'h3a == architecturalRegMap_8 | (6'h3a ==
    architecturalRegMap_7 | (6'h3a == architecturalRegMap_6 | (6'h3a == architecturalRegMap_5 | (6'h3a ==
    architecturalRegMap_4 | (6'h3a == architecturalRegMap_3 | (6'h3a == architecturalRegMap_2 | (6'h3a ==
    architecturalRegMap_1 | _GEN_1260)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3181 = 6'h3b == architecturalRegMap_15 | (6'h3b == architecturalRegMap_14 | (6'h3b ==
    architecturalRegMap_13 | (6'h3b == architecturalRegMap_12 | (6'h3b == architecturalRegMap_11 | (6'h3b ==
    architecturalRegMap_10 | (6'h3b == architecturalRegMap_9 | (6'h3b == architecturalRegMap_8 | (6'h3b ==
    architecturalRegMap_7 | (6'h3b == architecturalRegMap_6 | (6'h3b == architecturalRegMap_5 | (6'h3b ==
    architecturalRegMap_4 | (6'h3b == architecturalRegMap_3 | (6'h3b == architecturalRegMap_2 | (6'h3b ==
    architecturalRegMap_1 | _GEN_1261)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3182 = 6'h3c == architecturalRegMap_15 | (6'h3c == architecturalRegMap_14 | (6'h3c ==
    architecturalRegMap_13 | (6'h3c == architecturalRegMap_12 | (6'h3c == architecturalRegMap_11 | (6'h3c ==
    architecturalRegMap_10 | (6'h3c == architecturalRegMap_9 | (6'h3c == architecturalRegMap_8 | (6'h3c ==
    architecturalRegMap_7 | (6'h3c == architecturalRegMap_6 | (6'h3c == architecturalRegMap_5 | (6'h3c ==
    architecturalRegMap_4 | (6'h3c == architecturalRegMap_3 | (6'h3c == architecturalRegMap_2 | (6'h3c ==
    architecturalRegMap_1 | _GEN_1262)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3183 = 6'h3d == architecturalRegMap_15 | (6'h3d == architecturalRegMap_14 | (6'h3d ==
    architecturalRegMap_13 | (6'h3d == architecturalRegMap_12 | (6'h3d == architecturalRegMap_11 | (6'h3d ==
    architecturalRegMap_10 | (6'h3d == architecturalRegMap_9 | (6'h3d == architecturalRegMap_8 | (6'h3d ==
    architecturalRegMap_7 | (6'h3d == architecturalRegMap_6 | (6'h3d == architecturalRegMap_5 | (6'h3d ==
    architecturalRegMap_4 | (6'h3d == architecturalRegMap_3 | (6'h3d == architecturalRegMap_2 | (6'h3d ==
    architecturalRegMap_1 | _GEN_1263)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3184 = 6'h3e == architecturalRegMap_15 | (6'h3e == architecturalRegMap_14 | (6'h3e ==
    architecturalRegMap_13 | (6'h3e == architecturalRegMap_12 | (6'h3e == architecturalRegMap_11 | (6'h3e ==
    architecturalRegMap_10 | (6'h3e == architecturalRegMap_9 | (6'h3e == architecturalRegMap_8 | (6'h3e ==
    architecturalRegMap_7 | (6'h3e == architecturalRegMap_6 | (6'h3e == architecturalRegMap_5 | (6'h3e ==
    architecturalRegMap_4 | (6'h3e == architecturalRegMap_3 | (6'h3e == architecturalRegMap_2 | (6'h3e ==
    architecturalRegMap_1 | _GEN_1264)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3185 = 6'h3f == architecturalRegMap_15 | (6'h3f == architecturalRegMap_14 | (6'h3f ==
    architecturalRegMap_13 | (6'h3f == architecturalRegMap_12 | (6'h3f == architecturalRegMap_11 | (6'h3f ==
    architecturalRegMap_10 | (6'h3f == architecturalRegMap_9 | (6'h3f == architecturalRegMap_8 | (6'h3f ==
    architecturalRegMap_7 | (6'h3f == architecturalRegMap_6 | (6'h3f == architecturalRegMap_5 | (6'h3f ==
    architecturalRegMap_4 | (6'h3f == architecturalRegMap_3 | (6'h3f == architecturalRegMap_2 | (6'h3f ==
    architecturalRegMap_1 | _GEN_1265)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_3186 = 6'h0 == architecturalRegMap_15 ? 1'h0 : _GEN_3058; // @[decode.scala 393:{46,46}]
  wire  _GEN_3187 = 6'h1 == architecturalRegMap_15 ? 1'h0 : _GEN_3059; // @[decode.scala 393:{46,46}]
  wire  _GEN_3188 = 6'h2 == architecturalRegMap_15 ? 1'h0 : _GEN_3060; // @[decode.scala 393:{46,46}]
  wire  _GEN_3189 = 6'h3 == architecturalRegMap_15 ? 1'h0 : _GEN_3061; // @[decode.scala 393:{46,46}]
  wire  _GEN_3190 = 6'h4 == architecturalRegMap_15 ? 1'h0 : _GEN_3062; // @[decode.scala 393:{46,46}]
  wire  _GEN_3191 = 6'h5 == architecturalRegMap_15 ? 1'h0 : _GEN_3063; // @[decode.scala 393:{46,46}]
  wire  _GEN_3192 = 6'h6 == architecturalRegMap_15 ? 1'h0 : _GEN_3064; // @[decode.scala 393:{46,46}]
  wire  _GEN_3193 = 6'h7 == architecturalRegMap_15 ? 1'h0 : _GEN_3065; // @[decode.scala 393:{46,46}]
  wire  _GEN_3194 = 6'h8 == architecturalRegMap_15 ? 1'h0 : _GEN_3066; // @[decode.scala 393:{46,46}]
  wire  _GEN_3195 = 6'h9 == architecturalRegMap_15 ? 1'h0 : _GEN_3067; // @[decode.scala 393:{46,46}]
  wire  _GEN_3196 = 6'ha == architecturalRegMap_15 ? 1'h0 : _GEN_3068; // @[decode.scala 393:{46,46}]
  wire  _GEN_3197 = 6'hb == architecturalRegMap_15 ? 1'h0 : _GEN_3069; // @[decode.scala 393:{46,46}]
  wire  _GEN_3198 = 6'hc == architecturalRegMap_15 ? 1'h0 : _GEN_3070; // @[decode.scala 393:{46,46}]
  wire  _GEN_3199 = 6'hd == architecturalRegMap_15 ? 1'h0 : _GEN_3071; // @[decode.scala 393:{46,46}]
  wire  _GEN_3200 = 6'he == architecturalRegMap_15 ? 1'h0 : _GEN_3072; // @[decode.scala 393:{46,46}]
  wire  _GEN_3201 = 6'hf == architecturalRegMap_15 ? 1'h0 : _GEN_3073; // @[decode.scala 393:{46,46}]
  wire  _GEN_3202 = 6'h10 == architecturalRegMap_15 ? 1'h0 : _GEN_3074; // @[decode.scala 393:{46,46}]
  wire  _GEN_3203 = 6'h11 == architecturalRegMap_15 ? 1'h0 : _GEN_3075; // @[decode.scala 393:{46,46}]
  wire  _GEN_3204 = 6'h12 == architecturalRegMap_15 ? 1'h0 : _GEN_3076; // @[decode.scala 393:{46,46}]
  wire  _GEN_3205 = 6'h13 == architecturalRegMap_15 ? 1'h0 : _GEN_3077; // @[decode.scala 393:{46,46}]
  wire  _GEN_3206 = 6'h14 == architecturalRegMap_15 ? 1'h0 : _GEN_3078; // @[decode.scala 393:{46,46}]
  wire  _GEN_3207 = 6'h15 == architecturalRegMap_15 ? 1'h0 : _GEN_3079; // @[decode.scala 393:{46,46}]
  wire  _GEN_3208 = 6'h16 == architecturalRegMap_15 ? 1'h0 : _GEN_3080; // @[decode.scala 393:{46,46}]
  wire  _GEN_3209 = 6'h17 == architecturalRegMap_15 ? 1'h0 : _GEN_3081; // @[decode.scala 393:{46,46}]
  wire  _GEN_3210 = 6'h18 == architecturalRegMap_15 ? 1'h0 : _GEN_3082; // @[decode.scala 393:{46,46}]
  wire  _GEN_3211 = 6'h19 == architecturalRegMap_15 ? 1'h0 : _GEN_3083; // @[decode.scala 393:{46,46}]
  wire  _GEN_3212 = 6'h1a == architecturalRegMap_15 ? 1'h0 : _GEN_3084; // @[decode.scala 393:{46,46}]
  wire  _GEN_3213 = 6'h1b == architecturalRegMap_15 ? 1'h0 : _GEN_3085; // @[decode.scala 393:{46,46}]
  wire  _GEN_3214 = 6'h1c == architecturalRegMap_15 ? 1'h0 : _GEN_3086; // @[decode.scala 393:{46,46}]
  wire  _GEN_3215 = 6'h1d == architecturalRegMap_15 ? 1'h0 : _GEN_3087; // @[decode.scala 393:{46,46}]
  wire  _GEN_3216 = 6'h1e == architecturalRegMap_15 ? 1'h0 : _GEN_3088; // @[decode.scala 393:{46,46}]
  wire  _GEN_3217 = 6'h1f == architecturalRegMap_15 ? 1'h0 : _GEN_3089; // @[decode.scala 393:{46,46}]
  wire  _GEN_3218 = 6'h20 == architecturalRegMap_15 ? 1'h0 : _GEN_3090; // @[decode.scala 393:{46,46}]
  wire  _GEN_3219 = 6'h21 == architecturalRegMap_15 ? 1'h0 : _GEN_3091; // @[decode.scala 393:{46,46}]
  wire  _GEN_3220 = 6'h22 == architecturalRegMap_15 ? 1'h0 : _GEN_3092; // @[decode.scala 393:{46,46}]
  wire  _GEN_3221 = 6'h23 == architecturalRegMap_15 ? 1'h0 : _GEN_3093; // @[decode.scala 393:{46,46}]
  wire  _GEN_3222 = 6'h24 == architecturalRegMap_15 ? 1'h0 : _GEN_3094; // @[decode.scala 393:{46,46}]
  wire  _GEN_3223 = 6'h25 == architecturalRegMap_15 ? 1'h0 : _GEN_3095; // @[decode.scala 393:{46,46}]
  wire  _GEN_3224 = 6'h26 == architecturalRegMap_15 ? 1'h0 : _GEN_3096; // @[decode.scala 393:{46,46}]
  wire  _GEN_3225 = 6'h27 == architecturalRegMap_15 ? 1'h0 : _GEN_3097; // @[decode.scala 393:{46,46}]
  wire  _GEN_3226 = 6'h28 == architecturalRegMap_15 ? 1'h0 : _GEN_3098; // @[decode.scala 393:{46,46}]
  wire  _GEN_3227 = 6'h29 == architecturalRegMap_15 ? 1'h0 : _GEN_3099; // @[decode.scala 393:{46,46}]
  wire  _GEN_3228 = 6'h2a == architecturalRegMap_15 ? 1'h0 : _GEN_3100; // @[decode.scala 393:{46,46}]
  wire  _GEN_3229 = 6'h2b == architecturalRegMap_15 ? 1'h0 : _GEN_3101; // @[decode.scala 393:{46,46}]
  wire  _GEN_3230 = 6'h2c == architecturalRegMap_15 ? 1'h0 : _GEN_3102; // @[decode.scala 393:{46,46}]
  wire  _GEN_3231 = 6'h2d == architecturalRegMap_15 ? 1'h0 : _GEN_3103; // @[decode.scala 393:{46,46}]
  wire  _GEN_3232 = 6'h2e == architecturalRegMap_15 ? 1'h0 : _GEN_3104; // @[decode.scala 393:{46,46}]
  wire  _GEN_3233 = 6'h2f == architecturalRegMap_15 ? 1'h0 : _GEN_3105; // @[decode.scala 393:{46,46}]
  wire  _GEN_3234 = 6'h30 == architecturalRegMap_15 ? 1'h0 : _GEN_3106; // @[decode.scala 393:{46,46}]
  wire  _GEN_3235 = 6'h31 == architecturalRegMap_15 ? 1'h0 : _GEN_3107; // @[decode.scala 393:{46,46}]
  wire  _GEN_3236 = 6'h32 == architecturalRegMap_15 ? 1'h0 : _GEN_3108; // @[decode.scala 393:{46,46}]
  wire  _GEN_3237 = 6'h33 == architecturalRegMap_15 ? 1'h0 : _GEN_3109; // @[decode.scala 393:{46,46}]
  wire  _GEN_3238 = 6'h34 == architecturalRegMap_15 ? 1'h0 : _GEN_3110; // @[decode.scala 393:{46,46}]
  wire  _GEN_3239 = 6'h35 == architecturalRegMap_15 ? 1'h0 : _GEN_3111; // @[decode.scala 393:{46,46}]
  wire  _GEN_3240 = 6'h36 == architecturalRegMap_15 ? 1'h0 : _GEN_3112; // @[decode.scala 393:{46,46}]
  wire  _GEN_3241 = 6'h37 == architecturalRegMap_15 ? 1'h0 : _GEN_3113; // @[decode.scala 393:{46,46}]
  wire  _GEN_3242 = 6'h38 == architecturalRegMap_15 ? 1'h0 : _GEN_3114; // @[decode.scala 393:{46,46}]
  wire  _GEN_3243 = 6'h39 == architecturalRegMap_15 ? 1'h0 : _GEN_3115; // @[decode.scala 393:{46,46}]
  wire  _GEN_3244 = 6'h3a == architecturalRegMap_15 ? 1'h0 : _GEN_3116; // @[decode.scala 393:{46,46}]
  wire  _GEN_3245 = 6'h3b == architecturalRegMap_15 ? 1'h0 : _GEN_3117; // @[decode.scala 393:{46,46}]
  wire  _GEN_3246 = 6'h3c == architecturalRegMap_15 ? 1'h0 : _GEN_3118; // @[decode.scala 393:{46,46}]
  wire  _GEN_3247 = 6'h3d == architecturalRegMap_15 ? 1'h0 : _GEN_3119; // @[decode.scala 393:{46,46}]
  wire  _GEN_3248 = 6'h3e == architecturalRegMap_15 ? 1'h0 : _GEN_3120; // @[decode.scala 393:{46,46}]
  wire  _GEN_3314 = 6'h0 == architecturalRegMap_16 ? 1'h0 : _GEN_3186; // @[decode.scala 393:{46,46}]
  wire  _GEN_3315 = 6'h1 == architecturalRegMap_16 ? 1'h0 : _GEN_3187; // @[decode.scala 393:{46,46}]
  wire  _GEN_3316 = 6'h2 == architecturalRegMap_16 ? 1'h0 : _GEN_3188; // @[decode.scala 393:{46,46}]
  wire  _GEN_3317 = 6'h3 == architecturalRegMap_16 ? 1'h0 : _GEN_3189; // @[decode.scala 393:{46,46}]
  wire  _GEN_3318 = 6'h4 == architecturalRegMap_16 ? 1'h0 : _GEN_3190; // @[decode.scala 393:{46,46}]
  wire  _GEN_3319 = 6'h5 == architecturalRegMap_16 ? 1'h0 : _GEN_3191; // @[decode.scala 393:{46,46}]
  wire  _GEN_3320 = 6'h6 == architecturalRegMap_16 ? 1'h0 : _GEN_3192; // @[decode.scala 393:{46,46}]
  wire  _GEN_3321 = 6'h7 == architecturalRegMap_16 ? 1'h0 : _GEN_3193; // @[decode.scala 393:{46,46}]
  wire  _GEN_3322 = 6'h8 == architecturalRegMap_16 ? 1'h0 : _GEN_3194; // @[decode.scala 393:{46,46}]
  wire  _GEN_3323 = 6'h9 == architecturalRegMap_16 ? 1'h0 : _GEN_3195; // @[decode.scala 393:{46,46}]
  wire  _GEN_3324 = 6'ha == architecturalRegMap_16 ? 1'h0 : _GEN_3196; // @[decode.scala 393:{46,46}]
  wire  _GEN_3325 = 6'hb == architecturalRegMap_16 ? 1'h0 : _GEN_3197; // @[decode.scala 393:{46,46}]
  wire  _GEN_3326 = 6'hc == architecturalRegMap_16 ? 1'h0 : _GEN_3198; // @[decode.scala 393:{46,46}]
  wire  _GEN_3327 = 6'hd == architecturalRegMap_16 ? 1'h0 : _GEN_3199; // @[decode.scala 393:{46,46}]
  wire  _GEN_3328 = 6'he == architecturalRegMap_16 ? 1'h0 : _GEN_3200; // @[decode.scala 393:{46,46}]
  wire  _GEN_3329 = 6'hf == architecturalRegMap_16 ? 1'h0 : _GEN_3201; // @[decode.scala 393:{46,46}]
  wire  _GEN_3330 = 6'h10 == architecturalRegMap_16 ? 1'h0 : _GEN_3202; // @[decode.scala 393:{46,46}]
  wire  _GEN_3331 = 6'h11 == architecturalRegMap_16 ? 1'h0 : _GEN_3203; // @[decode.scala 393:{46,46}]
  wire  _GEN_3332 = 6'h12 == architecturalRegMap_16 ? 1'h0 : _GEN_3204; // @[decode.scala 393:{46,46}]
  wire  _GEN_3333 = 6'h13 == architecturalRegMap_16 ? 1'h0 : _GEN_3205; // @[decode.scala 393:{46,46}]
  wire  _GEN_3334 = 6'h14 == architecturalRegMap_16 ? 1'h0 : _GEN_3206; // @[decode.scala 393:{46,46}]
  wire  _GEN_3335 = 6'h15 == architecturalRegMap_16 ? 1'h0 : _GEN_3207; // @[decode.scala 393:{46,46}]
  wire  _GEN_3336 = 6'h16 == architecturalRegMap_16 ? 1'h0 : _GEN_3208; // @[decode.scala 393:{46,46}]
  wire  _GEN_3337 = 6'h17 == architecturalRegMap_16 ? 1'h0 : _GEN_3209; // @[decode.scala 393:{46,46}]
  wire  _GEN_3338 = 6'h18 == architecturalRegMap_16 ? 1'h0 : _GEN_3210; // @[decode.scala 393:{46,46}]
  wire  _GEN_3339 = 6'h19 == architecturalRegMap_16 ? 1'h0 : _GEN_3211; // @[decode.scala 393:{46,46}]
  wire  _GEN_3340 = 6'h1a == architecturalRegMap_16 ? 1'h0 : _GEN_3212; // @[decode.scala 393:{46,46}]
  wire  _GEN_3341 = 6'h1b == architecturalRegMap_16 ? 1'h0 : _GEN_3213; // @[decode.scala 393:{46,46}]
  wire  _GEN_3342 = 6'h1c == architecturalRegMap_16 ? 1'h0 : _GEN_3214; // @[decode.scala 393:{46,46}]
  wire  _GEN_3343 = 6'h1d == architecturalRegMap_16 ? 1'h0 : _GEN_3215; // @[decode.scala 393:{46,46}]
  wire  _GEN_3344 = 6'h1e == architecturalRegMap_16 ? 1'h0 : _GEN_3216; // @[decode.scala 393:{46,46}]
  wire  _GEN_3345 = 6'h1f == architecturalRegMap_16 ? 1'h0 : _GEN_3217; // @[decode.scala 393:{46,46}]
  wire  _GEN_3346 = 6'h20 == architecturalRegMap_16 ? 1'h0 : _GEN_3218; // @[decode.scala 393:{46,46}]
  wire  _GEN_3347 = 6'h21 == architecturalRegMap_16 ? 1'h0 : _GEN_3219; // @[decode.scala 393:{46,46}]
  wire  _GEN_3348 = 6'h22 == architecturalRegMap_16 ? 1'h0 : _GEN_3220; // @[decode.scala 393:{46,46}]
  wire  _GEN_3349 = 6'h23 == architecturalRegMap_16 ? 1'h0 : _GEN_3221; // @[decode.scala 393:{46,46}]
  wire  _GEN_3350 = 6'h24 == architecturalRegMap_16 ? 1'h0 : _GEN_3222; // @[decode.scala 393:{46,46}]
  wire  _GEN_3351 = 6'h25 == architecturalRegMap_16 ? 1'h0 : _GEN_3223; // @[decode.scala 393:{46,46}]
  wire  _GEN_3352 = 6'h26 == architecturalRegMap_16 ? 1'h0 : _GEN_3224; // @[decode.scala 393:{46,46}]
  wire  _GEN_3353 = 6'h27 == architecturalRegMap_16 ? 1'h0 : _GEN_3225; // @[decode.scala 393:{46,46}]
  wire  _GEN_3354 = 6'h28 == architecturalRegMap_16 ? 1'h0 : _GEN_3226; // @[decode.scala 393:{46,46}]
  wire  _GEN_3355 = 6'h29 == architecturalRegMap_16 ? 1'h0 : _GEN_3227; // @[decode.scala 393:{46,46}]
  wire  _GEN_3356 = 6'h2a == architecturalRegMap_16 ? 1'h0 : _GEN_3228; // @[decode.scala 393:{46,46}]
  wire  _GEN_3357 = 6'h2b == architecturalRegMap_16 ? 1'h0 : _GEN_3229; // @[decode.scala 393:{46,46}]
  wire  _GEN_3358 = 6'h2c == architecturalRegMap_16 ? 1'h0 : _GEN_3230; // @[decode.scala 393:{46,46}]
  wire  _GEN_3359 = 6'h2d == architecturalRegMap_16 ? 1'h0 : _GEN_3231; // @[decode.scala 393:{46,46}]
  wire  _GEN_3360 = 6'h2e == architecturalRegMap_16 ? 1'h0 : _GEN_3232; // @[decode.scala 393:{46,46}]
  wire  _GEN_3361 = 6'h2f == architecturalRegMap_16 ? 1'h0 : _GEN_3233; // @[decode.scala 393:{46,46}]
  wire  _GEN_3362 = 6'h30 == architecturalRegMap_16 ? 1'h0 : _GEN_3234; // @[decode.scala 393:{46,46}]
  wire  _GEN_3363 = 6'h31 == architecturalRegMap_16 ? 1'h0 : _GEN_3235; // @[decode.scala 393:{46,46}]
  wire  _GEN_3364 = 6'h32 == architecturalRegMap_16 ? 1'h0 : _GEN_3236; // @[decode.scala 393:{46,46}]
  wire  _GEN_3365 = 6'h33 == architecturalRegMap_16 ? 1'h0 : _GEN_3237; // @[decode.scala 393:{46,46}]
  wire  _GEN_3366 = 6'h34 == architecturalRegMap_16 ? 1'h0 : _GEN_3238; // @[decode.scala 393:{46,46}]
  wire  _GEN_3367 = 6'h35 == architecturalRegMap_16 ? 1'h0 : _GEN_3239; // @[decode.scala 393:{46,46}]
  wire  _GEN_3368 = 6'h36 == architecturalRegMap_16 ? 1'h0 : _GEN_3240; // @[decode.scala 393:{46,46}]
  wire  _GEN_3369 = 6'h37 == architecturalRegMap_16 ? 1'h0 : _GEN_3241; // @[decode.scala 393:{46,46}]
  wire  _GEN_3370 = 6'h38 == architecturalRegMap_16 ? 1'h0 : _GEN_3242; // @[decode.scala 393:{46,46}]
  wire  _GEN_3371 = 6'h39 == architecturalRegMap_16 ? 1'h0 : _GEN_3243; // @[decode.scala 393:{46,46}]
  wire  _GEN_3372 = 6'h3a == architecturalRegMap_16 ? 1'h0 : _GEN_3244; // @[decode.scala 393:{46,46}]
  wire  _GEN_3373 = 6'h3b == architecturalRegMap_16 ? 1'h0 : _GEN_3245; // @[decode.scala 393:{46,46}]
  wire  _GEN_3374 = 6'h3c == architecturalRegMap_16 ? 1'h0 : _GEN_3246; // @[decode.scala 393:{46,46}]
  wire  _GEN_3375 = 6'h3d == architecturalRegMap_16 ? 1'h0 : _GEN_3247; // @[decode.scala 393:{46,46}]
  wire  _GEN_3376 = 6'h3e == architecturalRegMap_16 ? 1'h0 : _GEN_3248; // @[decode.scala 393:{46,46}]
  wire  _GEN_3442 = 6'h0 == architecturalRegMap_17 ? 1'h0 : _GEN_3314; // @[decode.scala 393:{46,46}]
  wire  _GEN_3443 = 6'h1 == architecturalRegMap_17 ? 1'h0 : _GEN_3315; // @[decode.scala 393:{46,46}]
  wire  _GEN_3444 = 6'h2 == architecturalRegMap_17 ? 1'h0 : _GEN_3316; // @[decode.scala 393:{46,46}]
  wire  _GEN_3445 = 6'h3 == architecturalRegMap_17 ? 1'h0 : _GEN_3317; // @[decode.scala 393:{46,46}]
  wire  _GEN_3446 = 6'h4 == architecturalRegMap_17 ? 1'h0 : _GEN_3318; // @[decode.scala 393:{46,46}]
  wire  _GEN_3447 = 6'h5 == architecturalRegMap_17 ? 1'h0 : _GEN_3319; // @[decode.scala 393:{46,46}]
  wire  _GEN_3448 = 6'h6 == architecturalRegMap_17 ? 1'h0 : _GEN_3320; // @[decode.scala 393:{46,46}]
  wire  _GEN_3449 = 6'h7 == architecturalRegMap_17 ? 1'h0 : _GEN_3321; // @[decode.scala 393:{46,46}]
  wire  _GEN_3450 = 6'h8 == architecturalRegMap_17 ? 1'h0 : _GEN_3322; // @[decode.scala 393:{46,46}]
  wire  _GEN_3451 = 6'h9 == architecturalRegMap_17 ? 1'h0 : _GEN_3323; // @[decode.scala 393:{46,46}]
  wire  _GEN_3452 = 6'ha == architecturalRegMap_17 ? 1'h0 : _GEN_3324; // @[decode.scala 393:{46,46}]
  wire  _GEN_3453 = 6'hb == architecturalRegMap_17 ? 1'h0 : _GEN_3325; // @[decode.scala 393:{46,46}]
  wire  _GEN_3454 = 6'hc == architecturalRegMap_17 ? 1'h0 : _GEN_3326; // @[decode.scala 393:{46,46}]
  wire  _GEN_3455 = 6'hd == architecturalRegMap_17 ? 1'h0 : _GEN_3327; // @[decode.scala 393:{46,46}]
  wire  _GEN_3456 = 6'he == architecturalRegMap_17 ? 1'h0 : _GEN_3328; // @[decode.scala 393:{46,46}]
  wire  _GEN_3457 = 6'hf == architecturalRegMap_17 ? 1'h0 : _GEN_3329; // @[decode.scala 393:{46,46}]
  wire  _GEN_3458 = 6'h10 == architecturalRegMap_17 ? 1'h0 : _GEN_3330; // @[decode.scala 393:{46,46}]
  wire  _GEN_3459 = 6'h11 == architecturalRegMap_17 ? 1'h0 : _GEN_3331; // @[decode.scala 393:{46,46}]
  wire  _GEN_3460 = 6'h12 == architecturalRegMap_17 ? 1'h0 : _GEN_3332; // @[decode.scala 393:{46,46}]
  wire  _GEN_3461 = 6'h13 == architecturalRegMap_17 ? 1'h0 : _GEN_3333; // @[decode.scala 393:{46,46}]
  wire  _GEN_3462 = 6'h14 == architecturalRegMap_17 ? 1'h0 : _GEN_3334; // @[decode.scala 393:{46,46}]
  wire  _GEN_3463 = 6'h15 == architecturalRegMap_17 ? 1'h0 : _GEN_3335; // @[decode.scala 393:{46,46}]
  wire  _GEN_3464 = 6'h16 == architecturalRegMap_17 ? 1'h0 : _GEN_3336; // @[decode.scala 393:{46,46}]
  wire  _GEN_3465 = 6'h17 == architecturalRegMap_17 ? 1'h0 : _GEN_3337; // @[decode.scala 393:{46,46}]
  wire  _GEN_3466 = 6'h18 == architecturalRegMap_17 ? 1'h0 : _GEN_3338; // @[decode.scala 393:{46,46}]
  wire  _GEN_3467 = 6'h19 == architecturalRegMap_17 ? 1'h0 : _GEN_3339; // @[decode.scala 393:{46,46}]
  wire  _GEN_3468 = 6'h1a == architecturalRegMap_17 ? 1'h0 : _GEN_3340; // @[decode.scala 393:{46,46}]
  wire  _GEN_3469 = 6'h1b == architecturalRegMap_17 ? 1'h0 : _GEN_3341; // @[decode.scala 393:{46,46}]
  wire  _GEN_3470 = 6'h1c == architecturalRegMap_17 ? 1'h0 : _GEN_3342; // @[decode.scala 393:{46,46}]
  wire  _GEN_3471 = 6'h1d == architecturalRegMap_17 ? 1'h0 : _GEN_3343; // @[decode.scala 393:{46,46}]
  wire  _GEN_3472 = 6'h1e == architecturalRegMap_17 ? 1'h0 : _GEN_3344; // @[decode.scala 393:{46,46}]
  wire  _GEN_3473 = 6'h1f == architecturalRegMap_17 ? 1'h0 : _GEN_3345; // @[decode.scala 393:{46,46}]
  wire  _GEN_3474 = 6'h20 == architecturalRegMap_17 ? 1'h0 : _GEN_3346; // @[decode.scala 393:{46,46}]
  wire  _GEN_3475 = 6'h21 == architecturalRegMap_17 ? 1'h0 : _GEN_3347; // @[decode.scala 393:{46,46}]
  wire  _GEN_3476 = 6'h22 == architecturalRegMap_17 ? 1'h0 : _GEN_3348; // @[decode.scala 393:{46,46}]
  wire  _GEN_3477 = 6'h23 == architecturalRegMap_17 ? 1'h0 : _GEN_3349; // @[decode.scala 393:{46,46}]
  wire  _GEN_3478 = 6'h24 == architecturalRegMap_17 ? 1'h0 : _GEN_3350; // @[decode.scala 393:{46,46}]
  wire  _GEN_3479 = 6'h25 == architecturalRegMap_17 ? 1'h0 : _GEN_3351; // @[decode.scala 393:{46,46}]
  wire  _GEN_3480 = 6'h26 == architecturalRegMap_17 ? 1'h0 : _GEN_3352; // @[decode.scala 393:{46,46}]
  wire  _GEN_3481 = 6'h27 == architecturalRegMap_17 ? 1'h0 : _GEN_3353; // @[decode.scala 393:{46,46}]
  wire  _GEN_3482 = 6'h28 == architecturalRegMap_17 ? 1'h0 : _GEN_3354; // @[decode.scala 393:{46,46}]
  wire  _GEN_3483 = 6'h29 == architecturalRegMap_17 ? 1'h0 : _GEN_3355; // @[decode.scala 393:{46,46}]
  wire  _GEN_3484 = 6'h2a == architecturalRegMap_17 ? 1'h0 : _GEN_3356; // @[decode.scala 393:{46,46}]
  wire  _GEN_3485 = 6'h2b == architecturalRegMap_17 ? 1'h0 : _GEN_3357; // @[decode.scala 393:{46,46}]
  wire  _GEN_3486 = 6'h2c == architecturalRegMap_17 ? 1'h0 : _GEN_3358; // @[decode.scala 393:{46,46}]
  wire  _GEN_3487 = 6'h2d == architecturalRegMap_17 ? 1'h0 : _GEN_3359; // @[decode.scala 393:{46,46}]
  wire  _GEN_3488 = 6'h2e == architecturalRegMap_17 ? 1'h0 : _GEN_3360; // @[decode.scala 393:{46,46}]
  wire  _GEN_3489 = 6'h2f == architecturalRegMap_17 ? 1'h0 : _GEN_3361; // @[decode.scala 393:{46,46}]
  wire  _GEN_3490 = 6'h30 == architecturalRegMap_17 ? 1'h0 : _GEN_3362; // @[decode.scala 393:{46,46}]
  wire  _GEN_3491 = 6'h31 == architecturalRegMap_17 ? 1'h0 : _GEN_3363; // @[decode.scala 393:{46,46}]
  wire  _GEN_3492 = 6'h32 == architecturalRegMap_17 ? 1'h0 : _GEN_3364; // @[decode.scala 393:{46,46}]
  wire  _GEN_3493 = 6'h33 == architecturalRegMap_17 ? 1'h0 : _GEN_3365; // @[decode.scala 393:{46,46}]
  wire  _GEN_3494 = 6'h34 == architecturalRegMap_17 ? 1'h0 : _GEN_3366; // @[decode.scala 393:{46,46}]
  wire  _GEN_3495 = 6'h35 == architecturalRegMap_17 ? 1'h0 : _GEN_3367; // @[decode.scala 393:{46,46}]
  wire  _GEN_3496 = 6'h36 == architecturalRegMap_17 ? 1'h0 : _GEN_3368; // @[decode.scala 393:{46,46}]
  wire  _GEN_3497 = 6'h37 == architecturalRegMap_17 ? 1'h0 : _GEN_3369; // @[decode.scala 393:{46,46}]
  wire  _GEN_3498 = 6'h38 == architecturalRegMap_17 ? 1'h0 : _GEN_3370; // @[decode.scala 393:{46,46}]
  wire  _GEN_3499 = 6'h39 == architecturalRegMap_17 ? 1'h0 : _GEN_3371; // @[decode.scala 393:{46,46}]
  wire  _GEN_3500 = 6'h3a == architecturalRegMap_17 ? 1'h0 : _GEN_3372; // @[decode.scala 393:{46,46}]
  wire  _GEN_3501 = 6'h3b == architecturalRegMap_17 ? 1'h0 : _GEN_3373; // @[decode.scala 393:{46,46}]
  wire  _GEN_3502 = 6'h3c == architecturalRegMap_17 ? 1'h0 : _GEN_3374; // @[decode.scala 393:{46,46}]
  wire  _GEN_3503 = 6'h3d == architecturalRegMap_17 ? 1'h0 : _GEN_3375; // @[decode.scala 393:{46,46}]
  wire  _GEN_3504 = 6'h3e == architecturalRegMap_17 ? 1'h0 : _GEN_3376; // @[decode.scala 393:{46,46}]
  wire  _GEN_3570 = 6'h0 == architecturalRegMap_18 ? 1'h0 : _GEN_3442; // @[decode.scala 393:{46,46}]
  wire  _GEN_3571 = 6'h1 == architecturalRegMap_18 ? 1'h0 : _GEN_3443; // @[decode.scala 393:{46,46}]
  wire  _GEN_3572 = 6'h2 == architecturalRegMap_18 ? 1'h0 : _GEN_3444; // @[decode.scala 393:{46,46}]
  wire  _GEN_3573 = 6'h3 == architecturalRegMap_18 ? 1'h0 : _GEN_3445; // @[decode.scala 393:{46,46}]
  wire  _GEN_3574 = 6'h4 == architecturalRegMap_18 ? 1'h0 : _GEN_3446; // @[decode.scala 393:{46,46}]
  wire  _GEN_3575 = 6'h5 == architecturalRegMap_18 ? 1'h0 : _GEN_3447; // @[decode.scala 393:{46,46}]
  wire  _GEN_3576 = 6'h6 == architecturalRegMap_18 ? 1'h0 : _GEN_3448; // @[decode.scala 393:{46,46}]
  wire  _GEN_3577 = 6'h7 == architecturalRegMap_18 ? 1'h0 : _GEN_3449; // @[decode.scala 393:{46,46}]
  wire  _GEN_3578 = 6'h8 == architecturalRegMap_18 ? 1'h0 : _GEN_3450; // @[decode.scala 393:{46,46}]
  wire  _GEN_3579 = 6'h9 == architecturalRegMap_18 ? 1'h0 : _GEN_3451; // @[decode.scala 393:{46,46}]
  wire  _GEN_3580 = 6'ha == architecturalRegMap_18 ? 1'h0 : _GEN_3452; // @[decode.scala 393:{46,46}]
  wire  _GEN_3581 = 6'hb == architecturalRegMap_18 ? 1'h0 : _GEN_3453; // @[decode.scala 393:{46,46}]
  wire  _GEN_3582 = 6'hc == architecturalRegMap_18 ? 1'h0 : _GEN_3454; // @[decode.scala 393:{46,46}]
  wire  _GEN_3583 = 6'hd == architecturalRegMap_18 ? 1'h0 : _GEN_3455; // @[decode.scala 393:{46,46}]
  wire  _GEN_3584 = 6'he == architecturalRegMap_18 ? 1'h0 : _GEN_3456; // @[decode.scala 393:{46,46}]
  wire  _GEN_3585 = 6'hf == architecturalRegMap_18 ? 1'h0 : _GEN_3457; // @[decode.scala 393:{46,46}]
  wire  _GEN_3586 = 6'h10 == architecturalRegMap_18 ? 1'h0 : _GEN_3458; // @[decode.scala 393:{46,46}]
  wire  _GEN_3587 = 6'h11 == architecturalRegMap_18 ? 1'h0 : _GEN_3459; // @[decode.scala 393:{46,46}]
  wire  _GEN_3588 = 6'h12 == architecturalRegMap_18 ? 1'h0 : _GEN_3460; // @[decode.scala 393:{46,46}]
  wire  _GEN_3589 = 6'h13 == architecturalRegMap_18 ? 1'h0 : _GEN_3461; // @[decode.scala 393:{46,46}]
  wire  _GEN_3590 = 6'h14 == architecturalRegMap_18 ? 1'h0 : _GEN_3462; // @[decode.scala 393:{46,46}]
  wire  _GEN_3591 = 6'h15 == architecturalRegMap_18 ? 1'h0 : _GEN_3463; // @[decode.scala 393:{46,46}]
  wire  _GEN_3592 = 6'h16 == architecturalRegMap_18 ? 1'h0 : _GEN_3464; // @[decode.scala 393:{46,46}]
  wire  _GEN_3593 = 6'h17 == architecturalRegMap_18 ? 1'h0 : _GEN_3465; // @[decode.scala 393:{46,46}]
  wire  _GEN_3594 = 6'h18 == architecturalRegMap_18 ? 1'h0 : _GEN_3466; // @[decode.scala 393:{46,46}]
  wire  _GEN_3595 = 6'h19 == architecturalRegMap_18 ? 1'h0 : _GEN_3467; // @[decode.scala 393:{46,46}]
  wire  _GEN_3596 = 6'h1a == architecturalRegMap_18 ? 1'h0 : _GEN_3468; // @[decode.scala 393:{46,46}]
  wire  _GEN_3597 = 6'h1b == architecturalRegMap_18 ? 1'h0 : _GEN_3469; // @[decode.scala 393:{46,46}]
  wire  _GEN_3598 = 6'h1c == architecturalRegMap_18 ? 1'h0 : _GEN_3470; // @[decode.scala 393:{46,46}]
  wire  _GEN_3599 = 6'h1d == architecturalRegMap_18 ? 1'h0 : _GEN_3471; // @[decode.scala 393:{46,46}]
  wire  _GEN_3600 = 6'h1e == architecturalRegMap_18 ? 1'h0 : _GEN_3472; // @[decode.scala 393:{46,46}]
  wire  _GEN_3601 = 6'h1f == architecturalRegMap_18 ? 1'h0 : _GEN_3473; // @[decode.scala 393:{46,46}]
  wire  _GEN_3602 = 6'h20 == architecturalRegMap_18 ? 1'h0 : _GEN_3474; // @[decode.scala 393:{46,46}]
  wire  _GEN_3603 = 6'h21 == architecturalRegMap_18 ? 1'h0 : _GEN_3475; // @[decode.scala 393:{46,46}]
  wire  _GEN_3604 = 6'h22 == architecturalRegMap_18 ? 1'h0 : _GEN_3476; // @[decode.scala 393:{46,46}]
  wire  _GEN_3605 = 6'h23 == architecturalRegMap_18 ? 1'h0 : _GEN_3477; // @[decode.scala 393:{46,46}]
  wire  _GEN_3606 = 6'h24 == architecturalRegMap_18 ? 1'h0 : _GEN_3478; // @[decode.scala 393:{46,46}]
  wire  _GEN_3607 = 6'h25 == architecturalRegMap_18 ? 1'h0 : _GEN_3479; // @[decode.scala 393:{46,46}]
  wire  _GEN_3608 = 6'h26 == architecturalRegMap_18 ? 1'h0 : _GEN_3480; // @[decode.scala 393:{46,46}]
  wire  _GEN_3609 = 6'h27 == architecturalRegMap_18 ? 1'h0 : _GEN_3481; // @[decode.scala 393:{46,46}]
  wire  _GEN_3610 = 6'h28 == architecturalRegMap_18 ? 1'h0 : _GEN_3482; // @[decode.scala 393:{46,46}]
  wire  _GEN_3611 = 6'h29 == architecturalRegMap_18 ? 1'h0 : _GEN_3483; // @[decode.scala 393:{46,46}]
  wire  _GEN_3612 = 6'h2a == architecturalRegMap_18 ? 1'h0 : _GEN_3484; // @[decode.scala 393:{46,46}]
  wire  _GEN_3613 = 6'h2b == architecturalRegMap_18 ? 1'h0 : _GEN_3485; // @[decode.scala 393:{46,46}]
  wire  _GEN_3614 = 6'h2c == architecturalRegMap_18 ? 1'h0 : _GEN_3486; // @[decode.scala 393:{46,46}]
  wire  _GEN_3615 = 6'h2d == architecturalRegMap_18 ? 1'h0 : _GEN_3487; // @[decode.scala 393:{46,46}]
  wire  _GEN_3616 = 6'h2e == architecturalRegMap_18 ? 1'h0 : _GEN_3488; // @[decode.scala 393:{46,46}]
  wire  _GEN_3617 = 6'h2f == architecturalRegMap_18 ? 1'h0 : _GEN_3489; // @[decode.scala 393:{46,46}]
  wire  _GEN_3618 = 6'h30 == architecturalRegMap_18 ? 1'h0 : _GEN_3490; // @[decode.scala 393:{46,46}]
  wire  _GEN_3619 = 6'h31 == architecturalRegMap_18 ? 1'h0 : _GEN_3491; // @[decode.scala 393:{46,46}]
  wire  _GEN_3620 = 6'h32 == architecturalRegMap_18 ? 1'h0 : _GEN_3492; // @[decode.scala 393:{46,46}]
  wire  _GEN_3621 = 6'h33 == architecturalRegMap_18 ? 1'h0 : _GEN_3493; // @[decode.scala 393:{46,46}]
  wire  _GEN_3622 = 6'h34 == architecturalRegMap_18 ? 1'h0 : _GEN_3494; // @[decode.scala 393:{46,46}]
  wire  _GEN_3623 = 6'h35 == architecturalRegMap_18 ? 1'h0 : _GEN_3495; // @[decode.scala 393:{46,46}]
  wire  _GEN_3624 = 6'h36 == architecturalRegMap_18 ? 1'h0 : _GEN_3496; // @[decode.scala 393:{46,46}]
  wire  _GEN_3625 = 6'h37 == architecturalRegMap_18 ? 1'h0 : _GEN_3497; // @[decode.scala 393:{46,46}]
  wire  _GEN_3626 = 6'h38 == architecturalRegMap_18 ? 1'h0 : _GEN_3498; // @[decode.scala 393:{46,46}]
  wire  _GEN_3627 = 6'h39 == architecturalRegMap_18 ? 1'h0 : _GEN_3499; // @[decode.scala 393:{46,46}]
  wire  _GEN_3628 = 6'h3a == architecturalRegMap_18 ? 1'h0 : _GEN_3500; // @[decode.scala 393:{46,46}]
  wire  _GEN_3629 = 6'h3b == architecturalRegMap_18 ? 1'h0 : _GEN_3501; // @[decode.scala 393:{46,46}]
  wire  _GEN_3630 = 6'h3c == architecturalRegMap_18 ? 1'h0 : _GEN_3502; // @[decode.scala 393:{46,46}]
  wire  _GEN_3631 = 6'h3d == architecturalRegMap_18 ? 1'h0 : _GEN_3503; // @[decode.scala 393:{46,46}]
  wire  _GEN_3632 = 6'h3e == architecturalRegMap_18 ? 1'h0 : _GEN_3504; // @[decode.scala 393:{46,46}]
  wire  _GEN_3698 = 6'h0 == architecturalRegMap_19 ? 1'h0 : _GEN_3570; // @[decode.scala 393:{46,46}]
  wire  _GEN_3699 = 6'h1 == architecturalRegMap_19 ? 1'h0 : _GEN_3571; // @[decode.scala 393:{46,46}]
  wire  _GEN_3700 = 6'h2 == architecturalRegMap_19 ? 1'h0 : _GEN_3572; // @[decode.scala 393:{46,46}]
  wire  _GEN_3701 = 6'h3 == architecturalRegMap_19 ? 1'h0 : _GEN_3573; // @[decode.scala 393:{46,46}]
  wire  _GEN_3702 = 6'h4 == architecturalRegMap_19 ? 1'h0 : _GEN_3574; // @[decode.scala 393:{46,46}]
  wire  _GEN_3703 = 6'h5 == architecturalRegMap_19 ? 1'h0 : _GEN_3575; // @[decode.scala 393:{46,46}]
  wire  _GEN_3704 = 6'h6 == architecturalRegMap_19 ? 1'h0 : _GEN_3576; // @[decode.scala 393:{46,46}]
  wire  _GEN_3705 = 6'h7 == architecturalRegMap_19 ? 1'h0 : _GEN_3577; // @[decode.scala 393:{46,46}]
  wire  _GEN_3706 = 6'h8 == architecturalRegMap_19 ? 1'h0 : _GEN_3578; // @[decode.scala 393:{46,46}]
  wire  _GEN_3707 = 6'h9 == architecturalRegMap_19 ? 1'h0 : _GEN_3579; // @[decode.scala 393:{46,46}]
  wire  _GEN_3708 = 6'ha == architecturalRegMap_19 ? 1'h0 : _GEN_3580; // @[decode.scala 393:{46,46}]
  wire  _GEN_3709 = 6'hb == architecturalRegMap_19 ? 1'h0 : _GEN_3581; // @[decode.scala 393:{46,46}]
  wire  _GEN_3710 = 6'hc == architecturalRegMap_19 ? 1'h0 : _GEN_3582; // @[decode.scala 393:{46,46}]
  wire  _GEN_3711 = 6'hd == architecturalRegMap_19 ? 1'h0 : _GEN_3583; // @[decode.scala 393:{46,46}]
  wire  _GEN_3712 = 6'he == architecturalRegMap_19 ? 1'h0 : _GEN_3584; // @[decode.scala 393:{46,46}]
  wire  _GEN_3713 = 6'hf == architecturalRegMap_19 ? 1'h0 : _GEN_3585; // @[decode.scala 393:{46,46}]
  wire  _GEN_3714 = 6'h10 == architecturalRegMap_19 ? 1'h0 : _GEN_3586; // @[decode.scala 393:{46,46}]
  wire  _GEN_3715 = 6'h11 == architecturalRegMap_19 ? 1'h0 : _GEN_3587; // @[decode.scala 393:{46,46}]
  wire  _GEN_3716 = 6'h12 == architecturalRegMap_19 ? 1'h0 : _GEN_3588; // @[decode.scala 393:{46,46}]
  wire  _GEN_3717 = 6'h13 == architecturalRegMap_19 ? 1'h0 : _GEN_3589; // @[decode.scala 393:{46,46}]
  wire  _GEN_3718 = 6'h14 == architecturalRegMap_19 ? 1'h0 : _GEN_3590; // @[decode.scala 393:{46,46}]
  wire  _GEN_3719 = 6'h15 == architecturalRegMap_19 ? 1'h0 : _GEN_3591; // @[decode.scala 393:{46,46}]
  wire  _GEN_3720 = 6'h16 == architecturalRegMap_19 ? 1'h0 : _GEN_3592; // @[decode.scala 393:{46,46}]
  wire  _GEN_3721 = 6'h17 == architecturalRegMap_19 ? 1'h0 : _GEN_3593; // @[decode.scala 393:{46,46}]
  wire  _GEN_3722 = 6'h18 == architecturalRegMap_19 ? 1'h0 : _GEN_3594; // @[decode.scala 393:{46,46}]
  wire  _GEN_3723 = 6'h19 == architecturalRegMap_19 ? 1'h0 : _GEN_3595; // @[decode.scala 393:{46,46}]
  wire  _GEN_3724 = 6'h1a == architecturalRegMap_19 ? 1'h0 : _GEN_3596; // @[decode.scala 393:{46,46}]
  wire  _GEN_3725 = 6'h1b == architecturalRegMap_19 ? 1'h0 : _GEN_3597; // @[decode.scala 393:{46,46}]
  wire  _GEN_3726 = 6'h1c == architecturalRegMap_19 ? 1'h0 : _GEN_3598; // @[decode.scala 393:{46,46}]
  wire  _GEN_3727 = 6'h1d == architecturalRegMap_19 ? 1'h0 : _GEN_3599; // @[decode.scala 393:{46,46}]
  wire  _GEN_3728 = 6'h1e == architecturalRegMap_19 ? 1'h0 : _GEN_3600; // @[decode.scala 393:{46,46}]
  wire  _GEN_3729 = 6'h1f == architecturalRegMap_19 ? 1'h0 : _GEN_3601; // @[decode.scala 393:{46,46}]
  wire  _GEN_3730 = 6'h20 == architecturalRegMap_19 ? 1'h0 : _GEN_3602; // @[decode.scala 393:{46,46}]
  wire  _GEN_3731 = 6'h21 == architecturalRegMap_19 ? 1'h0 : _GEN_3603; // @[decode.scala 393:{46,46}]
  wire  _GEN_3732 = 6'h22 == architecturalRegMap_19 ? 1'h0 : _GEN_3604; // @[decode.scala 393:{46,46}]
  wire  _GEN_3733 = 6'h23 == architecturalRegMap_19 ? 1'h0 : _GEN_3605; // @[decode.scala 393:{46,46}]
  wire  _GEN_3734 = 6'h24 == architecturalRegMap_19 ? 1'h0 : _GEN_3606; // @[decode.scala 393:{46,46}]
  wire  _GEN_3735 = 6'h25 == architecturalRegMap_19 ? 1'h0 : _GEN_3607; // @[decode.scala 393:{46,46}]
  wire  _GEN_3736 = 6'h26 == architecturalRegMap_19 ? 1'h0 : _GEN_3608; // @[decode.scala 393:{46,46}]
  wire  _GEN_3737 = 6'h27 == architecturalRegMap_19 ? 1'h0 : _GEN_3609; // @[decode.scala 393:{46,46}]
  wire  _GEN_3738 = 6'h28 == architecturalRegMap_19 ? 1'h0 : _GEN_3610; // @[decode.scala 393:{46,46}]
  wire  _GEN_3739 = 6'h29 == architecturalRegMap_19 ? 1'h0 : _GEN_3611; // @[decode.scala 393:{46,46}]
  wire  _GEN_3740 = 6'h2a == architecturalRegMap_19 ? 1'h0 : _GEN_3612; // @[decode.scala 393:{46,46}]
  wire  _GEN_3741 = 6'h2b == architecturalRegMap_19 ? 1'h0 : _GEN_3613; // @[decode.scala 393:{46,46}]
  wire  _GEN_3742 = 6'h2c == architecturalRegMap_19 ? 1'h0 : _GEN_3614; // @[decode.scala 393:{46,46}]
  wire  _GEN_3743 = 6'h2d == architecturalRegMap_19 ? 1'h0 : _GEN_3615; // @[decode.scala 393:{46,46}]
  wire  _GEN_3744 = 6'h2e == architecturalRegMap_19 ? 1'h0 : _GEN_3616; // @[decode.scala 393:{46,46}]
  wire  _GEN_3745 = 6'h2f == architecturalRegMap_19 ? 1'h0 : _GEN_3617; // @[decode.scala 393:{46,46}]
  wire  _GEN_3746 = 6'h30 == architecturalRegMap_19 ? 1'h0 : _GEN_3618; // @[decode.scala 393:{46,46}]
  wire  _GEN_3747 = 6'h31 == architecturalRegMap_19 ? 1'h0 : _GEN_3619; // @[decode.scala 393:{46,46}]
  wire  _GEN_3748 = 6'h32 == architecturalRegMap_19 ? 1'h0 : _GEN_3620; // @[decode.scala 393:{46,46}]
  wire  _GEN_3749 = 6'h33 == architecturalRegMap_19 ? 1'h0 : _GEN_3621; // @[decode.scala 393:{46,46}]
  wire  _GEN_3750 = 6'h34 == architecturalRegMap_19 ? 1'h0 : _GEN_3622; // @[decode.scala 393:{46,46}]
  wire  _GEN_3751 = 6'h35 == architecturalRegMap_19 ? 1'h0 : _GEN_3623; // @[decode.scala 393:{46,46}]
  wire  _GEN_3752 = 6'h36 == architecturalRegMap_19 ? 1'h0 : _GEN_3624; // @[decode.scala 393:{46,46}]
  wire  _GEN_3753 = 6'h37 == architecturalRegMap_19 ? 1'h0 : _GEN_3625; // @[decode.scala 393:{46,46}]
  wire  _GEN_3754 = 6'h38 == architecturalRegMap_19 ? 1'h0 : _GEN_3626; // @[decode.scala 393:{46,46}]
  wire  _GEN_3755 = 6'h39 == architecturalRegMap_19 ? 1'h0 : _GEN_3627; // @[decode.scala 393:{46,46}]
  wire  _GEN_3756 = 6'h3a == architecturalRegMap_19 ? 1'h0 : _GEN_3628; // @[decode.scala 393:{46,46}]
  wire  _GEN_3757 = 6'h3b == architecturalRegMap_19 ? 1'h0 : _GEN_3629; // @[decode.scala 393:{46,46}]
  wire  _GEN_3758 = 6'h3c == architecturalRegMap_19 ? 1'h0 : _GEN_3630; // @[decode.scala 393:{46,46}]
  wire  _GEN_3759 = 6'h3d == architecturalRegMap_19 ? 1'h0 : _GEN_3631; // @[decode.scala 393:{46,46}]
  wire  _GEN_3760 = 6'h3e == architecturalRegMap_19 ? 1'h0 : _GEN_3632; // @[decode.scala 393:{46,46}]
  wire  _GEN_3826 = 6'h0 == architecturalRegMap_20 ? 1'h0 : _GEN_3698; // @[decode.scala 393:{46,46}]
  wire  _GEN_3827 = 6'h1 == architecturalRegMap_20 ? 1'h0 : _GEN_3699; // @[decode.scala 393:{46,46}]
  wire  _GEN_3828 = 6'h2 == architecturalRegMap_20 ? 1'h0 : _GEN_3700; // @[decode.scala 393:{46,46}]
  wire  _GEN_3829 = 6'h3 == architecturalRegMap_20 ? 1'h0 : _GEN_3701; // @[decode.scala 393:{46,46}]
  wire  _GEN_3830 = 6'h4 == architecturalRegMap_20 ? 1'h0 : _GEN_3702; // @[decode.scala 393:{46,46}]
  wire  _GEN_3831 = 6'h5 == architecturalRegMap_20 ? 1'h0 : _GEN_3703; // @[decode.scala 393:{46,46}]
  wire  _GEN_3832 = 6'h6 == architecturalRegMap_20 ? 1'h0 : _GEN_3704; // @[decode.scala 393:{46,46}]
  wire  _GEN_3833 = 6'h7 == architecturalRegMap_20 ? 1'h0 : _GEN_3705; // @[decode.scala 393:{46,46}]
  wire  _GEN_3834 = 6'h8 == architecturalRegMap_20 ? 1'h0 : _GEN_3706; // @[decode.scala 393:{46,46}]
  wire  _GEN_3835 = 6'h9 == architecturalRegMap_20 ? 1'h0 : _GEN_3707; // @[decode.scala 393:{46,46}]
  wire  _GEN_3836 = 6'ha == architecturalRegMap_20 ? 1'h0 : _GEN_3708; // @[decode.scala 393:{46,46}]
  wire  _GEN_3837 = 6'hb == architecturalRegMap_20 ? 1'h0 : _GEN_3709; // @[decode.scala 393:{46,46}]
  wire  _GEN_3838 = 6'hc == architecturalRegMap_20 ? 1'h0 : _GEN_3710; // @[decode.scala 393:{46,46}]
  wire  _GEN_3839 = 6'hd == architecturalRegMap_20 ? 1'h0 : _GEN_3711; // @[decode.scala 393:{46,46}]
  wire  _GEN_3840 = 6'he == architecturalRegMap_20 ? 1'h0 : _GEN_3712; // @[decode.scala 393:{46,46}]
  wire  _GEN_3841 = 6'hf == architecturalRegMap_20 ? 1'h0 : _GEN_3713; // @[decode.scala 393:{46,46}]
  wire  _GEN_3842 = 6'h10 == architecturalRegMap_20 ? 1'h0 : _GEN_3714; // @[decode.scala 393:{46,46}]
  wire  _GEN_3843 = 6'h11 == architecturalRegMap_20 ? 1'h0 : _GEN_3715; // @[decode.scala 393:{46,46}]
  wire  _GEN_3844 = 6'h12 == architecturalRegMap_20 ? 1'h0 : _GEN_3716; // @[decode.scala 393:{46,46}]
  wire  _GEN_3845 = 6'h13 == architecturalRegMap_20 ? 1'h0 : _GEN_3717; // @[decode.scala 393:{46,46}]
  wire  _GEN_3846 = 6'h14 == architecturalRegMap_20 ? 1'h0 : _GEN_3718; // @[decode.scala 393:{46,46}]
  wire  _GEN_3847 = 6'h15 == architecturalRegMap_20 ? 1'h0 : _GEN_3719; // @[decode.scala 393:{46,46}]
  wire  _GEN_3848 = 6'h16 == architecturalRegMap_20 ? 1'h0 : _GEN_3720; // @[decode.scala 393:{46,46}]
  wire  _GEN_3849 = 6'h17 == architecturalRegMap_20 ? 1'h0 : _GEN_3721; // @[decode.scala 393:{46,46}]
  wire  _GEN_3850 = 6'h18 == architecturalRegMap_20 ? 1'h0 : _GEN_3722; // @[decode.scala 393:{46,46}]
  wire  _GEN_3851 = 6'h19 == architecturalRegMap_20 ? 1'h0 : _GEN_3723; // @[decode.scala 393:{46,46}]
  wire  _GEN_3852 = 6'h1a == architecturalRegMap_20 ? 1'h0 : _GEN_3724; // @[decode.scala 393:{46,46}]
  wire  _GEN_3853 = 6'h1b == architecturalRegMap_20 ? 1'h0 : _GEN_3725; // @[decode.scala 393:{46,46}]
  wire  _GEN_3854 = 6'h1c == architecturalRegMap_20 ? 1'h0 : _GEN_3726; // @[decode.scala 393:{46,46}]
  wire  _GEN_3855 = 6'h1d == architecturalRegMap_20 ? 1'h0 : _GEN_3727; // @[decode.scala 393:{46,46}]
  wire  _GEN_3856 = 6'h1e == architecturalRegMap_20 ? 1'h0 : _GEN_3728; // @[decode.scala 393:{46,46}]
  wire  _GEN_3857 = 6'h1f == architecturalRegMap_20 ? 1'h0 : _GEN_3729; // @[decode.scala 393:{46,46}]
  wire  _GEN_3858 = 6'h20 == architecturalRegMap_20 ? 1'h0 : _GEN_3730; // @[decode.scala 393:{46,46}]
  wire  _GEN_3859 = 6'h21 == architecturalRegMap_20 ? 1'h0 : _GEN_3731; // @[decode.scala 393:{46,46}]
  wire  _GEN_3860 = 6'h22 == architecturalRegMap_20 ? 1'h0 : _GEN_3732; // @[decode.scala 393:{46,46}]
  wire  _GEN_3861 = 6'h23 == architecturalRegMap_20 ? 1'h0 : _GEN_3733; // @[decode.scala 393:{46,46}]
  wire  _GEN_3862 = 6'h24 == architecturalRegMap_20 ? 1'h0 : _GEN_3734; // @[decode.scala 393:{46,46}]
  wire  _GEN_3863 = 6'h25 == architecturalRegMap_20 ? 1'h0 : _GEN_3735; // @[decode.scala 393:{46,46}]
  wire  _GEN_3864 = 6'h26 == architecturalRegMap_20 ? 1'h0 : _GEN_3736; // @[decode.scala 393:{46,46}]
  wire  _GEN_3865 = 6'h27 == architecturalRegMap_20 ? 1'h0 : _GEN_3737; // @[decode.scala 393:{46,46}]
  wire  _GEN_3866 = 6'h28 == architecturalRegMap_20 ? 1'h0 : _GEN_3738; // @[decode.scala 393:{46,46}]
  wire  _GEN_3867 = 6'h29 == architecturalRegMap_20 ? 1'h0 : _GEN_3739; // @[decode.scala 393:{46,46}]
  wire  _GEN_3868 = 6'h2a == architecturalRegMap_20 ? 1'h0 : _GEN_3740; // @[decode.scala 393:{46,46}]
  wire  _GEN_3869 = 6'h2b == architecturalRegMap_20 ? 1'h0 : _GEN_3741; // @[decode.scala 393:{46,46}]
  wire  _GEN_3870 = 6'h2c == architecturalRegMap_20 ? 1'h0 : _GEN_3742; // @[decode.scala 393:{46,46}]
  wire  _GEN_3871 = 6'h2d == architecturalRegMap_20 ? 1'h0 : _GEN_3743; // @[decode.scala 393:{46,46}]
  wire  _GEN_3872 = 6'h2e == architecturalRegMap_20 ? 1'h0 : _GEN_3744; // @[decode.scala 393:{46,46}]
  wire  _GEN_3873 = 6'h2f == architecturalRegMap_20 ? 1'h0 : _GEN_3745; // @[decode.scala 393:{46,46}]
  wire  _GEN_3874 = 6'h30 == architecturalRegMap_20 ? 1'h0 : _GEN_3746; // @[decode.scala 393:{46,46}]
  wire  _GEN_3875 = 6'h31 == architecturalRegMap_20 ? 1'h0 : _GEN_3747; // @[decode.scala 393:{46,46}]
  wire  _GEN_3876 = 6'h32 == architecturalRegMap_20 ? 1'h0 : _GEN_3748; // @[decode.scala 393:{46,46}]
  wire  _GEN_3877 = 6'h33 == architecturalRegMap_20 ? 1'h0 : _GEN_3749; // @[decode.scala 393:{46,46}]
  wire  _GEN_3878 = 6'h34 == architecturalRegMap_20 ? 1'h0 : _GEN_3750; // @[decode.scala 393:{46,46}]
  wire  _GEN_3879 = 6'h35 == architecturalRegMap_20 ? 1'h0 : _GEN_3751; // @[decode.scala 393:{46,46}]
  wire  _GEN_3880 = 6'h36 == architecturalRegMap_20 ? 1'h0 : _GEN_3752; // @[decode.scala 393:{46,46}]
  wire  _GEN_3881 = 6'h37 == architecturalRegMap_20 ? 1'h0 : _GEN_3753; // @[decode.scala 393:{46,46}]
  wire  _GEN_3882 = 6'h38 == architecturalRegMap_20 ? 1'h0 : _GEN_3754; // @[decode.scala 393:{46,46}]
  wire  _GEN_3883 = 6'h39 == architecturalRegMap_20 ? 1'h0 : _GEN_3755; // @[decode.scala 393:{46,46}]
  wire  _GEN_3884 = 6'h3a == architecturalRegMap_20 ? 1'h0 : _GEN_3756; // @[decode.scala 393:{46,46}]
  wire  _GEN_3885 = 6'h3b == architecturalRegMap_20 ? 1'h0 : _GEN_3757; // @[decode.scala 393:{46,46}]
  wire  _GEN_3886 = 6'h3c == architecturalRegMap_20 ? 1'h0 : _GEN_3758; // @[decode.scala 393:{46,46}]
  wire  _GEN_3887 = 6'h3d == architecturalRegMap_20 ? 1'h0 : _GEN_3759; // @[decode.scala 393:{46,46}]
  wire  _GEN_3888 = 6'h3e == architecturalRegMap_20 ? 1'h0 : _GEN_3760; // @[decode.scala 393:{46,46}]
  wire  _GEN_3954 = 6'h0 == architecturalRegMap_21 ? 1'h0 : _GEN_3826; // @[decode.scala 393:{46,46}]
  wire  _GEN_3955 = 6'h1 == architecturalRegMap_21 ? 1'h0 : _GEN_3827; // @[decode.scala 393:{46,46}]
  wire  _GEN_3956 = 6'h2 == architecturalRegMap_21 ? 1'h0 : _GEN_3828; // @[decode.scala 393:{46,46}]
  wire  _GEN_3957 = 6'h3 == architecturalRegMap_21 ? 1'h0 : _GEN_3829; // @[decode.scala 393:{46,46}]
  wire  _GEN_3958 = 6'h4 == architecturalRegMap_21 ? 1'h0 : _GEN_3830; // @[decode.scala 393:{46,46}]
  wire  _GEN_3959 = 6'h5 == architecturalRegMap_21 ? 1'h0 : _GEN_3831; // @[decode.scala 393:{46,46}]
  wire  _GEN_3960 = 6'h6 == architecturalRegMap_21 ? 1'h0 : _GEN_3832; // @[decode.scala 393:{46,46}]
  wire  _GEN_3961 = 6'h7 == architecturalRegMap_21 ? 1'h0 : _GEN_3833; // @[decode.scala 393:{46,46}]
  wire  _GEN_3962 = 6'h8 == architecturalRegMap_21 ? 1'h0 : _GEN_3834; // @[decode.scala 393:{46,46}]
  wire  _GEN_3963 = 6'h9 == architecturalRegMap_21 ? 1'h0 : _GEN_3835; // @[decode.scala 393:{46,46}]
  wire  _GEN_3964 = 6'ha == architecturalRegMap_21 ? 1'h0 : _GEN_3836; // @[decode.scala 393:{46,46}]
  wire  _GEN_3965 = 6'hb == architecturalRegMap_21 ? 1'h0 : _GEN_3837; // @[decode.scala 393:{46,46}]
  wire  _GEN_3966 = 6'hc == architecturalRegMap_21 ? 1'h0 : _GEN_3838; // @[decode.scala 393:{46,46}]
  wire  _GEN_3967 = 6'hd == architecturalRegMap_21 ? 1'h0 : _GEN_3839; // @[decode.scala 393:{46,46}]
  wire  _GEN_3968 = 6'he == architecturalRegMap_21 ? 1'h0 : _GEN_3840; // @[decode.scala 393:{46,46}]
  wire  _GEN_3969 = 6'hf == architecturalRegMap_21 ? 1'h0 : _GEN_3841; // @[decode.scala 393:{46,46}]
  wire  _GEN_3970 = 6'h10 == architecturalRegMap_21 ? 1'h0 : _GEN_3842; // @[decode.scala 393:{46,46}]
  wire  _GEN_3971 = 6'h11 == architecturalRegMap_21 ? 1'h0 : _GEN_3843; // @[decode.scala 393:{46,46}]
  wire  _GEN_3972 = 6'h12 == architecturalRegMap_21 ? 1'h0 : _GEN_3844; // @[decode.scala 393:{46,46}]
  wire  _GEN_3973 = 6'h13 == architecturalRegMap_21 ? 1'h0 : _GEN_3845; // @[decode.scala 393:{46,46}]
  wire  _GEN_3974 = 6'h14 == architecturalRegMap_21 ? 1'h0 : _GEN_3846; // @[decode.scala 393:{46,46}]
  wire  _GEN_3975 = 6'h15 == architecturalRegMap_21 ? 1'h0 : _GEN_3847; // @[decode.scala 393:{46,46}]
  wire  _GEN_3976 = 6'h16 == architecturalRegMap_21 ? 1'h0 : _GEN_3848; // @[decode.scala 393:{46,46}]
  wire  _GEN_3977 = 6'h17 == architecturalRegMap_21 ? 1'h0 : _GEN_3849; // @[decode.scala 393:{46,46}]
  wire  _GEN_3978 = 6'h18 == architecturalRegMap_21 ? 1'h0 : _GEN_3850; // @[decode.scala 393:{46,46}]
  wire  _GEN_3979 = 6'h19 == architecturalRegMap_21 ? 1'h0 : _GEN_3851; // @[decode.scala 393:{46,46}]
  wire  _GEN_3980 = 6'h1a == architecturalRegMap_21 ? 1'h0 : _GEN_3852; // @[decode.scala 393:{46,46}]
  wire  _GEN_3981 = 6'h1b == architecturalRegMap_21 ? 1'h0 : _GEN_3853; // @[decode.scala 393:{46,46}]
  wire  _GEN_3982 = 6'h1c == architecturalRegMap_21 ? 1'h0 : _GEN_3854; // @[decode.scala 393:{46,46}]
  wire  _GEN_3983 = 6'h1d == architecturalRegMap_21 ? 1'h0 : _GEN_3855; // @[decode.scala 393:{46,46}]
  wire  _GEN_3984 = 6'h1e == architecturalRegMap_21 ? 1'h0 : _GEN_3856; // @[decode.scala 393:{46,46}]
  wire  _GEN_3985 = 6'h1f == architecturalRegMap_21 ? 1'h0 : _GEN_3857; // @[decode.scala 393:{46,46}]
  wire  _GEN_3986 = 6'h20 == architecturalRegMap_21 ? 1'h0 : _GEN_3858; // @[decode.scala 393:{46,46}]
  wire  _GEN_3987 = 6'h21 == architecturalRegMap_21 ? 1'h0 : _GEN_3859; // @[decode.scala 393:{46,46}]
  wire  _GEN_3988 = 6'h22 == architecturalRegMap_21 ? 1'h0 : _GEN_3860; // @[decode.scala 393:{46,46}]
  wire  _GEN_3989 = 6'h23 == architecturalRegMap_21 ? 1'h0 : _GEN_3861; // @[decode.scala 393:{46,46}]
  wire  _GEN_3990 = 6'h24 == architecturalRegMap_21 ? 1'h0 : _GEN_3862; // @[decode.scala 393:{46,46}]
  wire  _GEN_3991 = 6'h25 == architecturalRegMap_21 ? 1'h0 : _GEN_3863; // @[decode.scala 393:{46,46}]
  wire  _GEN_3992 = 6'h26 == architecturalRegMap_21 ? 1'h0 : _GEN_3864; // @[decode.scala 393:{46,46}]
  wire  _GEN_3993 = 6'h27 == architecturalRegMap_21 ? 1'h0 : _GEN_3865; // @[decode.scala 393:{46,46}]
  wire  _GEN_3994 = 6'h28 == architecturalRegMap_21 ? 1'h0 : _GEN_3866; // @[decode.scala 393:{46,46}]
  wire  _GEN_3995 = 6'h29 == architecturalRegMap_21 ? 1'h0 : _GEN_3867; // @[decode.scala 393:{46,46}]
  wire  _GEN_3996 = 6'h2a == architecturalRegMap_21 ? 1'h0 : _GEN_3868; // @[decode.scala 393:{46,46}]
  wire  _GEN_3997 = 6'h2b == architecturalRegMap_21 ? 1'h0 : _GEN_3869; // @[decode.scala 393:{46,46}]
  wire  _GEN_3998 = 6'h2c == architecturalRegMap_21 ? 1'h0 : _GEN_3870; // @[decode.scala 393:{46,46}]
  wire  _GEN_3999 = 6'h2d == architecturalRegMap_21 ? 1'h0 : _GEN_3871; // @[decode.scala 393:{46,46}]
  wire  _GEN_4000 = 6'h2e == architecturalRegMap_21 ? 1'h0 : _GEN_3872; // @[decode.scala 393:{46,46}]
  wire  _GEN_4001 = 6'h2f == architecturalRegMap_21 ? 1'h0 : _GEN_3873; // @[decode.scala 393:{46,46}]
  wire  _GEN_4002 = 6'h30 == architecturalRegMap_21 ? 1'h0 : _GEN_3874; // @[decode.scala 393:{46,46}]
  wire  _GEN_4003 = 6'h31 == architecturalRegMap_21 ? 1'h0 : _GEN_3875; // @[decode.scala 393:{46,46}]
  wire  _GEN_4004 = 6'h32 == architecturalRegMap_21 ? 1'h0 : _GEN_3876; // @[decode.scala 393:{46,46}]
  wire  _GEN_4005 = 6'h33 == architecturalRegMap_21 ? 1'h0 : _GEN_3877; // @[decode.scala 393:{46,46}]
  wire  _GEN_4006 = 6'h34 == architecturalRegMap_21 ? 1'h0 : _GEN_3878; // @[decode.scala 393:{46,46}]
  wire  _GEN_4007 = 6'h35 == architecturalRegMap_21 ? 1'h0 : _GEN_3879; // @[decode.scala 393:{46,46}]
  wire  _GEN_4008 = 6'h36 == architecturalRegMap_21 ? 1'h0 : _GEN_3880; // @[decode.scala 393:{46,46}]
  wire  _GEN_4009 = 6'h37 == architecturalRegMap_21 ? 1'h0 : _GEN_3881; // @[decode.scala 393:{46,46}]
  wire  _GEN_4010 = 6'h38 == architecturalRegMap_21 ? 1'h0 : _GEN_3882; // @[decode.scala 393:{46,46}]
  wire  _GEN_4011 = 6'h39 == architecturalRegMap_21 ? 1'h0 : _GEN_3883; // @[decode.scala 393:{46,46}]
  wire  _GEN_4012 = 6'h3a == architecturalRegMap_21 ? 1'h0 : _GEN_3884; // @[decode.scala 393:{46,46}]
  wire  _GEN_4013 = 6'h3b == architecturalRegMap_21 ? 1'h0 : _GEN_3885; // @[decode.scala 393:{46,46}]
  wire  _GEN_4014 = 6'h3c == architecturalRegMap_21 ? 1'h0 : _GEN_3886; // @[decode.scala 393:{46,46}]
  wire  _GEN_4015 = 6'h3d == architecturalRegMap_21 ? 1'h0 : _GEN_3887; // @[decode.scala 393:{46,46}]
  wire  _GEN_4016 = 6'h3e == architecturalRegMap_21 ? 1'h0 : _GEN_3888; // @[decode.scala 393:{46,46}]
  wire  _GEN_4082 = 6'h0 == architecturalRegMap_22 ? 1'h0 : _GEN_3954; // @[decode.scala 393:{46,46}]
  wire  _GEN_4083 = 6'h1 == architecturalRegMap_22 ? 1'h0 : _GEN_3955; // @[decode.scala 393:{46,46}]
  wire  _GEN_4084 = 6'h2 == architecturalRegMap_22 ? 1'h0 : _GEN_3956; // @[decode.scala 393:{46,46}]
  wire  _GEN_4085 = 6'h3 == architecturalRegMap_22 ? 1'h0 : _GEN_3957; // @[decode.scala 393:{46,46}]
  wire  _GEN_4086 = 6'h4 == architecturalRegMap_22 ? 1'h0 : _GEN_3958; // @[decode.scala 393:{46,46}]
  wire  _GEN_4087 = 6'h5 == architecturalRegMap_22 ? 1'h0 : _GEN_3959; // @[decode.scala 393:{46,46}]
  wire  _GEN_4088 = 6'h6 == architecturalRegMap_22 ? 1'h0 : _GEN_3960; // @[decode.scala 393:{46,46}]
  wire  _GEN_4089 = 6'h7 == architecturalRegMap_22 ? 1'h0 : _GEN_3961; // @[decode.scala 393:{46,46}]
  wire  _GEN_4090 = 6'h8 == architecturalRegMap_22 ? 1'h0 : _GEN_3962; // @[decode.scala 393:{46,46}]
  wire  _GEN_4091 = 6'h9 == architecturalRegMap_22 ? 1'h0 : _GEN_3963; // @[decode.scala 393:{46,46}]
  wire  _GEN_4092 = 6'ha == architecturalRegMap_22 ? 1'h0 : _GEN_3964; // @[decode.scala 393:{46,46}]
  wire  _GEN_4093 = 6'hb == architecturalRegMap_22 ? 1'h0 : _GEN_3965; // @[decode.scala 393:{46,46}]
  wire  _GEN_4094 = 6'hc == architecturalRegMap_22 ? 1'h0 : _GEN_3966; // @[decode.scala 393:{46,46}]
  wire  _GEN_4095 = 6'hd == architecturalRegMap_22 ? 1'h0 : _GEN_3967; // @[decode.scala 393:{46,46}]
  wire  _GEN_4096 = 6'he == architecturalRegMap_22 ? 1'h0 : _GEN_3968; // @[decode.scala 393:{46,46}]
  wire  _GEN_4097 = 6'hf == architecturalRegMap_22 ? 1'h0 : _GEN_3969; // @[decode.scala 393:{46,46}]
  wire  _GEN_4098 = 6'h10 == architecturalRegMap_22 ? 1'h0 : _GEN_3970; // @[decode.scala 393:{46,46}]
  wire  _GEN_4099 = 6'h11 == architecturalRegMap_22 ? 1'h0 : _GEN_3971; // @[decode.scala 393:{46,46}]
  wire  _GEN_4100 = 6'h12 == architecturalRegMap_22 ? 1'h0 : _GEN_3972; // @[decode.scala 393:{46,46}]
  wire  _GEN_4101 = 6'h13 == architecturalRegMap_22 ? 1'h0 : _GEN_3973; // @[decode.scala 393:{46,46}]
  wire  _GEN_4102 = 6'h14 == architecturalRegMap_22 ? 1'h0 : _GEN_3974; // @[decode.scala 393:{46,46}]
  wire  _GEN_4103 = 6'h15 == architecturalRegMap_22 ? 1'h0 : _GEN_3975; // @[decode.scala 393:{46,46}]
  wire  _GEN_4104 = 6'h16 == architecturalRegMap_22 ? 1'h0 : _GEN_3976; // @[decode.scala 393:{46,46}]
  wire  _GEN_4105 = 6'h17 == architecturalRegMap_22 ? 1'h0 : _GEN_3977; // @[decode.scala 393:{46,46}]
  wire  _GEN_4106 = 6'h18 == architecturalRegMap_22 ? 1'h0 : _GEN_3978; // @[decode.scala 393:{46,46}]
  wire  _GEN_4107 = 6'h19 == architecturalRegMap_22 ? 1'h0 : _GEN_3979; // @[decode.scala 393:{46,46}]
  wire  _GEN_4108 = 6'h1a == architecturalRegMap_22 ? 1'h0 : _GEN_3980; // @[decode.scala 393:{46,46}]
  wire  _GEN_4109 = 6'h1b == architecturalRegMap_22 ? 1'h0 : _GEN_3981; // @[decode.scala 393:{46,46}]
  wire  _GEN_4110 = 6'h1c == architecturalRegMap_22 ? 1'h0 : _GEN_3982; // @[decode.scala 393:{46,46}]
  wire  _GEN_4111 = 6'h1d == architecturalRegMap_22 ? 1'h0 : _GEN_3983; // @[decode.scala 393:{46,46}]
  wire  _GEN_4112 = 6'h1e == architecturalRegMap_22 ? 1'h0 : _GEN_3984; // @[decode.scala 393:{46,46}]
  wire  _GEN_4113 = 6'h1f == architecturalRegMap_22 ? 1'h0 : _GEN_3985; // @[decode.scala 393:{46,46}]
  wire  _GEN_4114 = 6'h20 == architecturalRegMap_22 ? 1'h0 : _GEN_3986; // @[decode.scala 393:{46,46}]
  wire  _GEN_4115 = 6'h21 == architecturalRegMap_22 ? 1'h0 : _GEN_3987; // @[decode.scala 393:{46,46}]
  wire  _GEN_4116 = 6'h22 == architecturalRegMap_22 ? 1'h0 : _GEN_3988; // @[decode.scala 393:{46,46}]
  wire  _GEN_4117 = 6'h23 == architecturalRegMap_22 ? 1'h0 : _GEN_3989; // @[decode.scala 393:{46,46}]
  wire  _GEN_4118 = 6'h24 == architecturalRegMap_22 ? 1'h0 : _GEN_3990; // @[decode.scala 393:{46,46}]
  wire  _GEN_4119 = 6'h25 == architecturalRegMap_22 ? 1'h0 : _GEN_3991; // @[decode.scala 393:{46,46}]
  wire  _GEN_4120 = 6'h26 == architecturalRegMap_22 ? 1'h0 : _GEN_3992; // @[decode.scala 393:{46,46}]
  wire  _GEN_4121 = 6'h27 == architecturalRegMap_22 ? 1'h0 : _GEN_3993; // @[decode.scala 393:{46,46}]
  wire  _GEN_4122 = 6'h28 == architecturalRegMap_22 ? 1'h0 : _GEN_3994; // @[decode.scala 393:{46,46}]
  wire  _GEN_4123 = 6'h29 == architecturalRegMap_22 ? 1'h0 : _GEN_3995; // @[decode.scala 393:{46,46}]
  wire  _GEN_4124 = 6'h2a == architecturalRegMap_22 ? 1'h0 : _GEN_3996; // @[decode.scala 393:{46,46}]
  wire  _GEN_4125 = 6'h2b == architecturalRegMap_22 ? 1'h0 : _GEN_3997; // @[decode.scala 393:{46,46}]
  wire  _GEN_4126 = 6'h2c == architecturalRegMap_22 ? 1'h0 : _GEN_3998; // @[decode.scala 393:{46,46}]
  wire  _GEN_4127 = 6'h2d == architecturalRegMap_22 ? 1'h0 : _GEN_3999; // @[decode.scala 393:{46,46}]
  wire  _GEN_4128 = 6'h2e == architecturalRegMap_22 ? 1'h0 : _GEN_4000; // @[decode.scala 393:{46,46}]
  wire  _GEN_4129 = 6'h2f == architecturalRegMap_22 ? 1'h0 : _GEN_4001; // @[decode.scala 393:{46,46}]
  wire  _GEN_4130 = 6'h30 == architecturalRegMap_22 ? 1'h0 : _GEN_4002; // @[decode.scala 393:{46,46}]
  wire  _GEN_4131 = 6'h31 == architecturalRegMap_22 ? 1'h0 : _GEN_4003; // @[decode.scala 393:{46,46}]
  wire  _GEN_4132 = 6'h32 == architecturalRegMap_22 ? 1'h0 : _GEN_4004; // @[decode.scala 393:{46,46}]
  wire  _GEN_4133 = 6'h33 == architecturalRegMap_22 ? 1'h0 : _GEN_4005; // @[decode.scala 393:{46,46}]
  wire  _GEN_4134 = 6'h34 == architecturalRegMap_22 ? 1'h0 : _GEN_4006; // @[decode.scala 393:{46,46}]
  wire  _GEN_4135 = 6'h35 == architecturalRegMap_22 ? 1'h0 : _GEN_4007; // @[decode.scala 393:{46,46}]
  wire  _GEN_4136 = 6'h36 == architecturalRegMap_22 ? 1'h0 : _GEN_4008; // @[decode.scala 393:{46,46}]
  wire  _GEN_4137 = 6'h37 == architecturalRegMap_22 ? 1'h0 : _GEN_4009; // @[decode.scala 393:{46,46}]
  wire  _GEN_4138 = 6'h38 == architecturalRegMap_22 ? 1'h0 : _GEN_4010; // @[decode.scala 393:{46,46}]
  wire  _GEN_4139 = 6'h39 == architecturalRegMap_22 ? 1'h0 : _GEN_4011; // @[decode.scala 393:{46,46}]
  wire  _GEN_4140 = 6'h3a == architecturalRegMap_22 ? 1'h0 : _GEN_4012; // @[decode.scala 393:{46,46}]
  wire  _GEN_4141 = 6'h3b == architecturalRegMap_22 ? 1'h0 : _GEN_4013; // @[decode.scala 393:{46,46}]
  wire  _GEN_4142 = 6'h3c == architecturalRegMap_22 ? 1'h0 : _GEN_4014; // @[decode.scala 393:{46,46}]
  wire  _GEN_4143 = 6'h3d == architecturalRegMap_22 ? 1'h0 : _GEN_4015; // @[decode.scala 393:{46,46}]
  wire  _GEN_4144 = 6'h3e == architecturalRegMap_22 ? 1'h0 : _GEN_4016; // @[decode.scala 393:{46,46}]
  wire  _GEN_4210 = 6'h0 == architecturalRegMap_23 ? 1'h0 : _GEN_4082; // @[decode.scala 393:{46,46}]
  wire  _GEN_4211 = 6'h1 == architecturalRegMap_23 ? 1'h0 : _GEN_4083; // @[decode.scala 393:{46,46}]
  wire  _GEN_4212 = 6'h2 == architecturalRegMap_23 ? 1'h0 : _GEN_4084; // @[decode.scala 393:{46,46}]
  wire  _GEN_4213 = 6'h3 == architecturalRegMap_23 ? 1'h0 : _GEN_4085; // @[decode.scala 393:{46,46}]
  wire  _GEN_4214 = 6'h4 == architecturalRegMap_23 ? 1'h0 : _GEN_4086; // @[decode.scala 393:{46,46}]
  wire  _GEN_4215 = 6'h5 == architecturalRegMap_23 ? 1'h0 : _GEN_4087; // @[decode.scala 393:{46,46}]
  wire  _GEN_4216 = 6'h6 == architecturalRegMap_23 ? 1'h0 : _GEN_4088; // @[decode.scala 393:{46,46}]
  wire  _GEN_4217 = 6'h7 == architecturalRegMap_23 ? 1'h0 : _GEN_4089; // @[decode.scala 393:{46,46}]
  wire  _GEN_4218 = 6'h8 == architecturalRegMap_23 ? 1'h0 : _GEN_4090; // @[decode.scala 393:{46,46}]
  wire  _GEN_4219 = 6'h9 == architecturalRegMap_23 ? 1'h0 : _GEN_4091; // @[decode.scala 393:{46,46}]
  wire  _GEN_4220 = 6'ha == architecturalRegMap_23 ? 1'h0 : _GEN_4092; // @[decode.scala 393:{46,46}]
  wire  _GEN_4221 = 6'hb == architecturalRegMap_23 ? 1'h0 : _GEN_4093; // @[decode.scala 393:{46,46}]
  wire  _GEN_4222 = 6'hc == architecturalRegMap_23 ? 1'h0 : _GEN_4094; // @[decode.scala 393:{46,46}]
  wire  _GEN_4223 = 6'hd == architecturalRegMap_23 ? 1'h0 : _GEN_4095; // @[decode.scala 393:{46,46}]
  wire  _GEN_4224 = 6'he == architecturalRegMap_23 ? 1'h0 : _GEN_4096; // @[decode.scala 393:{46,46}]
  wire  _GEN_4225 = 6'hf == architecturalRegMap_23 ? 1'h0 : _GEN_4097; // @[decode.scala 393:{46,46}]
  wire  _GEN_4226 = 6'h10 == architecturalRegMap_23 ? 1'h0 : _GEN_4098; // @[decode.scala 393:{46,46}]
  wire  _GEN_4227 = 6'h11 == architecturalRegMap_23 ? 1'h0 : _GEN_4099; // @[decode.scala 393:{46,46}]
  wire  _GEN_4228 = 6'h12 == architecturalRegMap_23 ? 1'h0 : _GEN_4100; // @[decode.scala 393:{46,46}]
  wire  _GEN_4229 = 6'h13 == architecturalRegMap_23 ? 1'h0 : _GEN_4101; // @[decode.scala 393:{46,46}]
  wire  _GEN_4230 = 6'h14 == architecturalRegMap_23 ? 1'h0 : _GEN_4102; // @[decode.scala 393:{46,46}]
  wire  _GEN_4231 = 6'h15 == architecturalRegMap_23 ? 1'h0 : _GEN_4103; // @[decode.scala 393:{46,46}]
  wire  _GEN_4232 = 6'h16 == architecturalRegMap_23 ? 1'h0 : _GEN_4104; // @[decode.scala 393:{46,46}]
  wire  _GEN_4233 = 6'h17 == architecturalRegMap_23 ? 1'h0 : _GEN_4105; // @[decode.scala 393:{46,46}]
  wire  _GEN_4234 = 6'h18 == architecturalRegMap_23 ? 1'h0 : _GEN_4106; // @[decode.scala 393:{46,46}]
  wire  _GEN_4235 = 6'h19 == architecturalRegMap_23 ? 1'h0 : _GEN_4107; // @[decode.scala 393:{46,46}]
  wire  _GEN_4236 = 6'h1a == architecturalRegMap_23 ? 1'h0 : _GEN_4108; // @[decode.scala 393:{46,46}]
  wire  _GEN_4237 = 6'h1b == architecturalRegMap_23 ? 1'h0 : _GEN_4109; // @[decode.scala 393:{46,46}]
  wire  _GEN_4238 = 6'h1c == architecturalRegMap_23 ? 1'h0 : _GEN_4110; // @[decode.scala 393:{46,46}]
  wire  _GEN_4239 = 6'h1d == architecturalRegMap_23 ? 1'h0 : _GEN_4111; // @[decode.scala 393:{46,46}]
  wire  _GEN_4240 = 6'h1e == architecturalRegMap_23 ? 1'h0 : _GEN_4112; // @[decode.scala 393:{46,46}]
  wire  _GEN_4241 = 6'h1f == architecturalRegMap_23 ? 1'h0 : _GEN_4113; // @[decode.scala 393:{46,46}]
  wire  _GEN_4242 = 6'h20 == architecturalRegMap_23 ? 1'h0 : _GEN_4114; // @[decode.scala 393:{46,46}]
  wire  _GEN_4243 = 6'h21 == architecturalRegMap_23 ? 1'h0 : _GEN_4115; // @[decode.scala 393:{46,46}]
  wire  _GEN_4244 = 6'h22 == architecturalRegMap_23 ? 1'h0 : _GEN_4116; // @[decode.scala 393:{46,46}]
  wire  _GEN_4245 = 6'h23 == architecturalRegMap_23 ? 1'h0 : _GEN_4117; // @[decode.scala 393:{46,46}]
  wire  _GEN_4246 = 6'h24 == architecturalRegMap_23 ? 1'h0 : _GEN_4118; // @[decode.scala 393:{46,46}]
  wire  _GEN_4247 = 6'h25 == architecturalRegMap_23 ? 1'h0 : _GEN_4119; // @[decode.scala 393:{46,46}]
  wire  _GEN_4248 = 6'h26 == architecturalRegMap_23 ? 1'h0 : _GEN_4120; // @[decode.scala 393:{46,46}]
  wire  _GEN_4249 = 6'h27 == architecturalRegMap_23 ? 1'h0 : _GEN_4121; // @[decode.scala 393:{46,46}]
  wire  _GEN_4250 = 6'h28 == architecturalRegMap_23 ? 1'h0 : _GEN_4122; // @[decode.scala 393:{46,46}]
  wire  _GEN_4251 = 6'h29 == architecturalRegMap_23 ? 1'h0 : _GEN_4123; // @[decode.scala 393:{46,46}]
  wire  _GEN_4252 = 6'h2a == architecturalRegMap_23 ? 1'h0 : _GEN_4124; // @[decode.scala 393:{46,46}]
  wire  _GEN_4253 = 6'h2b == architecturalRegMap_23 ? 1'h0 : _GEN_4125; // @[decode.scala 393:{46,46}]
  wire  _GEN_4254 = 6'h2c == architecturalRegMap_23 ? 1'h0 : _GEN_4126; // @[decode.scala 393:{46,46}]
  wire  _GEN_4255 = 6'h2d == architecturalRegMap_23 ? 1'h0 : _GEN_4127; // @[decode.scala 393:{46,46}]
  wire  _GEN_4256 = 6'h2e == architecturalRegMap_23 ? 1'h0 : _GEN_4128; // @[decode.scala 393:{46,46}]
  wire  _GEN_4257 = 6'h2f == architecturalRegMap_23 ? 1'h0 : _GEN_4129; // @[decode.scala 393:{46,46}]
  wire  _GEN_4258 = 6'h30 == architecturalRegMap_23 ? 1'h0 : _GEN_4130; // @[decode.scala 393:{46,46}]
  wire  _GEN_4259 = 6'h31 == architecturalRegMap_23 ? 1'h0 : _GEN_4131; // @[decode.scala 393:{46,46}]
  wire  _GEN_4260 = 6'h32 == architecturalRegMap_23 ? 1'h0 : _GEN_4132; // @[decode.scala 393:{46,46}]
  wire  _GEN_4261 = 6'h33 == architecturalRegMap_23 ? 1'h0 : _GEN_4133; // @[decode.scala 393:{46,46}]
  wire  _GEN_4262 = 6'h34 == architecturalRegMap_23 ? 1'h0 : _GEN_4134; // @[decode.scala 393:{46,46}]
  wire  _GEN_4263 = 6'h35 == architecturalRegMap_23 ? 1'h0 : _GEN_4135; // @[decode.scala 393:{46,46}]
  wire  _GEN_4264 = 6'h36 == architecturalRegMap_23 ? 1'h0 : _GEN_4136; // @[decode.scala 393:{46,46}]
  wire  _GEN_4265 = 6'h37 == architecturalRegMap_23 ? 1'h0 : _GEN_4137; // @[decode.scala 393:{46,46}]
  wire  _GEN_4266 = 6'h38 == architecturalRegMap_23 ? 1'h0 : _GEN_4138; // @[decode.scala 393:{46,46}]
  wire  _GEN_4267 = 6'h39 == architecturalRegMap_23 ? 1'h0 : _GEN_4139; // @[decode.scala 393:{46,46}]
  wire  _GEN_4268 = 6'h3a == architecturalRegMap_23 ? 1'h0 : _GEN_4140; // @[decode.scala 393:{46,46}]
  wire  _GEN_4269 = 6'h3b == architecturalRegMap_23 ? 1'h0 : _GEN_4141; // @[decode.scala 393:{46,46}]
  wire  _GEN_4270 = 6'h3c == architecturalRegMap_23 ? 1'h0 : _GEN_4142; // @[decode.scala 393:{46,46}]
  wire  _GEN_4271 = 6'h3d == architecturalRegMap_23 ? 1'h0 : _GEN_4143; // @[decode.scala 393:{46,46}]
  wire  _GEN_4272 = 6'h3e == architecturalRegMap_23 ? 1'h0 : _GEN_4144; // @[decode.scala 393:{46,46}]
  wire  _GEN_4338 = 6'h0 == architecturalRegMap_24 ? 1'h0 : _GEN_4210; // @[decode.scala 393:{46,46}]
  wire  _GEN_4339 = 6'h1 == architecturalRegMap_24 ? 1'h0 : _GEN_4211; // @[decode.scala 393:{46,46}]
  wire  _GEN_4340 = 6'h2 == architecturalRegMap_24 ? 1'h0 : _GEN_4212; // @[decode.scala 393:{46,46}]
  wire  _GEN_4341 = 6'h3 == architecturalRegMap_24 ? 1'h0 : _GEN_4213; // @[decode.scala 393:{46,46}]
  wire  _GEN_4342 = 6'h4 == architecturalRegMap_24 ? 1'h0 : _GEN_4214; // @[decode.scala 393:{46,46}]
  wire  _GEN_4343 = 6'h5 == architecturalRegMap_24 ? 1'h0 : _GEN_4215; // @[decode.scala 393:{46,46}]
  wire  _GEN_4344 = 6'h6 == architecturalRegMap_24 ? 1'h0 : _GEN_4216; // @[decode.scala 393:{46,46}]
  wire  _GEN_4345 = 6'h7 == architecturalRegMap_24 ? 1'h0 : _GEN_4217; // @[decode.scala 393:{46,46}]
  wire  _GEN_4346 = 6'h8 == architecturalRegMap_24 ? 1'h0 : _GEN_4218; // @[decode.scala 393:{46,46}]
  wire  _GEN_4347 = 6'h9 == architecturalRegMap_24 ? 1'h0 : _GEN_4219; // @[decode.scala 393:{46,46}]
  wire  _GEN_4348 = 6'ha == architecturalRegMap_24 ? 1'h0 : _GEN_4220; // @[decode.scala 393:{46,46}]
  wire  _GEN_4349 = 6'hb == architecturalRegMap_24 ? 1'h0 : _GEN_4221; // @[decode.scala 393:{46,46}]
  wire  _GEN_4350 = 6'hc == architecturalRegMap_24 ? 1'h0 : _GEN_4222; // @[decode.scala 393:{46,46}]
  wire  _GEN_4351 = 6'hd == architecturalRegMap_24 ? 1'h0 : _GEN_4223; // @[decode.scala 393:{46,46}]
  wire  _GEN_4352 = 6'he == architecturalRegMap_24 ? 1'h0 : _GEN_4224; // @[decode.scala 393:{46,46}]
  wire  _GEN_4353 = 6'hf == architecturalRegMap_24 ? 1'h0 : _GEN_4225; // @[decode.scala 393:{46,46}]
  wire  _GEN_4354 = 6'h10 == architecturalRegMap_24 ? 1'h0 : _GEN_4226; // @[decode.scala 393:{46,46}]
  wire  _GEN_4355 = 6'h11 == architecturalRegMap_24 ? 1'h0 : _GEN_4227; // @[decode.scala 393:{46,46}]
  wire  _GEN_4356 = 6'h12 == architecturalRegMap_24 ? 1'h0 : _GEN_4228; // @[decode.scala 393:{46,46}]
  wire  _GEN_4357 = 6'h13 == architecturalRegMap_24 ? 1'h0 : _GEN_4229; // @[decode.scala 393:{46,46}]
  wire  _GEN_4358 = 6'h14 == architecturalRegMap_24 ? 1'h0 : _GEN_4230; // @[decode.scala 393:{46,46}]
  wire  _GEN_4359 = 6'h15 == architecturalRegMap_24 ? 1'h0 : _GEN_4231; // @[decode.scala 393:{46,46}]
  wire  _GEN_4360 = 6'h16 == architecturalRegMap_24 ? 1'h0 : _GEN_4232; // @[decode.scala 393:{46,46}]
  wire  _GEN_4361 = 6'h17 == architecturalRegMap_24 ? 1'h0 : _GEN_4233; // @[decode.scala 393:{46,46}]
  wire  _GEN_4362 = 6'h18 == architecturalRegMap_24 ? 1'h0 : _GEN_4234; // @[decode.scala 393:{46,46}]
  wire  _GEN_4363 = 6'h19 == architecturalRegMap_24 ? 1'h0 : _GEN_4235; // @[decode.scala 393:{46,46}]
  wire  _GEN_4364 = 6'h1a == architecturalRegMap_24 ? 1'h0 : _GEN_4236; // @[decode.scala 393:{46,46}]
  wire  _GEN_4365 = 6'h1b == architecturalRegMap_24 ? 1'h0 : _GEN_4237; // @[decode.scala 393:{46,46}]
  wire  _GEN_4366 = 6'h1c == architecturalRegMap_24 ? 1'h0 : _GEN_4238; // @[decode.scala 393:{46,46}]
  wire  _GEN_4367 = 6'h1d == architecturalRegMap_24 ? 1'h0 : _GEN_4239; // @[decode.scala 393:{46,46}]
  wire  _GEN_4368 = 6'h1e == architecturalRegMap_24 ? 1'h0 : _GEN_4240; // @[decode.scala 393:{46,46}]
  wire  _GEN_4369 = 6'h1f == architecturalRegMap_24 ? 1'h0 : _GEN_4241; // @[decode.scala 393:{46,46}]
  wire  _GEN_4370 = 6'h20 == architecturalRegMap_24 ? 1'h0 : _GEN_4242; // @[decode.scala 393:{46,46}]
  wire  _GEN_4371 = 6'h21 == architecturalRegMap_24 ? 1'h0 : _GEN_4243; // @[decode.scala 393:{46,46}]
  wire  _GEN_4372 = 6'h22 == architecturalRegMap_24 ? 1'h0 : _GEN_4244; // @[decode.scala 393:{46,46}]
  wire  _GEN_4373 = 6'h23 == architecturalRegMap_24 ? 1'h0 : _GEN_4245; // @[decode.scala 393:{46,46}]
  wire  _GEN_4374 = 6'h24 == architecturalRegMap_24 ? 1'h0 : _GEN_4246; // @[decode.scala 393:{46,46}]
  wire  _GEN_4375 = 6'h25 == architecturalRegMap_24 ? 1'h0 : _GEN_4247; // @[decode.scala 393:{46,46}]
  wire  _GEN_4376 = 6'h26 == architecturalRegMap_24 ? 1'h0 : _GEN_4248; // @[decode.scala 393:{46,46}]
  wire  _GEN_4377 = 6'h27 == architecturalRegMap_24 ? 1'h0 : _GEN_4249; // @[decode.scala 393:{46,46}]
  wire  _GEN_4378 = 6'h28 == architecturalRegMap_24 ? 1'h0 : _GEN_4250; // @[decode.scala 393:{46,46}]
  wire  _GEN_4379 = 6'h29 == architecturalRegMap_24 ? 1'h0 : _GEN_4251; // @[decode.scala 393:{46,46}]
  wire  _GEN_4380 = 6'h2a == architecturalRegMap_24 ? 1'h0 : _GEN_4252; // @[decode.scala 393:{46,46}]
  wire  _GEN_4381 = 6'h2b == architecturalRegMap_24 ? 1'h0 : _GEN_4253; // @[decode.scala 393:{46,46}]
  wire  _GEN_4382 = 6'h2c == architecturalRegMap_24 ? 1'h0 : _GEN_4254; // @[decode.scala 393:{46,46}]
  wire  _GEN_4383 = 6'h2d == architecturalRegMap_24 ? 1'h0 : _GEN_4255; // @[decode.scala 393:{46,46}]
  wire  _GEN_4384 = 6'h2e == architecturalRegMap_24 ? 1'h0 : _GEN_4256; // @[decode.scala 393:{46,46}]
  wire  _GEN_4385 = 6'h2f == architecturalRegMap_24 ? 1'h0 : _GEN_4257; // @[decode.scala 393:{46,46}]
  wire  _GEN_4386 = 6'h30 == architecturalRegMap_24 ? 1'h0 : _GEN_4258; // @[decode.scala 393:{46,46}]
  wire  _GEN_4387 = 6'h31 == architecturalRegMap_24 ? 1'h0 : _GEN_4259; // @[decode.scala 393:{46,46}]
  wire  _GEN_4388 = 6'h32 == architecturalRegMap_24 ? 1'h0 : _GEN_4260; // @[decode.scala 393:{46,46}]
  wire  _GEN_4389 = 6'h33 == architecturalRegMap_24 ? 1'h0 : _GEN_4261; // @[decode.scala 393:{46,46}]
  wire  _GEN_4390 = 6'h34 == architecturalRegMap_24 ? 1'h0 : _GEN_4262; // @[decode.scala 393:{46,46}]
  wire  _GEN_4391 = 6'h35 == architecturalRegMap_24 ? 1'h0 : _GEN_4263; // @[decode.scala 393:{46,46}]
  wire  _GEN_4392 = 6'h36 == architecturalRegMap_24 ? 1'h0 : _GEN_4264; // @[decode.scala 393:{46,46}]
  wire  _GEN_4393 = 6'h37 == architecturalRegMap_24 ? 1'h0 : _GEN_4265; // @[decode.scala 393:{46,46}]
  wire  _GEN_4394 = 6'h38 == architecturalRegMap_24 ? 1'h0 : _GEN_4266; // @[decode.scala 393:{46,46}]
  wire  _GEN_4395 = 6'h39 == architecturalRegMap_24 ? 1'h0 : _GEN_4267; // @[decode.scala 393:{46,46}]
  wire  _GEN_4396 = 6'h3a == architecturalRegMap_24 ? 1'h0 : _GEN_4268; // @[decode.scala 393:{46,46}]
  wire  _GEN_4397 = 6'h3b == architecturalRegMap_24 ? 1'h0 : _GEN_4269; // @[decode.scala 393:{46,46}]
  wire  _GEN_4398 = 6'h3c == architecturalRegMap_24 ? 1'h0 : _GEN_4270; // @[decode.scala 393:{46,46}]
  wire  _GEN_4399 = 6'h3d == architecturalRegMap_24 ? 1'h0 : _GEN_4271; // @[decode.scala 393:{46,46}]
  wire  _GEN_4400 = 6'h3e == architecturalRegMap_24 ? 1'h0 : _GEN_4272; // @[decode.scala 393:{46,46}]
  wire  _GEN_4466 = 6'h0 == architecturalRegMap_25 ? 1'h0 : _GEN_4338; // @[decode.scala 393:{46,46}]
  wire  _GEN_4467 = 6'h1 == architecturalRegMap_25 ? 1'h0 : _GEN_4339; // @[decode.scala 393:{46,46}]
  wire  _GEN_4468 = 6'h2 == architecturalRegMap_25 ? 1'h0 : _GEN_4340; // @[decode.scala 393:{46,46}]
  wire  _GEN_4469 = 6'h3 == architecturalRegMap_25 ? 1'h0 : _GEN_4341; // @[decode.scala 393:{46,46}]
  wire  _GEN_4470 = 6'h4 == architecturalRegMap_25 ? 1'h0 : _GEN_4342; // @[decode.scala 393:{46,46}]
  wire  _GEN_4471 = 6'h5 == architecturalRegMap_25 ? 1'h0 : _GEN_4343; // @[decode.scala 393:{46,46}]
  wire  _GEN_4472 = 6'h6 == architecturalRegMap_25 ? 1'h0 : _GEN_4344; // @[decode.scala 393:{46,46}]
  wire  _GEN_4473 = 6'h7 == architecturalRegMap_25 ? 1'h0 : _GEN_4345; // @[decode.scala 393:{46,46}]
  wire  _GEN_4474 = 6'h8 == architecturalRegMap_25 ? 1'h0 : _GEN_4346; // @[decode.scala 393:{46,46}]
  wire  _GEN_4475 = 6'h9 == architecturalRegMap_25 ? 1'h0 : _GEN_4347; // @[decode.scala 393:{46,46}]
  wire  _GEN_4476 = 6'ha == architecturalRegMap_25 ? 1'h0 : _GEN_4348; // @[decode.scala 393:{46,46}]
  wire  _GEN_4477 = 6'hb == architecturalRegMap_25 ? 1'h0 : _GEN_4349; // @[decode.scala 393:{46,46}]
  wire  _GEN_4478 = 6'hc == architecturalRegMap_25 ? 1'h0 : _GEN_4350; // @[decode.scala 393:{46,46}]
  wire  _GEN_4479 = 6'hd == architecturalRegMap_25 ? 1'h0 : _GEN_4351; // @[decode.scala 393:{46,46}]
  wire  _GEN_4480 = 6'he == architecturalRegMap_25 ? 1'h0 : _GEN_4352; // @[decode.scala 393:{46,46}]
  wire  _GEN_4481 = 6'hf == architecturalRegMap_25 ? 1'h0 : _GEN_4353; // @[decode.scala 393:{46,46}]
  wire  _GEN_4482 = 6'h10 == architecturalRegMap_25 ? 1'h0 : _GEN_4354; // @[decode.scala 393:{46,46}]
  wire  _GEN_4483 = 6'h11 == architecturalRegMap_25 ? 1'h0 : _GEN_4355; // @[decode.scala 393:{46,46}]
  wire  _GEN_4484 = 6'h12 == architecturalRegMap_25 ? 1'h0 : _GEN_4356; // @[decode.scala 393:{46,46}]
  wire  _GEN_4485 = 6'h13 == architecturalRegMap_25 ? 1'h0 : _GEN_4357; // @[decode.scala 393:{46,46}]
  wire  _GEN_4486 = 6'h14 == architecturalRegMap_25 ? 1'h0 : _GEN_4358; // @[decode.scala 393:{46,46}]
  wire  _GEN_4487 = 6'h15 == architecturalRegMap_25 ? 1'h0 : _GEN_4359; // @[decode.scala 393:{46,46}]
  wire  _GEN_4488 = 6'h16 == architecturalRegMap_25 ? 1'h0 : _GEN_4360; // @[decode.scala 393:{46,46}]
  wire  _GEN_4489 = 6'h17 == architecturalRegMap_25 ? 1'h0 : _GEN_4361; // @[decode.scala 393:{46,46}]
  wire  _GEN_4490 = 6'h18 == architecturalRegMap_25 ? 1'h0 : _GEN_4362; // @[decode.scala 393:{46,46}]
  wire  _GEN_4491 = 6'h19 == architecturalRegMap_25 ? 1'h0 : _GEN_4363; // @[decode.scala 393:{46,46}]
  wire  _GEN_4492 = 6'h1a == architecturalRegMap_25 ? 1'h0 : _GEN_4364; // @[decode.scala 393:{46,46}]
  wire  _GEN_4493 = 6'h1b == architecturalRegMap_25 ? 1'h0 : _GEN_4365; // @[decode.scala 393:{46,46}]
  wire  _GEN_4494 = 6'h1c == architecturalRegMap_25 ? 1'h0 : _GEN_4366; // @[decode.scala 393:{46,46}]
  wire  _GEN_4495 = 6'h1d == architecturalRegMap_25 ? 1'h0 : _GEN_4367; // @[decode.scala 393:{46,46}]
  wire  _GEN_4496 = 6'h1e == architecturalRegMap_25 ? 1'h0 : _GEN_4368; // @[decode.scala 393:{46,46}]
  wire  _GEN_4497 = 6'h1f == architecturalRegMap_25 ? 1'h0 : _GEN_4369; // @[decode.scala 393:{46,46}]
  wire  _GEN_4498 = 6'h20 == architecturalRegMap_25 ? 1'h0 : _GEN_4370; // @[decode.scala 393:{46,46}]
  wire  _GEN_4499 = 6'h21 == architecturalRegMap_25 ? 1'h0 : _GEN_4371; // @[decode.scala 393:{46,46}]
  wire  _GEN_4500 = 6'h22 == architecturalRegMap_25 ? 1'h0 : _GEN_4372; // @[decode.scala 393:{46,46}]
  wire  _GEN_4501 = 6'h23 == architecturalRegMap_25 ? 1'h0 : _GEN_4373; // @[decode.scala 393:{46,46}]
  wire  _GEN_4502 = 6'h24 == architecturalRegMap_25 ? 1'h0 : _GEN_4374; // @[decode.scala 393:{46,46}]
  wire  _GEN_4503 = 6'h25 == architecturalRegMap_25 ? 1'h0 : _GEN_4375; // @[decode.scala 393:{46,46}]
  wire  _GEN_4504 = 6'h26 == architecturalRegMap_25 ? 1'h0 : _GEN_4376; // @[decode.scala 393:{46,46}]
  wire  _GEN_4505 = 6'h27 == architecturalRegMap_25 ? 1'h0 : _GEN_4377; // @[decode.scala 393:{46,46}]
  wire  _GEN_4506 = 6'h28 == architecturalRegMap_25 ? 1'h0 : _GEN_4378; // @[decode.scala 393:{46,46}]
  wire  _GEN_4507 = 6'h29 == architecturalRegMap_25 ? 1'h0 : _GEN_4379; // @[decode.scala 393:{46,46}]
  wire  _GEN_4508 = 6'h2a == architecturalRegMap_25 ? 1'h0 : _GEN_4380; // @[decode.scala 393:{46,46}]
  wire  _GEN_4509 = 6'h2b == architecturalRegMap_25 ? 1'h0 : _GEN_4381; // @[decode.scala 393:{46,46}]
  wire  _GEN_4510 = 6'h2c == architecturalRegMap_25 ? 1'h0 : _GEN_4382; // @[decode.scala 393:{46,46}]
  wire  _GEN_4511 = 6'h2d == architecturalRegMap_25 ? 1'h0 : _GEN_4383; // @[decode.scala 393:{46,46}]
  wire  _GEN_4512 = 6'h2e == architecturalRegMap_25 ? 1'h0 : _GEN_4384; // @[decode.scala 393:{46,46}]
  wire  _GEN_4513 = 6'h2f == architecturalRegMap_25 ? 1'h0 : _GEN_4385; // @[decode.scala 393:{46,46}]
  wire  _GEN_4514 = 6'h30 == architecturalRegMap_25 ? 1'h0 : _GEN_4386; // @[decode.scala 393:{46,46}]
  wire  _GEN_4515 = 6'h31 == architecturalRegMap_25 ? 1'h0 : _GEN_4387; // @[decode.scala 393:{46,46}]
  wire  _GEN_4516 = 6'h32 == architecturalRegMap_25 ? 1'h0 : _GEN_4388; // @[decode.scala 393:{46,46}]
  wire  _GEN_4517 = 6'h33 == architecturalRegMap_25 ? 1'h0 : _GEN_4389; // @[decode.scala 393:{46,46}]
  wire  _GEN_4518 = 6'h34 == architecturalRegMap_25 ? 1'h0 : _GEN_4390; // @[decode.scala 393:{46,46}]
  wire  _GEN_4519 = 6'h35 == architecturalRegMap_25 ? 1'h0 : _GEN_4391; // @[decode.scala 393:{46,46}]
  wire  _GEN_4520 = 6'h36 == architecturalRegMap_25 ? 1'h0 : _GEN_4392; // @[decode.scala 393:{46,46}]
  wire  _GEN_4521 = 6'h37 == architecturalRegMap_25 ? 1'h0 : _GEN_4393; // @[decode.scala 393:{46,46}]
  wire  _GEN_4522 = 6'h38 == architecturalRegMap_25 ? 1'h0 : _GEN_4394; // @[decode.scala 393:{46,46}]
  wire  _GEN_4523 = 6'h39 == architecturalRegMap_25 ? 1'h0 : _GEN_4395; // @[decode.scala 393:{46,46}]
  wire  _GEN_4524 = 6'h3a == architecturalRegMap_25 ? 1'h0 : _GEN_4396; // @[decode.scala 393:{46,46}]
  wire  _GEN_4525 = 6'h3b == architecturalRegMap_25 ? 1'h0 : _GEN_4397; // @[decode.scala 393:{46,46}]
  wire  _GEN_4526 = 6'h3c == architecturalRegMap_25 ? 1'h0 : _GEN_4398; // @[decode.scala 393:{46,46}]
  wire  _GEN_4527 = 6'h3d == architecturalRegMap_25 ? 1'h0 : _GEN_4399; // @[decode.scala 393:{46,46}]
  wire  _GEN_4528 = 6'h3e == architecturalRegMap_25 ? 1'h0 : _GEN_4400; // @[decode.scala 393:{46,46}]
  wire  _GEN_4594 = 6'h0 == architecturalRegMap_26 ? 1'h0 : _GEN_4466; // @[decode.scala 393:{46,46}]
  wire  _GEN_4595 = 6'h1 == architecturalRegMap_26 ? 1'h0 : _GEN_4467; // @[decode.scala 393:{46,46}]
  wire  _GEN_4596 = 6'h2 == architecturalRegMap_26 ? 1'h0 : _GEN_4468; // @[decode.scala 393:{46,46}]
  wire  _GEN_4597 = 6'h3 == architecturalRegMap_26 ? 1'h0 : _GEN_4469; // @[decode.scala 393:{46,46}]
  wire  _GEN_4598 = 6'h4 == architecturalRegMap_26 ? 1'h0 : _GEN_4470; // @[decode.scala 393:{46,46}]
  wire  _GEN_4599 = 6'h5 == architecturalRegMap_26 ? 1'h0 : _GEN_4471; // @[decode.scala 393:{46,46}]
  wire  _GEN_4600 = 6'h6 == architecturalRegMap_26 ? 1'h0 : _GEN_4472; // @[decode.scala 393:{46,46}]
  wire  _GEN_4601 = 6'h7 == architecturalRegMap_26 ? 1'h0 : _GEN_4473; // @[decode.scala 393:{46,46}]
  wire  _GEN_4602 = 6'h8 == architecturalRegMap_26 ? 1'h0 : _GEN_4474; // @[decode.scala 393:{46,46}]
  wire  _GEN_4603 = 6'h9 == architecturalRegMap_26 ? 1'h0 : _GEN_4475; // @[decode.scala 393:{46,46}]
  wire  _GEN_4604 = 6'ha == architecturalRegMap_26 ? 1'h0 : _GEN_4476; // @[decode.scala 393:{46,46}]
  wire  _GEN_4605 = 6'hb == architecturalRegMap_26 ? 1'h0 : _GEN_4477; // @[decode.scala 393:{46,46}]
  wire  _GEN_4606 = 6'hc == architecturalRegMap_26 ? 1'h0 : _GEN_4478; // @[decode.scala 393:{46,46}]
  wire  _GEN_4607 = 6'hd == architecturalRegMap_26 ? 1'h0 : _GEN_4479; // @[decode.scala 393:{46,46}]
  wire  _GEN_4608 = 6'he == architecturalRegMap_26 ? 1'h0 : _GEN_4480; // @[decode.scala 393:{46,46}]
  wire  _GEN_4609 = 6'hf == architecturalRegMap_26 ? 1'h0 : _GEN_4481; // @[decode.scala 393:{46,46}]
  wire  _GEN_4610 = 6'h10 == architecturalRegMap_26 ? 1'h0 : _GEN_4482; // @[decode.scala 393:{46,46}]
  wire  _GEN_4611 = 6'h11 == architecturalRegMap_26 ? 1'h0 : _GEN_4483; // @[decode.scala 393:{46,46}]
  wire  _GEN_4612 = 6'h12 == architecturalRegMap_26 ? 1'h0 : _GEN_4484; // @[decode.scala 393:{46,46}]
  wire  _GEN_4613 = 6'h13 == architecturalRegMap_26 ? 1'h0 : _GEN_4485; // @[decode.scala 393:{46,46}]
  wire  _GEN_4614 = 6'h14 == architecturalRegMap_26 ? 1'h0 : _GEN_4486; // @[decode.scala 393:{46,46}]
  wire  _GEN_4615 = 6'h15 == architecturalRegMap_26 ? 1'h0 : _GEN_4487; // @[decode.scala 393:{46,46}]
  wire  _GEN_4616 = 6'h16 == architecturalRegMap_26 ? 1'h0 : _GEN_4488; // @[decode.scala 393:{46,46}]
  wire  _GEN_4617 = 6'h17 == architecturalRegMap_26 ? 1'h0 : _GEN_4489; // @[decode.scala 393:{46,46}]
  wire  _GEN_4618 = 6'h18 == architecturalRegMap_26 ? 1'h0 : _GEN_4490; // @[decode.scala 393:{46,46}]
  wire  _GEN_4619 = 6'h19 == architecturalRegMap_26 ? 1'h0 : _GEN_4491; // @[decode.scala 393:{46,46}]
  wire  _GEN_4620 = 6'h1a == architecturalRegMap_26 ? 1'h0 : _GEN_4492; // @[decode.scala 393:{46,46}]
  wire  _GEN_4621 = 6'h1b == architecturalRegMap_26 ? 1'h0 : _GEN_4493; // @[decode.scala 393:{46,46}]
  wire  _GEN_4622 = 6'h1c == architecturalRegMap_26 ? 1'h0 : _GEN_4494; // @[decode.scala 393:{46,46}]
  wire  _GEN_4623 = 6'h1d == architecturalRegMap_26 ? 1'h0 : _GEN_4495; // @[decode.scala 393:{46,46}]
  wire  _GEN_4624 = 6'h1e == architecturalRegMap_26 ? 1'h0 : _GEN_4496; // @[decode.scala 393:{46,46}]
  wire  _GEN_4625 = 6'h1f == architecturalRegMap_26 ? 1'h0 : _GEN_4497; // @[decode.scala 393:{46,46}]
  wire  _GEN_4626 = 6'h20 == architecturalRegMap_26 ? 1'h0 : _GEN_4498; // @[decode.scala 393:{46,46}]
  wire  _GEN_4627 = 6'h21 == architecturalRegMap_26 ? 1'h0 : _GEN_4499; // @[decode.scala 393:{46,46}]
  wire  _GEN_4628 = 6'h22 == architecturalRegMap_26 ? 1'h0 : _GEN_4500; // @[decode.scala 393:{46,46}]
  wire  _GEN_4629 = 6'h23 == architecturalRegMap_26 ? 1'h0 : _GEN_4501; // @[decode.scala 393:{46,46}]
  wire  _GEN_4630 = 6'h24 == architecturalRegMap_26 ? 1'h0 : _GEN_4502; // @[decode.scala 393:{46,46}]
  wire  _GEN_4631 = 6'h25 == architecturalRegMap_26 ? 1'h0 : _GEN_4503; // @[decode.scala 393:{46,46}]
  wire  _GEN_4632 = 6'h26 == architecturalRegMap_26 ? 1'h0 : _GEN_4504; // @[decode.scala 393:{46,46}]
  wire  _GEN_4633 = 6'h27 == architecturalRegMap_26 ? 1'h0 : _GEN_4505; // @[decode.scala 393:{46,46}]
  wire  _GEN_4634 = 6'h28 == architecturalRegMap_26 ? 1'h0 : _GEN_4506; // @[decode.scala 393:{46,46}]
  wire  _GEN_4635 = 6'h29 == architecturalRegMap_26 ? 1'h0 : _GEN_4507; // @[decode.scala 393:{46,46}]
  wire  _GEN_4636 = 6'h2a == architecturalRegMap_26 ? 1'h0 : _GEN_4508; // @[decode.scala 393:{46,46}]
  wire  _GEN_4637 = 6'h2b == architecturalRegMap_26 ? 1'h0 : _GEN_4509; // @[decode.scala 393:{46,46}]
  wire  _GEN_4638 = 6'h2c == architecturalRegMap_26 ? 1'h0 : _GEN_4510; // @[decode.scala 393:{46,46}]
  wire  _GEN_4639 = 6'h2d == architecturalRegMap_26 ? 1'h0 : _GEN_4511; // @[decode.scala 393:{46,46}]
  wire  _GEN_4640 = 6'h2e == architecturalRegMap_26 ? 1'h0 : _GEN_4512; // @[decode.scala 393:{46,46}]
  wire  _GEN_4641 = 6'h2f == architecturalRegMap_26 ? 1'h0 : _GEN_4513; // @[decode.scala 393:{46,46}]
  wire  _GEN_4642 = 6'h30 == architecturalRegMap_26 ? 1'h0 : _GEN_4514; // @[decode.scala 393:{46,46}]
  wire  _GEN_4643 = 6'h31 == architecturalRegMap_26 ? 1'h0 : _GEN_4515; // @[decode.scala 393:{46,46}]
  wire  _GEN_4644 = 6'h32 == architecturalRegMap_26 ? 1'h0 : _GEN_4516; // @[decode.scala 393:{46,46}]
  wire  _GEN_4645 = 6'h33 == architecturalRegMap_26 ? 1'h0 : _GEN_4517; // @[decode.scala 393:{46,46}]
  wire  _GEN_4646 = 6'h34 == architecturalRegMap_26 ? 1'h0 : _GEN_4518; // @[decode.scala 393:{46,46}]
  wire  _GEN_4647 = 6'h35 == architecturalRegMap_26 ? 1'h0 : _GEN_4519; // @[decode.scala 393:{46,46}]
  wire  _GEN_4648 = 6'h36 == architecturalRegMap_26 ? 1'h0 : _GEN_4520; // @[decode.scala 393:{46,46}]
  wire  _GEN_4649 = 6'h37 == architecturalRegMap_26 ? 1'h0 : _GEN_4521; // @[decode.scala 393:{46,46}]
  wire  _GEN_4650 = 6'h38 == architecturalRegMap_26 ? 1'h0 : _GEN_4522; // @[decode.scala 393:{46,46}]
  wire  _GEN_4651 = 6'h39 == architecturalRegMap_26 ? 1'h0 : _GEN_4523; // @[decode.scala 393:{46,46}]
  wire  _GEN_4652 = 6'h3a == architecturalRegMap_26 ? 1'h0 : _GEN_4524; // @[decode.scala 393:{46,46}]
  wire  _GEN_4653 = 6'h3b == architecturalRegMap_26 ? 1'h0 : _GEN_4525; // @[decode.scala 393:{46,46}]
  wire  _GEN_4654 = 6'h3c == architecturalRegMap_26 ? 1'h0 : _GEN_4526; // @[decode.scala 393:{46,46}]
  wire  _GEN_4655 = 6'h3d == architecturalRegMap_26 ? 1'h0 : _GEN_4527; // @[decode.scala 393:{46,46}]
  wire  _GEN_4656 = 6'h3e == architecturalRegMap_26 ? 1'h0 : _GEN_4528; // @[decode.scala 393:{46,46}]
  wire  _GEN_4722 = 6'h0 == architecturalRegMap_27 ? 1'h0 : _GEN_4594; // @[decode.scala 393:{46,46}]
  wire  _GEN_4723 = 6'h1 == architecturalRegMap_27 ? 1'h0 : _GEN_4595; // @[decode.scala 393:{46,46}]
  wire  _GEN_4724 = 6'h2 == architecturalRegMap_27 ? 1'h0 : _GEN_4596; // @[decode.scala 393:{46,46}]
  wire  _GEN_4725 = 6'h3 == architecturalRegMap_27 ? 1'h0 : _GEN_4597; // @[decode.scala 393:{46,46}]
  wire  _GEN_4726 = 6'h4 == architecturalRegMap_27 ? 1'h0 : _GEN_4598; // @[decode.scala 393:{46,46}]
  wire  _GEN_4727 = 6'h5 == architecturalRegMap_27 ? 1'h0 : _GEN_4599; // @[decode.scala 393:{46,46}]
  wire  _GEN_4728 = 6'h6 == architecturalRegMap_27 ? 1'h0 : _GEN_4600; // @[decode.scala 393:{46,46}]
  wire  _GEN_4729 = 6'h7 == architecturalRegMap_27 ? 1'h0 : _GEN_4601; // @[decode.scala 393:{46,46}]
  wire  _GEN_4730 = 6'h8 == architecturalRegMap_27 ? 1'h0 : _GEN_4602; // @[decode.scala 393:{46,46}]
  wire  _GEN_4731 = 6'h9 == architecturalRegMap_27 ? 1'h0 : _GEN_4603; // @[decode.scala 393:{46,46}]
  wire  _GEN_4732 = 6'ha == architecturalRegMap_27 ? 1'h0 : _GEN_4604; // @[decode.scala 393:{46,46}]
  wire  _GEN_4733 = 6'hb == architecturalRegMap_27 ? 1'h0 : _GEN_4605; // @[decode.scala 393:{46,46}]
  wire  _GEN_4734 = 6'hc == architecturalRegMap_27 ? 1'h0 : _GEN_4606; // @[decode.scala 393:{46,46}]
  wire  _GEN_4735 = 6'hd == architecturalRegMap_27 ? 1'h0 : _GEN_4607; // @[decode.scala 393:{46,46}]
  wire  _GEN_4736 = 6'he == architecturalRegMap_27 ? 1'h0 : _GEN_4608; // @[decode.scala 393:{46,46}]
  wire  _GEN_4737 = 6'hf == architecturalRegMap_27 ? 1'h0 : _GEN_4609; // @[decode.scala 393:{46,46}]
  wire  _GEN_4738 = 6'h10 == architecturalRegMap_27 ? 1'h0 : _GEN_4610; // @[decode.scala 393:{46,46}]
  wire  _GEN_4739 = 6'h11 == architecturalRegMap_27 ? 1'h0 : _GEN_4611; // @[decode.scala 393:{46,46}]
  wire  _GEN_4740 = 6'h12 == architecturalRegMap_27 ? 1'h0 : _GEN_4612; // @[decode.scala 393:{46,46}]
  wire  _GEN_4741 = 6'h13 == architecturalRegMap_27 ? 1'h0 : _GEN_4613; // @[decode.scala 393:{46,46}]
  wire  _GEN_4742 = 6'h14 == architecturalRegMap_27 ? 1'h0 : _GEN_4614; // @[decode.scala 393:{46,46}]
  wire  _GEN_4743 = 6'h15 == architecturalRegMap_27 ? 1'h0 : _GEN_4615; // @[decode.scala 393:{46,46}]
  wire  _GEN_4744 = 6'h16 == architecturalRegMap_27 ? 1'h0 : _GEN_4616; // @[decode.scala 393:{46,46}]
  wire  _GEN_4745 = 6'h17 == architecturalRegMap_27 ? 1'h0 : _GEN_4617; // @[decode.scala 393:{46,46}]
  wire  _GEN_4746 = 6'h18 == architecturalRegMap_27 ? 1'h0 : _GEN_4618; // @[decode.scala 393:{46,46}]
  wire  _GEN_4747 = 6'h19 == architecturalRegMap_27 ? 1'h0 : _GEN_4619; // @[decode.scala 393:{46,46}]
  wire  _GEN_4748 = 6'h1a == architecturalRegMap_27 ? 1'h0 : _GEN_4620; // @[decode.scala 393:{46,46}]
  wire  _GEN_4749 = 6'h1b == architecturalRegMap_27 ? 1'h0 : _GEN_4621; // @[decode.scala 393:{46,46}]
  wire  _GEN_4750 = 6'h1c == architecturalRegMap_27 ? 1'h0 : _GEN_4622; // @[decode.scala 393:{46,46}]
  wire  _GEN_4751 = 6'h1d == architecturalRegMap_27 ? 1'h0 : _GEN_4623; // @[decode.scala 393:{46,46}]
  wire  _GEN_4752 = 6'h1e == architecturalRegMap_27 ? 1'h0 : _GEN_4624; // @[decode.scala 393:{46,46}]
  wire  _GEN_4753 = 6'h1f == architecturalRegMap_27 ? 1'h0 : _GEN_4625; // @[decode.scala 393:{46,46}]
  wire  _GEN_4754 = 6'h20 == architecturalRegMap_27 ? 1'h0 : _GEN_4626; // @[decode.scala 393:{46,46}]
  wire  _GEN_4755 = 6'h21 == architecturalRegMap_27 ? 1'h0 : _GEN_4627; // @[decode.scala 393:{46,46}]
  wire  _GEN_4756 = 6'h22 == architecturalRegMap_27 ? 1'h0 : _GEN_4628; // @[decode.scala 393:{46,46}]
  wire  _GEN_4757 = 6'h23 == architecturalRegMap_27 ? 1'h0 : _GEN_4629; // @[decode.scala 393:{46,46}]
  wire  _GEN_4758 = 6'h24 == architecturalRegMap_27 ? 1'h0 : _GEN_4630; // @[decode.scala 393:{46,46}]
  wire  _GEN_4759 = 6'h25 == architecturalRegMap_27 ? 1'h0 : _GEN_4631; // @[decode.scala 393:{46,46}]
  wire  _GEN_4760 = 6'h26 == architecturalRegMap_27 ? 1'h0 : _GEN_4632; // @[decode.scala 393:{46,46}]
  wire  _GEN_4761 = 6'h27 == architecturalRegMap_27 ? 1'h0 : _GEN_4633; // @[decode.scala 393:{46,46}]
  wire  _GEN_4762 = 6'h28 == architecturalRegMap_27 ? 1'h0 : _GEN_4634; // @[decode.scala 393:{46,46}]
  wire  _GEN_4763 = 6'h29 == architecturalRegMap_27 ? 1'h0 : _GEN_4635; // @[decode.scala 393:{46,46}]
  wire  _GEN_4764 = 6'h2a == architecturalRegMap_27 ? 1'h0 : _GEN_4636; // @[decode.scala 393:{46,46}]
  wire  _GEN_4765 = 6'h2b == architecturalRegMap_27 ? 1'h0 : _GEN_4637; // @[decode.scala 393:{46,46}]
  wire  _GEN_4766 = 6'h2c == architecturalRegMap_27 ? 1'h0 : _GEN_4638; // @[decode.scala 393:{46,46}]
  wire  _GEN_4767 = 6'h2d == architecturalRegMap_27 ? 1'h0 : _GEN_4639; // @[decode.scala 393:{46,46}]
  wire  _GEN_4768 = 6'h2e == architecturalRegMap_27 ? 1'h0 : _GEN_4640; // @[decode.scala 393:{46,46}]
  wire  _GEN_4769 = 6'h2f == architecturalRegMap_27 ? 1'h0 : _GEN_4641; // @[decode.scala 393:{46,46}]
  wire  _GEN_4770 = 6'h30 == architecturalRegMap_27 ? 1'h0 : _GEN_4642; // @[decode.scala 393:{46,46}]
  wire  _GEN_4771 = 6'h31 == architecturalRegMap_27 ? 1'h0 : _GEN_4643; // @[decode.scala 393:{46,46}]
  wire  _GEN_4772 = 6'h32 == architecturalRegMap_27 ? 1'h0 : _GEN_4644; // @[decode.scala 393:{46,46}]
  wire  _GEN_4773 = 6'h33 == architecturalRegMap_27 ? 1'h0 : _GEN_4645; // @[decode.scala 393:{46,46}]
  wire  _GEN_4774 = 6'h34 == architecturalRegMap_27 ? 1'h0 : _GEN_4646; // @[decode.scala 393:{46,46}]
  wire  _GEN_4775 = 6'h35 == architecturalRegMap_27 ? 1'h0 : _GEN_4647; // @[decode.scala 393:{46,46}]
  wire  _GEN_4776 = 6'h36 == architecturalRegMap_27 ? 1'h0 : _GEN_4648; // @[decode.scala 393:{46,46}]
  wire  _GEN_4777 = 6'h37 == architecturalRegMap_27 ? 1'h0 : _GEN_4649; // @[decode.scala 393:{46,46}]
  wire  _GEN_4778 = 6'h38 == architecturalRegMap_27 ? 1'h0 : _GEN_4650; // @[decode.scala 393:{46,46}]
  wire  _GEN_4779 = 6'h39 == architecturalRegMap_27 ? 1'h0 : _GEN_4651; // @[decode.scala 393:{46,46}]
  wire  _GEN_4780 = 6'h3a == architecturalRegMap_27 ? 1'h0 : _GEN_4652; // @[decode.scala 393:{46,46}]
  wire  _GEN_4781 = 6'h3b == architecturalRegMap_27 ? 1'h0 : _GEN_4653; // @[decode.scala 393:{46,46}]
  wire  _GEN_4782 = 6'h3c == architecturalRegMap_27 ? 1'h0 : _GEN_4654; // @[decode.scala 393:{46,46}]
  wire  _GEN_4783 = 6'h3d == architecturalRegMap_27 ? 1'h0 : _GEN_4655; // @[decode.scala 393:{46,46}]
  wire  _GEN_4784 = 6'h3e == architecturalRegMap_27 ? 1'h0 : _GEN_4656; // @[decode.scala 393:{46,46}]
  wire  _GEN_4850 = 6'h0 == architecturalRegMap_28 ? 1'h0 : _GEN_4722; // @[decode.scala 393:{46,46}]
  wire  _GEN_4851 = 6'h1 == architecturalRegMap_28 ? 1'h0 : _GEN_4723; // @[decode.scala 393:{46,46}]
  wire  _GEN_4852 = 6'h2 == architecturalRegMap_28 ? 1'h0 : _GEN_4724; // @[decode.scala 393:{46,46}]
  wire  _GEN_4853 = 6'h3 == architecturalRegMap_28 ? 1'h0 : _GEN_4725; // @[decode.scala 393:{46,46}]
  wire  _GEN_4854 = 6'h4 == architecturalRegMap_28 ? 1'h0 : _GEN_4726; // @[decode.scala 393:{46,46}]
  wire  _GEN_4855 = 6'h5 == architecturalRegMap_28 ? 1'h0 : _GEN_4727; // @[decode.scala 393:{46,46}]
  wire  _GEN_4856 = 6'h6 == architecturalRegMap_28 ? 1'h0 : _GEN_4728; // @[decode.scala 393:{46,46}]
  wire  _GEN_4857 = 6'h7 == architecturalRegMap_28 ? 1'h0 : _GEN_4729; // @[decode.scala 393:{46,46}]
  wire  _GEN_4858 = 6'h8 == architecturalRegMap_28 ? 1'h0 : _GEN_4730; // @[decode.scala 393:{46,46}]
  wire  _GEN_4859 = 6'h9 == architecturalRegMap_28 ? 1'h0 : _GEN_4731; // @[decode.scala 393:{46,46}]
  wire  _GEN_4860 = 6'ha == architecturalRegMap_28 ? 1'h0 : _GEN_4732; // @[decode.scala 393:{46,46}]
  wire  _GEN_4861 = 6'hb == architecturalRegMap_28 ? 1'h0 : _GEN_4733; // @[decode.scala 393:{46,46}]
  wire  _GEN_4862 = 6'hc == architecturalRegMap_28 ? 1'h0 : _GEN_4734; // @[decode.scala 393:{46,46}]
  wire  _GEN_4863 = 6'hd == architecturalRegMap_28 ? 1'h0 : _GEN_4735; // @[decode.scala 393:{46,46}]
  wire  _GEN_4864 = 6'he == architecturalRegMap_28 ? 1'h0 : _GEN_4736; // @[decode.scala 393:{46,46}]
  wire  _GEN_4865 = 6'hf == architecturalRegMap_28 ? 1'h0 : _GEN_4737; // @[decode.scala 393:{46,46}]
  wire  _GEN_4866 = 6'h10 == architecturalRegMap_28 ? 1'h0 : _GEN_4738; // @[decode.scala 393:{46,46}]
  wire  _GEN_4867 = 6'h11 == architecturalRegMap_28 ? 1'h0 : _GEN_4739; // @[decode.scala 393:{46,46}]
  wire  _GEN_4868 = 6'h12 == architecturalRegMap_28 ? 1'h0 : _GEN_4740; // @[decode.scala 393:{46,46}]
  wire  _GEN_4869 = 6'h13 == architecturalRegMap_28 ? 1'h0 : _GEN_4741; // @[decode.scala 393:{46,46}]
  wire  _GEN_4870 = 6'h14 == architecturalRegMap_28 ? 1'h0 : _GEN_4742; // @[decode.scala 393:{46,46}]
  wire  _GEN_4871 = 6'h15 == architecturalRegMap_28 ? 1'h0 : _GEN_4743; // @[decode.scala 393:{46,46}]
  wire  _GEN_4872 = 6'h16 == architecturalRegMap_28 ? 1'h0 : _GEN_4744; // @[decode.scala 393:{46,46}]
  wire  _GEN_4873 = 6'h17 == architecturalRegMap_28 ? 1'h0 : _GEN_4745; // @[decode.scala 393:{46,46}]
  wire  _GEN_4874 = 6'h18 == architecturalRegMap_28 ? 1'h0 : _GEN_4746; // @[decode.scala 393:{46,46}]
  wire  _GEN_4875 = 6'h19 == architecturalRegMap_28 ? 1'h0 : _GEN_4747; // @[decode.scala 393:{46,46}]
  wire  _GEN_4876 = 6'h1a == architecturalRegMap_28 ? 1'h0 : _GEN_4748; // @[decode.scala 393:{46,46}]
  wire  _GEN_4877 = 6'h1b == architecturalRegMap_28 ? 1'h0 : _GEN_4749; // @[decode.scala 393:{46,46}]
  wire  _GEN_4878 = 6'h1c == architecturalRegMap_28 ? 1'h0 : _GEN_4750; // @[decode.scala 393:{46,46}]
  wire  _GEN_4879 = 6'h1d == architecturalRegMap_28 ? 1'h0 : _GEN_4751; // @[decode.scala 393:{46,46}]
  wire  _GEN_4880 = 6'h1e == architecturalRegMap_28 ? 1'h0 : _GEN_4752; // @[decode.scala 393:{46,46}]
  wire  _GEN_4881 = 6'h1f == architecturalRegMap_28 ? 1'h0 : _GEN_4753; // @[decode.scala 393:{46,46}]
  wire  _GEN_4882 = 6'h20 == architecturalRegMap_28 ? 1'h0 : _GEN_4754; // @[decode.scala 393:{46,46}]
  wire  _GEN_4883 = 6'h21 == architecturalRegMap_28 ? 1'h0 : _GEN_4755; // @[decode.scala 393:{46,46}]
  wire  _GEN_4884 = 6'h22 == architecturalRegMap_28 ? 1'h0 : _GEN_4756; // @[decode.scala 393:{46,46}]
  wire  _GEN_4885 = 6'h23 == architecturalRegMap_28 ? 1'h0 : _GEN_4757; // @[decode.scala 393:{46,46}]
  wire  _GEN_4886 = 6'h24 == architecturalRegMap_28 ? 1'h0 : _GEN_4758; // @[decode.scala 393:{46,46}]
  wire  _GEN_4887 = 6'h25 == architecturalRegMap_28 ? 1'h0 : _GEN_4759; // @[decode.scala 393:{46,46}]
  wire  _GEN_4888 = 6'h26 == architecturalRegMap_28 ? 1'h0 : _GEN_4760; // @[decode.scala 393:{46,46}]
  wire  _GEN_4889 = 6'h27 == architecturalRegMap_28 ? 1'h0 : _GEN_4761; // @[decode.scala 393:{46,46}]
  wire  _GEN_4890 = 6'h28 == architecturalRegMap_28 ? 1'h0 : _GEN_4762; // @[decode.scala 393:{46,46}]
  wire  _GEN_4891 = 6'h29 == architecturalRegMap_28 ? 1'h0 : _GEN_4763; // @[decode.scala 393:{46,46}]
  wire  _GEN_4892 = 6'h2a == architecturalRegMap_28 ? 1'h0 : _GEN_4764; // @[decode.scala 393:{46,46}]
  wire  _GEN_4893 = 6'h2b == architecturalRegMap_28 ? 1'h0 : _GEN_4765; // @[decode.scala 393:{46,46}]
  wire  _GEN_4894 = 6'h2c == architecturalRegMap_28 ? 1'h0 : _GEN_4766; // @[decode.scala 393:{46,46}]
  wire  _GEN_4895 = 6'h2d == architecturalRegMap_28 ? 1'h0 : _GEN_4767; // @[decode.scala 393:{46,46}]
  wire  _GEN_4896 = 6'h2e == architecturalRegMap_28 ? 1'h0 : _GEN_4768; // @[decode.scala 393:{46,46}]
  wire  _GEN_4897 = 6'h2f == architecturalRegMap_28 ? 1'h0 : _GEN_4769; // @[decode.scala 393:{46,46}]
  wire  _GEN_4898 = 6'h30 == architecturalRegMap_28 ? 1'h0 : _GEN_4770; // @[decode.scala 393:{46,46}]
  wire  _GEN_4899 = 6'h31 == architecturalRegMap_28 ? 1'h0 : _GEN_4771; // @[decode.scala 393:{46,46}]
  wire  _GEN_4900 = 6'h32 == architecturalRegMap_28 ? 1'h0 : _GEN_4772; // @[decode.scala 393:{46,46}]
  wire  _GEN_4901 = 6'h33 == architecturalRegMap_28 ? 1'h0 : _GEN_4773; // @[decode.scala 393:{46,46}]
  wire  _GEN_4902 = 6'h34 == architecturalRegMap_28 ? 1'h0 : _GEN_4774; // @[decode.scala 393:{46,46}]
  wire  _GEN_4903 = 6'h35 == architecturalRegMap_28 ? 1'h0 : _GEN_4775; // @[decode.scala 393:{46,46}]
  wire  _GEN_4904 = 6'h36 == architecturalRegMap_28 ? 1'h0 : _GEN_4776; // @[decode.scala 393:{46,46}]
  wire  _GEN_4905 = 6'h37 == architecturalRegMap_28 ? 1'h0 : _GEN_4777; // @[decode.scala 393:{46,46}]
  wire  _GEN_4906 = 6'h38 == architecturalRegMap_28 ? 1'h0 : _GEN_4778; // @[decode.scala 393:{46,46}]
  wire  _GEN_4907 = 6'h39 == architecturalRegMap_28 ? 1'h0 : _GEN_4779; // @[decode.scala 393:{46,46}]
  wire  _GEN_4908 = 6'h3a == architecturalRegMap_28 ? 1'h0 : _GEN_4780; // @[decode.scala 393:{46,46}]
  wire  _GEN_4909 = 6'h3b == architecturalRegMap_28 ? 1'h0 : _GEN_4781; // @[decode.scala 393:{46,46}]
  wire  _GEN_4910 = 6'h3c == architecturalRegMap_28 ? 1'h0 : _GEN_4782; // @[decode.scala 393:{46,46}]
  wire  _GEN_4911 = 6'h3d == architecturalRegMap_28 ? 1'h0 : _GEN_4783; // @[decode.scala 393:{46,46}]
  wire  _GEN_4912 = 6'h3e == architecturalRegMap_28 ? 1'h0 : _GEN_4784; // @[decode.scala 393:{46,46}]
  wire  _GEN_4978 = 6'h0 == architecturalRegMap_29 ? 1'h0 : _GEN_4850; // @[decode.scala 393:{46,46}]
  wire  _GEN_4979 = 6'h1 == architecturalRegMap_29 ? 1'h0 : _GEN_4851; // @[decode.scala 393:{46,46}]
  wire  _GEN_4980 = 6'h2 == architecturalRegMap_29 ? 1'h0 : _GEN_4852; // @[decode.scala 393:{46,46}]
  wire  _GEN_4981 = 6'h3 == architecturalRegMap_29 ? 1'h0 : _GEN_4853; // @[decode.scala 393:{46,46}]
  wire  _GEN_4982 = 6'h4 == architecturalRegMap_29 ? 1'h0 : _GEN_4854; // @[decode.scala 393:{46,46}]
  wire  _GEN_4983 = 6'h5 == architecturalRegMap_29 ? 1'h0 : _GEN_4855; // @[decode.scala 393:{46,46}]
  wire  _GEN_4984 = 6'h6 == architecturalRegMap_29 ? 1'h0 : _GEN_4856; // @[decode.scala 393:{46,46}]
  wire  _GEN_4985 = 6'h7 == architecturalRegMap_29 ? 1'h0 : _GEN_4857; // @[decode.scala 393:{46,46}]
  wire  _GEN_4986 = 6'h8 == architecturalRegMap_29 ? 1'h0 : _GEN_4858; // @[decode.scala 393:{46,46}]
  wire  _GEN_4987 = 6'h9 == architecturalRegMap_29 ? 1'h0 : _GEN_4859; // @[decode.scala 393:{46,46}]
  wire  _GEN_4988 = 6'ha == architecturalRegMap_29 ? 1'h0 : _GEN_4860; // @[decode.scala 393:{46,46}]
  wire  _GEN_4989 = 6'hb == architecturalRegMap_29 ? 1'h0 : _GEN_4861; // @[decode.scala 393:{46,46}]
  wire  _GEN_4990 = 6'hc == architecturalRegMap_29 ? 1'h0 : _GEN_4862; // @[decode.scala 393:{46,46}]
  wire  _GEN_4991 = 6'hd == architecturalRegMap_29 ? 1'h0 : _GEN_4863; // @[decode.scala 393:{46,46}]
  wire  _GEN_4992 = 6'he == architecturalRegMap_29 ? 1'h0 : _GEN_4864; // @[decode.scala 393:{46,46}]
  wire  _GEN_4993 = 6'hf == architecturalRegMap_29 ? 1'h0 : _GEN_4865; // @[decode.scala 393:{46,46}]
  wire  _GEN_4994 = 6'h10 == architecturalRegMap_29 ? 1'h0 : _GEN_4866; // @[decode.scala 393:{46,46}]
  wire  _GEN_4995 = 6'h11 == architecturalRegMap_29 ? 1'h0 : _GEN_4867; // @[decode.scala 393:{46,46}]
  wire  _GEN_4996 = 6'h12 == architecturalRegMap_29 ? 1'h0 : _GEN_4868; // @[decode.scala 393:{46,46}]
  wire  _GEN_4997 = 6'h13 == architecturalRegMap_29 ? 1'h0 : _GEN_4869; // @[decode.scala 393:{46,46}]
  wire  _GEN_4998 = 6'h14 == architecturalRegMap_29 ? 1'h0 : _GEN_4870; // @[decode.scala 393:{46,46}]
  wire  _GEN_4999 = 6'h15 == architecturalRegMap_29 ? 1'h0 : _GEN_4871; // @[decode.scala 393:{46,46}]
  wire  _GEN_5000 = 6'h16 == architecturalRegMap_29 ? 1'h0 : _GEN_4872; // @[decode.scala 393:{46,46}]
  wire  _GEN_5001 = 6'h17 == architecturalRegMap_29 ? 1'h0 : _GEN_4873; // @[decode.scala 393:{46,46}]
  wire  _GEN_5002 = 6'h18 == architecturalRegMap_29 ? 1'h0 : _GEN_4874; // @[decode.scala 393:{46,46}]
  wire  _GEN_5003 = 6'h19 == architecturalRegMap_29 ? 1'h0 : _GEN_4875; // @[decode.scala 393:{46,46}]
  wire  _GEN_5004 = 6'h1a == architecturalRegMap_29 ? 1'h0 : _GEN_4876; // @[decode.scala 393:{46,46}]
  wire  _GEN_5005 = 6'h1b == architecturalRegMap_29 ? 1'h0 : _GEN_4877; // @[decode.scala 393:{46,46}]
  wire  _GEN_5006 = 6'h1c == architecturalRegMap_29 ? 1'h0 : _GEN_4878; // @[decode.scala 393:{46,46}]
  wire  _GEN_5007 = 6'h1d == architecturalRegMap_29 ? 1'h0 : _GEN_4879; // @[decode.scala 393:{46,46}]
  wire  _GEN_5008 = 6'h1e == architecturalRegMap_29 ? 1'h0 : _GEN_4880; // @[decode.scala 393:{46,46}]
  wire  _GEN_5009 = 6'h1f == architecturalRegMap_29 ? 1'h0 : _GEN_4881; // @[decode.scala 393:{46,46}]
  wire  _GEN_5010 = 6'h20 == architecturalRegMap_29 ? 1'h0 : _GEN_4882; // @[decode.scala 393:{46,46}]
  wire  _GEN_5011 = 6'h21 == architecturalRegMap_29 ? 1'h0 : _GEN_4883; // @[decode.scala 393:{46,46}]
  wire  _GEN_5012 = 6'h22 == architecturalRegMap_29 ? 1'h0 : _GEN_4884; // @[decode.scala 393:{46,46}]
  wire  _GEN_5013 = 6'h23 == architecturalRegMap_29 ? 1'h0 : _GEN_4885; // @[decode.scala 393:{46,46}]
  wire  _GEN_5014 = 6'h24 == architecturalRegMap_29 ? 1'h0 : _GEN_4886; // @[decode.scala 393:{46,46}]
  wire  _GEN_5015 = 6'h25 == architecturalRegMap_29 ? 1'h0 : _GEN_4887; // @[decode.scala 393:{46,46}]
  wire  _GEN_5016 = 6'h26 == architecturalRegMap_29 ? 1'h0 : _GEN_4888; // @[decode.scala 393:{46,46}]
  wire  _GEN_5017 = 6'h27 == architecturalRegMap_29 ? 1'h0 : _GEN_4889; // @[decode.scala 393:{46,46}]
  wire  _GEN_5018 = 6'h28 == architecturalRegMap_29 ? 1'h0 : _GEN_4890; // @[decode.scala 393:{46,46}]
  wire  _GEN_5019 = 6'h29 == architecturalRegMap_29 ? 1'h0 : _GEN_4891; // @[decode.scala 393:{46,46}]
  wire  _GEN_5020 = 6'h2a == architecturalRegMap_29 ? 1'h0 : _GEN_4892; // @[decode.scala 393:{46,46}]
  wire  _GEN_5021 = 6'h2b == architecturalRegMap_29 ? 1'h0 : _GEN_4893; // @[decode.scala 393:{46,46}]
  wire  _GEN_5022 = 6'h2c == architecturalRegMap_29 ? 1'h0 : _GEN_4894; // @[decode.scala 393:{46,46}]
  wire  _GEN_5023 = 6'h2d == architecturalRegMap_29 ? 1'h0 : _GEN_4895; // @[decode.scala 393:{46,46}]
  wire  _GEN_5024 = 6'h2e == architecturalRegMap_29 ? 1'h0 : _GEN_4896; // @[decode.scala 393:{46,46}]
  wire  _GEN_5025 = 6'h2f == architecturalRegMap_29 ? 1'h0 : _GEN_4897; // @[decode.scala 393:{46,46}]
  wire  _GEN_5026 = 6'h30 == architecturalRegMap_29 ? 1'h0 : _GEN_4898; // @[decode.scala 393:{46,46}]
  wire  _GEN_5027 = 6'h31 == architecturalRegMap_29 ? 1'h0 : _GEN_4899; // @[decode.scala 393:{46,46}]
  wire  _GEN_5028 = 6'h32 == architecturalRegMap_29 ? 1'h0 : _GEN_4900; // @[decode.scala 393:{46,46}]
  wire  _GEN_5029 = 6'h33 == architecturalRegMap_29 ? 1'h0 : _GEN_4901; // @[decode.scala 393:{46,46}]
  wire  _GEN_5030 = 6'h34 == architecturalRegMap_29 ? 1'h0 : _GEN_4902; // @[decode.scala 393:{46,46}]
  wire  _GEN_5031 = 6'h35 == architecturalRegMap_29 ? 1'h0 : _GEN_4903; // @[decode.scala 393:{46,46}]
  wire  _GEN_5032 = 6'h36 == architecturalRegMap_29 ? 1'h0 : _GEN_4904; // @[decode.scala 393:{46,46}]
  wire  _GEN_5033 = 6'h37 == architecturalRegMap_29 ? 1'h0 : _GEN_4905; // @[decode.scala 393:{46,46}]
  wire  _GEN_5034 = 6'h38 == architecturalRegMap_29 ? 1'h0 : _GEN_4906; // @[decode.scala 393:{46,46}]
  wire  _GEN_5035 = 6'h39 == architecturalRegMap_29 ? 1'h0 : _GEN_4907; // @[decode.scala 393:{46,46}]
  wire  _GEN_5036 = 6'h3a == architecturalRegMap_29 ? 1'h0 : _GEN_4908; // @[decode.scala 393:{46,46}]
  wire  _GEN_5037 = 6'h3b == architecturalRegMap_29 ? 1'h0 : _GEN_4909; // @[decode.scala 393:{46,46}]
  wire  _GEN_5038 = 6'h3c == architecturalRegMap_29 ? 1'h0 : _GEN_4910; // @[decode.scala 393:{46,46}]
  wire  _GEN_5039 = 6'h3d == architecturalRegMap_29 ? 1'h0 : _GEN_4911; // @[decode.scala 393:{46,46}]
  wire  _GEN_5040 = 6'h3e == architecturalRegMap_29 ? 1'h0 : _GEN_4912; // @[decode.scala 393:{46,46}]
  wire  _GEN_5042 = 6'h0 == architecturalRegMap_30 | (6'h0 == architecturalRegMap_29 | (6'h0 == architecturalRegMap_28
     | (6'h0 == architecturalRegMap_27 | (6'h0 == architecturalRegMap_26 | (6'h0 == architecturalRegMap_25 | (6'h0 ==
    architecturalRegMap_24 | (6'h0 == architecturalRegMap_23 | (6'h0 == architecturalRegMap_22 | (6'h0 ==
    architecturalRegMap_21 | (6'h0 == architecturalRegMap_20 | (6'h0 == architecturalRegMap_19 | (6'h0 ==
    architecturalRegMap_18 | (6'h0 == architecturalRegMap_17 | (6'h0 == architecturalRegMap_16 | _GEN_3122))))))))))))))
    ; // @[decode.scala 392:{47,47}]
  wire  _GEN_5043 = 6'h1 == architecturalRegMap_30 | (6'h1 == architecturalRegMap_29 | (6'h1 == architecturalRegMap_28
     | (6'h1 == architecturalRegMap_27 | (6'h1 == architecturalRegMap_26 | (6'h1 == architecturalRegMap_25 | (6'h1 ==
    architecturalRegMap_24 | (6'h1 == architecturalRegMap_23 | (6'h1 == architecturalRegMap_22 | (6'h1 ==
    architecturalRegMap_21 | (6'h1 == architecturalRegMap_20 | (6'h1 == architecturalRegMap_19 | (6'h1 ==
    architecturalRegMap_18 | (6'h1 == architecturalRegMap_17 | (6'h1 == architecturalRegMap_16 | _GEN_3123))))))))))))))
    ; // @[decode.scala 392:{47,47}]
  wire  _GEN_5044 = 6'h2 == architecturalRegMap_30 | (6'h2 == architecturalRegMap_29 | (6'h2 == architecturalRegMap_28
     | (6'h2 == architecturalRegMap_27 | (6'h2 == architecturalRegMap_26 | (6'h2 == architecturalRegMap_25 | (6'h2 ==
    architecturalRegMap_24 | (6'h2 == architecturalRegMap_23 | (6'h2 == architecturalRegMap_22 | (6'h2 ==
    architecturalRegMap_21 | (6'h2 == architecturalRegMap_20 | (6'h2 == architecturalRegMap_19 | (6'h2 ==
    architecturalRegMap_18 | (6'h2 == architecturalRegMap_17 | (6'h2 == architecturalRegMap_16 | _GEN_3124))))))))))))))
    ; // @[decode.scala 392:{47,47}]
  wire  _GEN_5045 = 6'h3 == architecturalRegMap_30 | (6'h3 == architecturalRegMap_29 | (6'h3 == architecturalRegMap_28
     | (6'h3 == architecturalRegMap_27 | (6'h3 == architecturalRegMap_26 | (6'h3 == architecturalRegMap_25 | (6'h3 ==
    architecturalRegMap_24 | (6'h3 == architecturalRegMap_23 | (6'h3 == architecturalRegMap_22 | (6'h3 ==
    architecturalRegMap_21 | (6'h3 == architecturalRegMap_20 | (6'h3 == architecturalRegMap_19 | (6'h3 ==
    architecturalRegMap_18 | (6'h3 == architecturalRegMap_17 | (6'h3 == architecturalRegMap_16 | _GEN_3125))))))))))))))
    ; // @[decode.scala 392:{47,47}]
  wire  _GEN_5046 = 6'h4 == architecturalRegMap_30 | (6'h4 == architecturalRegMap_29 | (6'h4 == architecturalRegMap_28
     | (6'h4 == architecturalRegMap_27 | (6'h4 == architecturalRegMap_26 | (6'h4 == architecturalRegMap_25 | (6'h4 ==
    architecturalRegMap_24 | (6'h4 == architecturalRegMap_23 | (6'h4 == architecturalRegMap_22 | (6'h4 ==
    architecturalRegMap_21 | (6'h4 == architecturalRegMap_20 | (6'h4 == architecturalRegMap_19 | (6'h4 ==
    architecturalRegMap_18 | (6'h4 == architecturalRegMap_17 | (6'h4 == architecturalRegMap_16 | _GEN_3126))))))))))))))
    ; // @[decode.scala 392:{47,47}]
  wire  _GEN_5047 = 6'h5 == architecturalRegMap_30 | (6'h5 == architecturalRegMap_29 | (6'h5 == architecturalRegMap_28
     | (6'h5 == architecturalRegMap_27 | (6'h5 == architecturalRegMap_26 | (6'h5 == architecturalRegMap_25 | (6'h5 ==
    architecturalRegMap_24 | (6'h5 == architecturalRegMap_23 | (6'h5 == architecturalRegMap_22 | (6'h5 ==
    architecturalRegMap_21 | (6'h5 == architecturalRegMap_20 | (6'h5 == architecturalRegMap_19 | (6'h5 ==
    architecturalRegMap_18 | (6'h5 == architecturalRegMap_17 | (6'h5 == architecturalRegMap_16 | _GEN_3127))))))))))))))
    ; // @[decode.scala 392:{47,47}]
  wire  _GEN_5048 = 6'h6 == architecturalRegMap_30 | (6'h6 == architecturalRegMap_29 | (6'h6 == architecturalRegMap_28
     | (6'h6 == architecturalRegMap_27 | (6'h6 == architecturalRegMap_26 | (6'h6 == architecturalRegMap_25 | (6'h6 ==
    architecturalRegMap_24 | (6'h6 == architecturalRegMap_23 | (6'h6 == architecturalRegMap_22 | (6'h6 ==
    architecturalRegMap_21 | (6'h6 == architecturalRegMap_20 | (6'h6 == architecturalRegMap_19 | (6'h6 ==
    architecturalRegMap_18 | (6'h6 == architecturalRegMap_17 | (6'h6 == architecturalRegMap_16 | _GEN_3128))))))))))))))
    ; // @[decode.scala 392:{47,47}]
  wire  _GEN_5049 = 6'h7 == architecturalRegMap_30 | (6'h7 == architecturalRegMap_29 | (6'h7 == architecturalRegMap_28
     | (6'h7 == architecturalRegMap_27 | (6'h7 == architecturalRegMap_26 | (6'h7 == architecturalRegMap_25 | (6'h7 ==
    architecturalRegMap_24 | (6'h7 == architecturalRegMap_23 | (6'h7 == architecturalRegMap_22 | (6'h7 ==
    architecturalRegMap_21 | (6'h7 == architecturalRegMap_20 | (6'h7 == architecturalRegMap_19 | (6'h7 ==
    architecturalRegMap_18 | (6'h7 == architecturalRegMap_17 | (6'h7 == architecturalRegMap_16 | _GEN_3129))))))))))))))
    ; // @[decode.scala 392:{47,47}]
  wire  _GEN_5050 = 6'h8 == architecturalRegMap_30 | (6'h8 == architecturalRegMap_29 | (6'h8 == architecturalRegMap_28
     | (6'h8 == architecturalRegMap_27 | (6'h8 == architecturalRegMap_26 | (6'h8 == architecturalRegMap_25 | (6'h8 ==
    architecturalRegMap_24 | (6'h8 == architecturalRegMap_23 | (6'h8 == architecturalRegMap_22 | (6'h8 ==
    architecturalRegMap_21 | (6'h8 == architecturalRegMap_20 | (6'h8 == architecturalRegMap_19 | (6'h8 ==
    architecturalRegMap_18 | (6'h8 == architecturalRegMap_17 | (6'h8 == architecturalRegMap_16 | _GEN_3130))))))))))))))
    ; // @[decode.scala 392:{47,47}]
  wire  _GEN_5051 = 6'h9 == architecturalRegMap_30 | (6'h9 == architecturalRegMap_29 | (6'h9 == architecturalRegMap_28
     | (6'h9 == architecturalRegMap_27 | (6'h9 == architecturalRegMap_26 | (6'h9 == architecturalRegMap_25 | (6'h9 ==
    architecturalRegMap_24 | (6'h9 == architecturalRegMap_23 | (6'h9 == architecturalRegMap_22 | (6'h9 ==
    architecturalRegMap_21 | (6'h9 == architecturalRegMap_20 | (6'h9 == architecturalRegMap_19 | (6'h9 ==
    architecturalRegMap_18 | (6'h9 == architecturalRegMap_17 | (6'h9 == architecturalRegMap_16 | _GEN_3131))))))))))))))
    ; // @[decode.scala 392:{47,47}]
  wire  _GEN_5052 = 6'ha == architecturalRegMap_30 | (6'ha == architecturalRegMap_29 | (6'ha == architecturalRegMap_28
     | (6'ha == architecturalRegMap_27 | (6'ha == architecturalRegMap_26 | (6'ha == architecturalRegMap_25 | (6'ha ==
    architecturalRegMap_24 | (6'ha == architecturalRegMap_23 | (6'ha == architecturalRegMap_22 | (6'ha ==
    architecturalRegMap_21 | (6'ha == architecturalRegMap_20 | (6'ha == architecturalRegMap_19 | (6'ha ==
    architecturalRegMap_18 | (6'ha == architecturalRegMap_17 | (6'ha == architecturalRegMap_16 | _GEN_3132))))))))))))))
    ; // @[decode.scala 392:{47,47}]
  wire  _GEN_5053 = 6'hb == architecturalRegMap_30 | (6'hb == architecturalRegMap_29 | (6'hb == architecturalRegMap_28
     | (6'hb == architecturalRegMap_27 | (6'hb == architecturalRegMap_26 | (6'hb == architecturalRegMap_25 | (6'hb ==
    architecturalRegMap_24 | (6'hb == architecturalRegMap_23 | (6'hb == architecturalRegMap_22 | (6'hb ==
    architecturalRegMap_21 | (6'hb == architecturalRegMap_20 | (6'hb == architecturalRegMap_19 | (6'hb ==
    architecturalRegMap_18 | (6'hb == architecturalRegMap_17 | (6'hb == architecturalRegMap_16 | _GEN_3133))))))))))))))
    ; // @[decode.scala 392:{47,47}]
  wire  _GEN_5054 = 6'hc == architecturalRegMap_30 | (6'hc == architecturalRegMap_29 | (6'hc == architecturalRegMap_28
     | (6'hc == architecturalRegMap_27 | (6'hc == architecturalRegMap_26 | (6'hc == architecturalRegMap_25 | (6'hc ==
    architecturalRegMap_24 | (6'hc == architecturalRegMap_23 | (6'hc == architecturalRegMap_22 | (6'hc ==
    architecturalRegMap_21 | (6'hc == architecturalRegMap_20 | (6'hc == architecturalRegMap_19 | (6'hc ==
    architecturalRegMap_18 | (6'hc == architecturalRegMap_17 | (6'hc == architecturalRegMap_16 | _GEN_3134))))))))))))))
    ; // @[decode.scala 392:{47,47}]
  wire  _GEN_5055 = 6'hd == architecturalRegMap_30 | (6'hd == architecturalRegMap_29 | (6'hd == architecturalRegMap_28
     | (6'hd == architecturalRegMap_27 | (6'hd == architecturalRegMap_26 | (6'hd == architecturalRegMap_25 | (6'hd ==
    architecturalRegMap_24 | (6'hd == architecturalRegMap_23 | (6'hd == architecturalRegMap_22 | (6'hd ==
    architecturalRegMap_21 | (6'hd == architecturalRegMap_20 | (6'hd == architecturalRegMap_19 | (6'hd ==
    architecturalRegMap_18 | (6'hd == architecturalRegMap_17 | (6'hd == architecturalRegMap_16 | _GEN_3135))))))))))))))
    ; // @[decode.scala 392:{47,47}]
  wire  _GEN_5056 = 6'he == architecturalRegMap_30 | (6'he == architecturalRegMap_29 | (6'he == architecturalRegMap_28
     | (6'he == architecturalRegMap_27 | (6'he == architecturalRegMap_26 | (6'he == architecturalRegMap_25 | (6'he ==
    architecturalRegMap_24 | (6'he == architecturalRegMap_23 | (6'he == architecturalRegMap_22 | (6'he ==
    architecturalRegMap_21 | (6'he == architecturalRegMap_20 | (6'he == architecturalRegMap_19 | (6'he ==
    architecturalRegMap_18 | (6'he == architecturalRegMap_17 | (6'he == architecturalRegMap_16 | _GEN_3136))))))))))))))
    ; // @[decode.scala 392:{47,47}]
  wire  _GEN_5057 = 6'hf == architecturalRegMap_30 | (6'hf == architecturalRegMap_29 | (6'hf == architecturalRegMap_28
     | (6'hf == architecturalRegMap_27 | (6'hf == architecturalRegMap_26 | (6'hf == architecturalRegMap_25 | (6'hf ==
    architecturalRegMap_24 | (6'hf == architecturalRegMap_23 | (6'hf == architecturalRegMap_22 | (6'hf ==
    architecturalRegMap_21 | (6'hf == architecturalRegMap_20 | (6'hf == architecturalRegMap_19 | (6'hf ==
    architecturalRegMap_18 | (6'hf == architecturalRegMap_17 | (6'hf == architecturalRegMap_16 | _GEN_3137))))))))))))))
    ; // @[decode.scala 392:{47,47}]
  wire  _GEN_5058 = 6'h10 == architecturalRegMap_30 | (6'h10 == architecturalRegMap_29 | (6'h10 ==
    architecturalRegMap_28 | (6'h10 == architecturalRegMap_27 | (6'h10 == architecturalRegMap_26 | (6'h10 ==
    architecturalRegMap_25 | (6'h10 == architecturalRegMap_24 | (6'h10 == architecturalRegMap_23 | (6'h10 ==
    architecturalRegMap_22 | (6'h10 == architecturalRegMap_21 | (6'h10 == architecturalRegMap_20 | (6'h10 ==
    architecturalRegMap_19 | (6'h10 == architecturalRegMap_18 | (6'h10 == architecturalRegMap_17 | (6'h10 ==
    architecturalRegMap_16 | _GEN_3138)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5059 = 6'h11 == architecturalRegMap_30 | (6'h11 == architecturalRegMap_29 | (6'h11 ==
    architecturalRegMap_28 | (6'h11 == architecturalRegMap_27 | (6'h11 == architecturalRegMap_26 | (6'h11 ==
    architecturalRegMap_25 | (6'h11 == architecturalRegMap_24 | (6'h11 == architecturalRegMap_23 | (6'h11 ==
    architecturalRegMap_22 | (6'h11 == architecturalRegMap_21 | (6'h11 == architecturalRegMap_20 | (6'h11 ==
    architecturalRegMap_19 | (6'h11 == architecturalRegMap_18 | (6'h11 == architecturalRegMap_17 | (6'h11 ==
    architecturalRegMap_16 | _GEN_3139)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5060 = 6'h12 == architecturalRegMap_30 | (6'h12 == architecturalRegMap_29 | (6'h12 ==
    architecturalRegMap_28 | (6'h12 == architecturalRegMap_27 | (6'h12 == architecturalRegMap_26 | (6'h12 ==
    architecturalRegMap_25 | (6'h12 == architecturalRegMap_24 | (6'h12 == architecturalRegMap_23 | (6'h12 ==
    architecturalRegMap_22 | (6'h12 == architecturalRegMap_21 | (6'h12 == architecturalRegMap_20 | (6'h12 ==
    architecturalRegMap_19 | (6'h12 == architecturalRegMap_18 | (6'h12 == architecturalRegMap_17 | (6'h12 ==
    architecturalRegMap_16 | _GEN_3140)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5061 = 6'h13 == architecturalRegMap_30 | (6'h13 == architecturalRegMap_29 | (6'h13 ==
    architecturalRegMap_28 | (6'h13 == architecturalRegMap_27 | (6'h13 == architecturalRegMap_26 | (6'h13 ==
    architecturalRegMap_25 | (6'h13 == architecturalRegMap_24 | (6'h13 == architecturalRegMap_23 | (6'h13 ==
    architecturalRegMap_22 | (6'h13 == architecturalRegMap_21 | (6'h13 == architecturalRegMap_20 | (6'h13 ==
    architecturalRegMap_19 | (6'h13 == architecturalRegMap_18 | (6'h13 == architecturalRegMap_17 | (6'h13 ==
    architecturalRegMap_16 | _GEN_3141)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5062 = 6'h14 == architecturalRegMap_30 | (6'h14 == architecturalRegMap_29 | (6'h14 ==
    architecturalRegMap_28 | (6'h14 == architecturalRegMap_27 | (6'h14 == architecturalRegMap_26 | (6'h14 ==
    architecturalRegMap_25 | (6'h14 == architecturalRegMap_24 | (6'h14 == architecturalRegMap_23 | (6'h14 ==
    architecturalRegMap_22 | (6'h14 == architecturalRegMap_21 | (6'h14 == architecturalRegMap_20 | (6'h14 ==
    architecturalRegMap_19 | (6'h14 == architecturalRegMap_18 | (6'h14 == architecturalRegMap_17 | (6'h14 ==
    architecturalRegMap_16 | _GEN_3142)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5063 = 6'h15 == architecturalRegMap_30 | (6'h15 == architecturalRegMap_29 | (6'h15 ==
    architecturalRegMap_28 | (6'h15 == architecturalRegMap_27 | (6'h15 == architecturalRegMap_26 | (6'h15 ==
    architecturalRegMap_25 | (6'h15 == architecturalRegMap_24 | (6'h15 == architecturalRegMap_23 | (6'h15 ==
    architecturalRegMap_22 | (6'h15 == architecturalRegMap_21 | (6'h15 == architecturalRegMap_20 | (6'h15 ==
    architecturalRegMap_19 | (6'h15 == architecturalRegMap_18 | (6'h15 == architecturalRegMap_17 | (6'h15 ==
    architecturalRegMap_16 | _GEN_3143)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5064 = 6'h16 == architecturalRegMap_30 | (6'h16 == architecturalRegMap_29 | (6'h16 ==
    architecturalRegMap_28 | (6'h16 == architecturalRegMap_27 | (6'h16 == architecturalRegMap_26 | (6'h16 ==
    architecturalRegMap_25 | (6'h16 == architecturalRegMap_24 | (6'h16 == architecturalRegMap_23 | (6'h16 ==
    architecturalRegMap_22 | (6'h16 == architecturalRegMap_21 | (6'h16 == architecturalRegMap_20 | (6'h16 ==
    architecturalRegMap_19 | (6'h16 == architecturalRegMap_18 | (6'h16 == architecturalRegMap_17 | (6'h16 ==
    architecturalRegMap_16 | _GEN_3144)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5065 = 6'h17 == architecturalRegMap_30 | (6'h17 == architecturalRegMap_29 | (6'h17 ==
    architecturalRegMap_28 | (6'h17 == architecturalRegMap_27 | (6'h17 == architecturalRegMap_26 | (6'h17 ==
    architecturalRegMap_25 | (6'h17 == architecturalRegMap_24 | (6'h17 == architecturalRegMap_23 | (6'h17 ==
    architecturalRegMap_22 | (6'h17 == architecturalRegMap_21 | (6'h17 == architecturalRegMap_20 | (6'h17 ==
    architecturalRegMap_19 | (6'h17 == architecturalRegMap_18 | (6'h17 == architecturalRegMap_17 | (6'h17 ==
    architecturalRegMap_16 | _GEN_3145)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5066 = 6'h18 == architecturalRegMap_30 | (6'h18 == architecturalRegMap_29 | (6'h18 ==
    architecturalRegMap_28 | (6'h18 == architecturalRegMap_27 | (6'h18 == architecturalRegMap_26 | (6'h18 ==
    architecturalRegMap_25 | (6'h18 == architecturalRegMap_24 | (6'h18 == architecturalRegMap_23 | (6'h18 ==
    architecturalRegMap_22 | (6'h18 == architecturalRegMap_21 | (6'h18 == architecturalRegMap_20 | (6'h18 ==
    architecturalRegMap_19 | (6'h18 == architecturalRegMap_18 | (6'h18 == architecturalRegMap_17 | (6'h18 ==
    architecturalRegMap_16 | _GEN_3146)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5067 = 6'h19 == architecturalRegMap_30 | (6'h19 == architecturalRegMap_29 | (6'h19 ==
    architecturalRegMap_28 | (6'h19 == architecturalRegMap_27 | (6'h19 == architecturalRegMap_26 | (6'h19 ==
    architecturalRegMap_25 | (6'h19 == architecturalRegMap_24 | (6'h19 == architecturalRegMap_23 | (6'h19 ==
    architecturalRegMap_22 | (6'h19 == architecturalRegMap_21 | (6'h19 == architecturalRegMap_20 | (6'h19 ==
    architecturalRegMap_19 | (6'h19 == architecturalRegMap_18 | (6'h19 == architecturalRegMap_17 | (6'h19 ==
    architecturalRegMap_16 | _GEN_3147)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5068 = 6'h1a == architecturalRegMap_30 | (6'h1a == architecturalRegMap_29 | (6'h1a ==
    architecturalRegMap_28 | (6'h1a == architecturalRegMap_27 | (6'h1a == architecturalRegMap_26 | (6'h1a ==
    architecturalRegMap_25 | (6'h1a == architecturalRegMap_24 | (6'h1a == architecturalRegMap_23 | (6'h1a ==
    architecturalRegMap_22 | (6'h1a == architecturalRegMap_21 | (6'h1a == architecturalRegMap_20 | (6'h1a ==
    architecturalRegMap_19 | (6'h1a == architecturalRegMap_18 | (6'h1a == architecturalRegMap_17 | (6'h1a ==
    architecturalRegMap_16 | _GEN_3148)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5069 = 6'h1b == architecturalRegMap_30 | (6'h1b == architecturalRegMap_29 | (6'h1b ==
    architecturalRegMap_28 | (6'h1b == architecturalRegMap_27 | (6'h1b == architecturalRegMap_26 | (6'h1b ==
    architecturalRegMap_25 | (6'h1b == architecturalRegMap_24 | (6'h1b == architecturalRegMap_23 | (6'h1b ==
    architecturalRegMap_22 | (6'h1b == architecturalRegMap_21 | (6'h1b == architecturalRegMap_20 | (6'h1b ==
    architecturalRegMap_19 | (6'h1b == architecturalRegMap_18 | (6'h1b == architecturalRegMap_17 | (6'h1b ==
    architecturalRegMap_16 | _GEN_3149)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5070 = 6'h1c == architecturalRegMap_30 | (6'h1c == architecturalRegMap_29 | (6'h1c ==
    architecturalRegMap_28 | (6'h1c == architecturalRegMap_27 | (6'h1c == architecturalRegMap_26 | (6'h1c ==
    architecturalRegMap_25 | (6'h1c == architecturalRegMap_24 | (6'h1c == architecturalRegMap_23 | (6'h1c ==
    architecturalRegMap_22 | (6'h1c == architecturalRegMap_21 | (6'h1c == architecturalRegMap_20 | (6'h1c ==
    architecturalRegMap_19 | (6'h1c == architecturalRegMap_18 | (6'h1c == architecturalRegMap_17 | (6'h1c ==
    architecturalRegMap_16 | _GEN_3150)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5071 = 6'h1d == architecturalRegMap_30 | (6'h1d == architecturalRegMap_29 | (6'h1d ==
    architecturalRegMap_28 | (6'h1d == architecturalRegMap_27 | (6'h1d == architecturalRegMap_26 | (6'h1d ==
    architecturalRegMap_25 | (6'h1d == architecturalRegMap_24 | (6'h1d == architecturalRegMap_23 | (6'h1d ==
    architecturalRegMap_22 | (6'h1d == architecturalRegMap_21 | (6'h1d == architecturalRegMap_20 | (6'h1d ==
    architecturalRegMap_19 | (6'h1d == architecturalRegMap_18 | (6'h1d == architecturalRegMap_17 | (6'h1d ==
    architecturalRegMap_16 | _GEN_3151)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5072 = 6'h1e == architecturalRegMap_30 | (6'h1e == architecturalRegMap_29 | (6'h1e ==
    architecturalRegMap_28 | (6'h1e == architecturalRegMap_27 | (6'h1e == architecturalRegMap_26 | (6'h1e ==
    architecturalRegMap_25 | (6'h1e == architecturalRegMap_24 | (6'h1e == architecturalRegMap_23 | (6'h1e ==
    architecturalRegMap_22 | (6'h1e == architecturalRegMap_21 | (6'h1e == architecturalRegMap_20 | (6'h1e ==
    architecturalRegMap_19 | (6'h1e == architecturalRegMap_18 | (6'h1e == architecturalRegMap_17 | (6'h1e ==
    architecturalRegMap_16 | _GEN_3152)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5073 = 6'h1f == architecturalRegMap_30 | (6'h1f == architecturalRegMap_29 | (6'h1f ==
    architecturalRegMap_28 | (6'h1f == architecturalRegMap_27 | (6'h1f == architecturalRegMap_26 | (6'h1f ==
    architecturalRegMap_25 | (6'h1f == architecturalRegMap_24 | (6'h1f == architecturalRegMap_23 | (6'h1f ==
    architecturalRegMap_22 | (6'h1f == architecturalRegMap_21 | (6'h1f == architecturalRegMap_20 | (6'h1f ==
    architecturalRegMap_19 | (6'h1f == architecturalRegMap_18 | (6'h1f == architecturalRegMap_17 | (6'h1f ==
    architecturalRegMap_16 | _GEN_3153)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5074 = 6'h20 == architecturalRegMap_30 | (6'h20 == architecturalRegMap_29 | (6'h20 ==
    architecturalRegMap_28 | (6'h20 == architecturalRegMap_27 | (6'h20 == architecturalRegMap_26 | (6'h20 ==
    architecturalRegMap_25 | (6'h20 == architecturalRegMap_24 | (6'h20 == architecturalRegMap_23 | (6'h20 ==
    architecturalRegMap_22 | (6'h20 == architecturalRegMap_21 | (6'h20 == architecturalRegMap_20 | (6'h20 ==
    architecturalRegMap_19 | (6'h20 == architecturalRegMap_18 | (6'h20 == architecturalRegMap_17 | (6'h20 ==
    architecturalRegMap_16 | _GEN_3154)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5075 = 6'h21 == architecturalRegMap_30 | (6'h21 == architecturalRegMap_29 | (6'h21 ==
    architecturalRegMap_28 | (6'h21 == architecturalRegMap_27 | (6'h21 == architecturalRegMap_26 | (6'h21 ==
    architecturalRegMap_25 | (6'h21 == architecturalRegMap_24 | (6'h21 == architecturalRegMap_23 | (6'h21 ==
    architecturalRegMap_22 | (6'h21 == architecturalRegMap_21 | (6'h21 == architecturalRegMap_20 | (6'h21 ==
    architecturalRegMap_19 | (6'h21 == architecturalRegMap_18 | (6'h21 == architecturalRegMap_17 | (6'h21 ==
    architecturalRegMap_16 | _GEN_3155)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5076 = 6'h22 == architecturalRegMap_30 | (6'h22 == architecturalRegMap_29 | (6'h22 ==
    architecturalRegMap_28 | (6'h22 == architecturalRegMap_27 | (6'h22 == architecturalRegMap_26 | (6'h22 ==
    architecturalRegMap_25 | (6'h22 == architecturalRegMap_24 | (6'h22 == architecturalRegMap_23 | (6'h22 ==
    architecturalRegMap_22 | (6'h22 == architecturalRegMap_21 | (6'h22 == architecturalRegMap_20 | (6'h22 ==
    architecturalRegMap_19 | (6'h22 == architecturalRegMap_18 | (6'h22 == architecturalRegMap_17 | (6'h22 ==
    architecturalRegMap_16 | _GEN_3156)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5077 = 6'h23 == architecturalRegMap_30 | (6'h23 == architecturalRegMap_29 | (6'h23 ==
    architecturalRegMap_28 | (6'h23 == architecturalRegMap_27 | (6'h23 == architecturalRegMap_26 | (6'h23 ==
    architecturalRegMap_25 | (6'h23 == architecturalRegMap_24 | (6'h23 == architecturalRegMap_23 | (6'h23 ==
    architecturalRegMap_22 | (6'h23 == architecturalRegMap_21 | (6'h23 == architecturalRegMap_20 | (6'h23 ==
    architecturalRegMap_19 | (6'h23 == architecturalRegMap_18 | (6'h23 == architecturalRegMap_17 | (6'h23 ==
    architecturalRegMap_16 | _GEN_3157)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5078 = 6'h24 == architecturalRegMap_30 | (6'h24 == architecturalRegMap_29 | (6'h24 ==
    architecturalRegMap_28 | (6'h24 == architecturalRegMap_27 | (6'h24 == architecturalRegMap_26 | (6'h24 ==
    architecturalRegMap_25 | (6'h24 == architecturalRegMap_24 | (6'h24 == architecturalRegMap_23 | (6'h24 ==
    architecturalRegMap_22 | (6'h24 == architecturalRegMap_21 | (6'h24 == architecturalRegMap_20 | (6'h24 ==
    architecturalRegMap_19 | (6'h24 == architecturalRegMap_18 | (6'h24 == architecturalRegMap_17 | (6'h24 ==
    architecturalRegMap_16 | _GEN_3158)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5079 = 6'h25 == architecturalRegMap_30 | (6'h25 == architecturalRegMap_29 | (6'h25 ==
    architecturalRegMap_28 | (6'h25 == architecturalRegMap_27 | (6'h25 == architecturalRegMap_26 | (6'h25 ==
    architecturalRegMap_25 | (6'h25 == architecturalRegMap_24 | (6'h25 == architecturalRegMap_23 | (6'h25 ==
    architecturalRegMap_22 | (6'h25 == architecturalRegMap_21 | (6'h25 == architecturalRegMap_20 | (6'h25 ==
    architecturalRegMap_19 | (6'h25 == architecturalRegMap_18 | (6'h25 == architecturalRegMap_17 | (6'h25 ==
    architecturalRegMap_16 | _GEN_3159)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5080 = 6'h26 == architecturalRegMap_30 | (6'h26 == architecturalRegMap_29 | (6'h26 ==
    architecturalRegMap_28 | (6'h26 == architecturalRegMap_27 | (6'h26 == architecturalRegMap_26 | (6'h26 ==
    architecturalRegMap_25 | (6'h26 == architecturalRegMap_24 | (6'h26 == architecturalRegMap_23 | (6'h26 ==
    architecturalRegMap_22 | (6'h26 == architecturalRegMap_21 | (6'h26 == architecturalRegMap_20 | (6'h26 ==
    architecturalRegMap_19 | (6'h26 == architecturalRegMap_18 | (6'h26 == architecturalRegMap_17 | (6'h26 ==
    architecturalRegMap_16 | _GEN_3160)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5081 = 6'h27 == architecturalRegMap_30 | (6'h27 == architecturalRegMap_29 | (6'h27 ==
    architecturalRegMap_28 | (6'h27 == architecturalRegMap_27 | (6'h27 == architecturalRegMap_26 | (6'h27 ==
    architecturalRegMap_25 | (6'h27 == architecturalRegMap_24 | (6'h27 == architecturalRegMap_23 | (6'h27 ==
    architecturalRegMap_22 | (6'h27 == architecturalRegMap_21 | (6'h27 == architecturalRegMap_20 | (6'h27 ==
    architecturalRegMap_19 | (6'h27 == architecturalRegMap_18 | (6'h27 == architecturalRegMap_17 | (6'h27 ==
    architecturalRegMap_16 | _GEN_3161)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5082 = 6'h28 == architecturalRegMap_30 | (6'h28 == architecturalRegMap_29 | (6'h28 ==
    architecturalRegMap_28 | (6'h28 == architecturalRegMap_27 | (6'h28 == architecturalRegMap_26 | (6'h28 ==
    architecturalRegMap_25 | (6'h28 == architecturalRegMap_24 | (6'h28 == architecturalRegMap_23 | (6'h28 ==
    architecturalRegMap_22 | (6'h28 == architecturalRegMap_21 | (6'h28 == architecturalRegMap_20 | (6'h28 ==
    architecturalRegMap_19 | (6'h28 == architecturalRegMap_18 | (6'h28 == architecturalRegMap_17 | (6'h28 ==
    architecturalRegMap_16 | _GEN_3162)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5083 = 6'h29 == architecturalRegMap_30 | (6'h29 == architecturalRegMap_29 | (6'h29 ==
    architecturalRegMap_28 | (6'h29 == architecturalRegMap_27 | (6'h29 == architecturalRegMap_26 | (6'h29 ==
    architecturalRegMap_25 | (6'h29 == architecturalRegMap_24 | (6'h29 == architecturalRegMap_23 | (6'h29 ==
    architecturalRegMap_22 | (6'h29 == architecturalRegMap_21 | (6'h29 == architecturalRegMap_20 | (6'h29 ==
    architecturalRegMap_19 | (6'h29 == architecturalRegMap_18 | (6'h29 == architecturalRegMap_17 | (6'h29 ==
    architecturalRegMap_16 | _GEN_3163)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5084 = 6'h2a == architecturalRegMap_30 | (6'h2a == architecturalRegMap_29 | (6'h2a ==
    architecturalRegMap_28 | (6'h2a == architecturalRegMap_27 | (6'h2a == architecturalRegMap_26 | (6'h2a ==
    architecturalRegMap_25 | (6'h2a == architecturalRegMap_24 | (6'h2a == architecturalRegMap_23 | (6'h2a ==
    architecturalRegMap_22 | (6'h2a == architecturalRegMap_21 | (6'h2a == architecturalRegMap_20 | (6'h2a ==
    architecturalRegMap_19 | (6'h2a == architecturalRegMap_18 | (6'h2a == architecturalRegMap_17 | (6'h2a ==
    architecturalRegMap_16 | _GEN_3164)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5085 = 6'h2b == architecturalRegMap_30 | (6'h2b == architecturalRegMap_29 | (6'h2b ==
    architecturalRegMap_28 | (6'h2b == architecturalRegMap_27 | (6'h2b == architecturalRegMap_26 | (6'h2b ==
    architecturalRegMap_25 | (6'h2b == architecturalRegMap_24 | (6'h2b == architecturalRegMap_23 | (6'h2b ==
    architecturalRegMap_22 | (6'h2b == architecturalRegMap_21 | (6'h2b == architecturalRegMap_20 | (6'h2b ==
    architecturalRegMap_19 | (6'h2b == architecturalRegMap_18 | (6'h2b == architecturalRegMap_17 | (6'h2b ==
    architecturalRegMap_16 | _GEN_3165)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5086 = 6'h2c == architecturalRegMap_30 | (6'h2c == architecturalRegMap_29 | (6'h2c ==
    architecturalRegMap_28 | (6'h2c == architecturalRegMap_27 | (6'h2c == architecturalRegMap_26 | (6'h2c ==
    architecturalRegMap_25 | (6'h2c == architecturalRegMap_24 | (6'h2c == architecturalRegMap_23 | (6'h2c ==
    architecturalRegMap_22 | (6'h2c == architecturalRegMap_21 | (6'h2c == architecturalRegMap_20 | (6'h2c ==
    architecturalRegMap_19 | (6'h2c == architecturalRegMap_18 | (6'h2c == architecturalRegMap_17 | (6'h2c ==
    architecturalRegMap_16 | _GEN_3166)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5087 = 6'h2d == architecturalRegMap_30 | (6'h2d == architecturalRegMap_29 | (6'h2d ==
    architecturalRegMap_28 | (6'h2d == architecturalRegMap_27 | (6'h2d == architecturalRegMap_26 | (6'h2d ==
    architecturalRegMap_25 | (6'h2d == architecturalRegMap_24 | (6'h2d == architecturalRegMap_23 | (6'h2d ==
    architecturalRegMap_22 | (6'h2d == architecturalRegMap_21 | (6'h2d == architecturalRegMap_20 | (6'h2d ==
    architecturalRegMap_19 | (6'h2d == architecturalRegMap_18 | (6'h2d == architecturalRegMap_17 | (6'h2d ==
    architecturalRegMap_16 | _GEN_3167)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5088 = 6'h2e == architecturalRegMap_30 | (6'h2e == architecturalRegMap_29 | (6'h2e ==
    architecturalRegMap_28 | (6'h2e == architecturalRegMap_27 | (6'h2e == architecturalRegMap_26 | (6'h2e ==
    architecturalRegMap_25 | (6'h2e == architecturalRegMap_24 | (6'h2e == architecturalRegMap_23 | (6'h2e ==
    architecturalRegMap_22 | (6'h2e == architecturalRegMap_21 | (6'h2e == architecturalRegMap_20 | (6'h2e ==
    architecturalRegMap_19 | (6'h2e == architecturalRegMap_18 | (6'h2e == architecturalRegMap_17 | (6'h2e ==
    architecturalRegMap_16 | _GEN_3168)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5089 = 6'h2f == architecturalRegMap_30 | (6'h2f == architecturalRegMap_29 | (6'h2f ==
    architecturalRegMap_28 | (6'h2f == architecturalRegMap_27 | (6'h2f == architecturalRegMap_26 | (6'h2f ==
    architecturalRegMap_25 | (6'h2f == architecturalRegMap_24 | (6'h2f == architecturalRegMap_23 | (6'h2f ==
    architecturalRegMap_22 | (6'h2f == architecturalRegMap_21 | (6'h2f == architecturalRegMap_20 | (6'h2f ==
    architecturalRegMap_19 | (6'h2f == architecturalRegMap_18 | (6'h2f == architecturalRegMap_17 | (6'h2f ==
    architecturalRegMap_16 | _GEN_3169)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5090 = 6'h30 == architecturalRegMap_30 | (6'h30 == architecturalRegMap_29 | (6'h30 ==
    architecturalRegMap_28 | (6'h30 == architecturalRegMap_27 | (6'h30 == architecturalRegMap_26 | (6'h30 ==
    architecturalRegMap_25 | (6'h30 == architecturalRegMap_24 | (6'h30 == architecturalRegMap_23 | (6'h30 ==
    architecturalRegMap_22 | (6'h30 == architecturalRegMap_21 | (6'h30 == architecturalRegMap_20 | (6'h30 ==
    architecturalRegMap_19 | (6'h30 == architecturalRegMap_18 | (6'h30 == architecturalRegMap_17 | (6'h30 ==
    architecturalRegMap_16 | _GEN_3170)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5091 = 6'h31 == architecturalRegMap_30 | (6'h31 == architecturalRegMap_29 | (6'h31 ==
    architecturalRegMap_28 | (6'h31 == architecturalRegMap_27 | (6'h31 == architecturalRegMap_26 | (6'h31 ==
    architecturalRegMap_25 | (6'h31 == architecturalRegMap_24 | (6'h31 == architecturalRegMap_23 | (6'h31 ==
    architecturalRegMap_22 | (6'h31 == architecturalRegMap_21 | (6'h31 == architecturalRegMap_20 | (6'h31 ==
    architecturalRegMap_19 | (6'h31 == architecturalRegMap_18 | (6'h31 == architecturalRegMap_17 | (6'h31 ==
    architecturalRegMap_16 | _GEN_3171)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5092 = 6'h32 == architecturalRegMap_30 | (6'h32 == architecturalRegMap_29 | (6'h32 ==
    architecturalRegMap_28 | (6'h32 == architecturalRegMap_27 | (6'h32 == architecturalRegMap_26 | (6'h32 ==
    architecturalRegMap_25 | (6'h32 == architecturalRegMap_24 | (6'h32 == architecturalRegMap_23 | (6'h32 ==
    architecturalRegMap_22 | (6'h32 == architecturalRegMap_21 | (6'h32 == architecturalRegMap_20 | (6'h32 ==
    architecturalRegMap_19 | (6'h32 == architecturalRegMap_18 | (6'h32 == architecturalRegMap_17 | (6'h32 ==
    architecturalRegMap_16 | _GEN_3172)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5093 = 6'h33 == architecturalRegMap_30 | (6'h33 == architecturalRegMap_29 | (6'h33 ==
    architecturalRegMap_28 | (6'h33 == architecturalRegMap_27 | (6'h33 == architecturalRegMap_26 | (6'h33 ==
    architecturalRegMap_25 | (6'h33 == architecturalRegMap_24 | (6'h33 == architecturalRegMap_23 | (6'h33 ==
    architecturalRegMap_22 | (6'h33 == architecturalRegMap_21 | (6'h33 == architecturalRegMap_20 | (6'h33 ==
    architecturalRegMap_19 | (6'h33 == architecturalRegMap_18 | (6'h33 == architecturalRegMap_17 | (6'h33 ==
    architecturalRegMap_16 | _GEN_3173)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5094 = 6'h34 == architecturalRegMap_30 | (6'h34 == architecturalRegMap_29 | (6'h34 ==
    architecturalRegMap_28 | (6'h34 == architecturalRegMap_27 | (6'h34 == architecturalRegMap_26 | (6'h34 ==
    architecturalRegMap_25 | (6'h34 == architecturalRegMap_24 | (6'h34 == architecturalRegMap_23 | (6'h34 ==
    architecturalRegMap_22 | (6'h34 == architecturalRegMap_21 | (6'h34 == architecturalRegMap_20 | (6'h34 ==
    architecturalRegMap_19 | (6'h34 == architecturalRegMap_18 | (6'h34 == architecturalRegMap_17 | (6'h34 ==
    architecturalRegMap_16 | _GEN_3174)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5095 = 6'h35 == architecturalRegMap_30 | (6'h35 == architecturalRegMap_29 | (6'h35 ==
    architecturalRegMap_28 | (6'h35 == architecturalRegMap_27 | (6'h35 == architecturalRegMap_26 | (6'h35 ==
    architecturalRegMap_25 | (6'h35 == architecturalRegMap_24 | (6'h35 == architecturalRegMap_23 | (6'h35 ==
    architecturalRegMap_22 | (6'h35 == architecturalRegMap_21 | (6'h35 == architecturalRegMap_20 | (6'h35 ==
    architecturalRegMap_19 | (6'h35 == architecturalRegMap_18 | (6'h35 == architecturalRegMap_17 | (6'h35 ==
    architecturalRegMap_16 | _GEN_3175)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5096 = 6'h36 == architecturalRegMap_30 | (6'h36 == architecturalRegMap_29 | (6'h36 ==
    architecturalRegMap_28 | (6'h36 == architecturalRegMap_27 | (6'h36 == architecturalRegMap_26 | (6'h36 ==
    architecturalRegMap_25 | (6'h36 == architecturalRegMap_24 | (6'h36 == architecturalRegMap_23 | (6'h36 ==
    architecturalRegMap_22 | (6'h36 == architecturalRegMap_21 | (6'h36 == architecturalRegMap_20 | (6'h36 ==
    architecturalRegMap_19 | (6'h36 == architecturalRegMap_18 | (6'h36 == architecturalRegMap_17 | (6'h36 ==
    architecturalRegMap_16 | _GEN_3176)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5097 = 6'h37 == architecturalRegMap_30 | (6'h37 == architecturalRegMap_29 | (6'h37 ==
    architecturalRegMap_28 | (6'h37 == architecturalRegMap_27 | (6'h37 == architecturalRegMap_26 | (6'h37 ==
    architecturalRegMap_25 | (6'h37 == architecturalRegMap_24 | (6'h37 == architecturalRegMap_23 | (6'h37 ==
    architecturalRegMap_22 | (6'h37 == architecturalRegMap_21 | (6'h37 == architecturalRegMap_20 | (6'h37 ==
    architecturalRegMap_19 | (6'h37 == architecturalRegMap_18 | (6'h37 == architecturalRegMap_17 | (6'h37 ==
    architecturalRegMap_16 | _GEN_3177)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5098 = 6'h38 == architecturalRegMap_30 | (6'h38 == architecturalRegMap_29 | (6'h38 ==
    architecturalRegMap_28 | (6'h38 == architecturalRegMap_27 | (6'h38 == architecturalRegMap_26 | (6'h38 ==
    architecturalRegMap_25 | (6'h38 == architecturalRegMap_24 | (6'h38 == architecturalRegMap_23 | (6'h38 ==
    architecturalRegMap_22 | (6'h38 == architecturalRegMap_21 | (6'h38 == architecturalRegMap_20 | (6'h38 ==
    architecturalRegMap_19 | (6'h38 == architecturalRegMap_18 | (6'h38 == architecturalRegMap_17 | (6'h38 ==
    architecturalRegMap_16 | _GEN_3178)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5099 = 6'h39 == architecturalRegMap_30 | (6'h39 == architecturalRegMap_29 | (6'h39 ==
    architecturalRegMap_28 | (6'h39 == architecturalRegMap_27 | (6'h39 == architecturalRegMap_26 | (6'h39 ==
    architecturalRegMap_25 | (6'h39 == architecturalRegMap_24 | (6'h39 == architecturalRegMap_23 | (6'h39 ==
    architecturalRegMap_22 | (6'h39 == architecturalRegMap_21 | (6'h39 == architecturalRegMap_20 | (6'h39 ==
    architecturalRegMap_19 | (6'h39 == architecturalRegMap_18 | (6'h39 == architecturalRegMap_17 | (6'h39 ==
    architecturalRegMap_16 | _GEN_3179)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5100 = 6'h3a == architecturalRegMap_30 | (6'h3a == architecturalRegMap_29 | (6'h3a ==
    architecturalRegMap_28 | (6'h3a == architecturalRegMap_27 | (6'h3a == architecturalRegMap_26 | (6'h3a ==
    architecturalRegMap_25 | (6'h3a == architecturalRegMap_24 | (6'h3a == architecturalRegMap_23 | (6'h3a ==
    architecturalRegMap_22 | (6'h3a == architecturalRegMap_21 | (6'h3a == architecturalRegMap_20 | (6'h3a ==
    architecturalRegMap_19 | (6'h3a == architecturalRegMap_18 | (6'h3a == architecturalRegMap_17 | (6'h3a ==
    architecturalRegMap_16 | _GEN_3180)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5101 = 6'h3b == architecturalRegMap_30 | (6'h3b == architecturalRegMap_29 | (6'h3b ==
    architecturalRegMap_28 | (6'h3b == architecturalRegMap_27 | (6'h3b == architecturalRegMap_26 | (6'h3b ==
    architecturalRegMap_25 | (6'h3b == architecturalRegMap_24 | (6'h3b == architecturalRegMap_23 | (6'h3b ==
    architecturalRegMap_22 | (6'h3b == architecturalRegMap_21 | (6'h3b == architecturalRegMap_20 | (6'h3b ==
    architecturalRegMap_19 | (6'h3b == architecturalRegMap_18 | (6'h3b == architecturalRegMap_17 | (6'h3b ==
    architecturalRegMap_16 | _GEN_3181)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5102 = 6'h3c == architecturalRegMap_30 | (6'h3c == architecturalRegMap_29 | (6'h3c ==
    architecturalRegMap_28 | (6'h3c == architecturalRegMap_27 | (6'h3c == architecturalRegMap_26 | (6'h3c ==
    architecturalRegMap_25 | (6'h3c == architecturalRegMap_24 | (6'h3c == architecturalRegMap_23 | (6'h3c ==
    architecturalRegMap_22 | (6'h3c == architecturalRegMap_21 | (6'h3c == architecturalRegMap_20 | (6'h3c ==
    architecturalRegMap_19 | (6'h3c == architecturalRegMap_18 | (6'h3c == architecturalRegMap_17 | (6'h3c ==
    architecturalRegMap_16 | _GEN_3182)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5103 = 6'h3d == architecturalRegMap_30 | (6'h3d == architecturalRegMap_29 | (6'h3d ==
    architecturalRegMap_28 | (6'h3d == architecturalRegMap_27 | (6'h3d == architecturalRegMap_26 | (6'h3d ==
    architecturalRegMap_25 | (6'h3d == architecturalRegMap_24 | (6'h3d == architecturalRegMap_23 | (6'h3d ==
    architecturalRegMap_22 | (6'h3d == architecturalRegMap_21 | (6'h3d == architecturalRegMap_20 | (6'h3d ==
    architecturalRegMap_19 | (6'h3d == architecturalRegMap_18 | (6'h3d == architecturalRegMap_17 | (6'h3d ==
    architecturalRegMap_16 | _GEN_3183)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5104 = 6'h3e == architecturalRegMap_30 | (6'h3e == architecturalRegMap_29 | (6'h3e ==
    architecturalRegMap_28 | (6'h3e == architecturalRegMap_27 | (6'h3e == architecturalRegMap_26 | (6'h3e ==
    architecturalRegMap_25 | (6'h3e == architecturalRegMap_24 | (6'h3e == architecturalRegMap_23 | (6'h3e ==
    architecturalRegMap_22 | (6'h3e == architecturalRegMap_21 | (6'h3e == architecturalRegMap_20 | (6'h3e ==
    architecturalRegMap_19 | (6'h3e == architecturalRegMap_18 | (6'h3e == architecturalRegMap_17 | (6'h3e ==
    architecturalRegMap_16 | _GEN_3184)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5105 = 6'h3f == architecturalRegMap_30 | (6'h3f == architecturalRegMap_29 | (6'h3f ==
    architecturalRegMap_28 | (6'h3f == architecturalRegMap_27 | (6'h3f == architecturalRegMap_26 | (6'h3f ==
    architecturalRegMap_25 | (6'h3f == architecturalRegMap_24 | (6'h3f == architecturalRegMap_23 | (6'h3f ==
    architecturalRegMap_22 | (6'h3f == architecturalRegMap_21 | (6'h3f == architecturalRegMap_20 | (6'h3f ==
    architecturalRegMap_19 | (6'h3f == architecturalRegMap_18 | (6'h3f == architecturalRegMap_17 | (6'h3f ==
    architecturalRegMap_16 | _GEN_3185)))))))))))))); // @[decode.scala 392:{47,47}]
  wire  _GEN_5106 = 6'h0 == architecturalRegMap_30 ? 1'h0 : _GEN_4978; // @[decode.scala 393:{46,46}]
  wire  _GEN_5107 = 6'h1 == architecturalRegMap_30 ? 1'h0 : _GEN_4979; // @[decode.scala 393:{46,46}]
  wire  _GEN_5108 = 6'h2 == architecturalRegMap_30 ? 1'h0 : _GEN_4980; // @[decode.scala 393:{46,46}]
  wire  _GEN_5109 = 6'h3 == architecturalRegMap_30 ? 1'h0 : _GEN_4981; // @[decode.scala 393:{46,46}]
  wire  _GEN_5110 = 6'h4 == architecturalRegMap_30 ? 1'h0 : _GEN_4982; // @[decode.scala 393:{46,46}]
  wire  _GEN_5111 = 6'h5 == architecturalRegMap_30 ? 1'h0 : _GEN_4983; // @[decode.scala 393:{46,46}]
  wire  _GEN_5112 = 6'h6 == architecturalRegMap_30 ? 1'h0 : _GEN_4984; // @[decode.scala 393:{46,46}]
  wire  _GEN_5113 = 6'h7 == architecturalRegMap_30 ? 1'h0 : _GEN_4985; // @[decode.scala 393:{46,46}]
  wire  _GEN_5114 = 6'h8 == architecturalRegMap_30 ? 1'h0 : _GEN_4986; // @[decode.scala 393:{46,46}]
  wire  _GEN_5115 = 6'h9 == architecturalRegMap_30 ? 1'h0 : _GEN_4987; // @[decode.scala 393:{46,46}]
  wire  _GEN_5116 = 6'ha == architecturalRegMap_30 ? 1'h0 : _GEN_4988; // @[decode.scala 393:{46,46}]
  wire  _GEN_5117 = 6'hb == architecturalRegMap_30 ? 1'h0 : _GEN_4989; // @[decode.scala 393:{46,46}]
  wire  _GEN_5118 = 6'hc == architecturalRegMap_30 ? 1'h0 : _GEN_4990; // @[decode.scala 393:{46,46}]
  wire  _GEN_5119 = 6'hd == architecturalRegMap_30 ? 1'h0 : _GEN_4991; // @[decode.scala 393:{46,46}]
  wire  _GEN_5120 = 6'he == architecturalRegMap_30 ? 1'h0 : _GEN_4992; // @[decode.scala 393:{46,46}]
  wire  _GEN_5121 = 6'hf == architecturalRegMap_30 ? 1'h0 : _GEN_4993; // @[decode.scala 393:{46,46}]
  wire  _GEN_5122 = 6'h10 == architecturalRegMap_30 ? 1'h0 : _GEN_4994; // @[decode.scala 393:{46,46}]
  wire  _GEN_5123 = 6'h11 == architecturalRegMap_30 ? 1'h0 : _GEN_4995; // @[decode.scala 393:{46,46}]
  wire  _GEN_5124 = 6'h12 == architecturalRegMap_30 ? 1'h0 : _GEN_4996; // @[decode.scala 393:{46,46}]
  wire  _GEN_5125 = 6'h13 == architecturalRegMap_30 ? 1'h0 : _GEN_4997; // @[decode.scala 393:{46,46}]
  wire  _GEN_5126 = 6'h14 == architecturalRegMap_30 ? 1'h0 : _GEN_4998; // @[decode.scala 393:{46,46}]
  wire  _GEN_5127 = 6'h15 == architecturalRegMap_30 ? 1'h0 : _GEN_4999; // @[decode.scala 393:{46,46}]
  wire  _GEN_5128 = 6'h16 == architecturalRegMap_30 ? 1'h0 : _GEN_5000; // @[decode.scala 393:{46,46}]
  wire  _GEN_5129 = 6'h17 == architecturalRegMap_30 ? 1'h0 : _GEN_5001; // @[decode.scala 393:{46,46}]
  wire  _GEN_5130 = 6'h18 == architecturalRegMap_30 ? 1'h0 : _GEN_5002; // @[decode.scala 393:{46,46}]
  wire  _GEN_5131 = 6'h19 == architecturalRegMap_30 ? 1'h0 : _GEN_5003; // @[decode.scala 393:{46,46}]
  wire  _GEN_5132 = 6'h1a == architecturalRegMap_30 ? 1'h0 : _GEN_5004; // @[decode.scala 393:{46,46}]
  wire  _GEN_5133 = 6'h1b == architecturalRegMap_30 ? 1'h0 : _GEN_5005; // @[decode.scala 393:{46,46}]
  wire  _GEN_5134 = 6'h1c == architecturalRegMap_30 ? 1'h0 : _GEN_5006; // @[decode.scala 393:{46,46}]
  wire  _GEN_5135 = 6'h1d == architecturalRegMap_30 ? 1'h0 : _GEN_5007; // @[decode.scala 393:{46,46}]
  wire  _GEN_5136 = 6'h1e == architecturalRegMap_30 ? 1'h0 : _GEN_5008; // @[decode.scala 393:{46,46}]
  wire  _GEN_5137 = 6'h1f == architecturalRegMap_30 ? 1'h0 : _GEN_5009; // @[decode.scala 393:{46,46}]
  wire  _GEN_5138 = 6'h20 == architecturalRegMap_30 ? 1'h0 : _GEN_5010; // @[decode.scala 393:{46,46}]
  wire  _GEN_5139 = 6'h21 == architecturalRegMap_30 ? 1'h0 : _GEN_5011; // @[decode.scala 393:{46,46}]
  wire  _GEN_5140 = 6'h22 == architecturalRegMap_30 ? 1'h0 : _GEN_5012; // @[decode.scala 393:{46,46}]
  wire  _GEN_5141 = 6'h23 == architecturalRegMap_30 ? 1'h0 : _GEN_5013; // @[decode.scala 393:{46,46}]
  wire  _GEN_5142 = 6'h24 == architecturalRegMap_30 ? 1'h0 : _GEN_5014; // @[decode.scala 393:{46,46}]
  wire  _GEN_5143 = 6'h25 == architecturalRegMap_30 ? 1'h0 : _GEN_5015; // @[decode.scala 393:{46,46}]
  wire  _GEN_5144 = 6'h26 == architecturalRegMap_30 ? 1'h0 : _GEN_5016; // @[decode.scala 393:{46,46}]
  wire  _GEN_5145 = 6'h27 == architecturalRegMap_30 ? 1'h0 : _GEN_5017; // @[decode.scala 393:{46,46}]
  wire  _GEN_5146 = 6'h28 == architecturalRegMap_30 ? 1'h0 : _GEN_5018; // @[decode.scala 393:{46,46}]
  wire  _GEN_5147 = 6'h29 == architecturalRegMap_30 ? 1'h0 : _GEN_5019; // @[decode.scala 393:{46,46}]
  wire  _GEN_5148 = 6'h2a == architecturalRegMap_30 ? 1'h0 : _GEN_5020; // @[decode.scala 393:{46,46}]
  wire  _GEN_5149 = 6'h2b == architecturalRegMap_30 ? 1'h0 : _GEN_5021; // @[decode.scala 393:{46,46}]
  wire  _GEN_5150 = 6'h2c == architecturalRegMap_30 ? 1'h0 : _GEN_5022; // @[decode.scala 393:{46,46}]
  wire  _GEN_5151 = 6'h2d == architecturalRegMap_30 ? 1'h0 : _GEN_5023; // @[decode.scala 393:{46,46}]
  wire  _GEN_5152 = 6'h2e == architecturalRegMap_30 ? 1'h0 : _GEN_5024; // @[decode.scala 393:{46,46}]
  wire  _GEN_5153 = 6'h2f == architecturalRegMap_30 ? 1'h0 : _GEN_5025; // @[decode.scala 393:{46,46}]
  wire  _GEN_5154 = 6'h30 == architecturalRegMap_30 ? 1'h0 : _GEN_5026; // @[decode.scala 393:{46,46}]
  wire  _GEN_5155 = 6'h31 == architecturalRegMap_30 ? 1'h0 : _GEN_5027; // @[decode.scala 393:{46,46}]
  wire  _GEN_5156 = 6'h32 == architecturalRegMap_30 ? 1'h0 : _GEN_5028; // @[decode.scala 393:{46,46}]
  wire  _GEN_5157 = 6'h33 == architecturalRegMap_30 ? 1'h0 : _GEN_5029; // @[decode.scala 393:{46,46}]
  wire  _GEN_5158 = 6'h34 == architecturalRegMap_30 ? 1'h0 : _GEN_5030; // @[decode.scala 393:{46,46}]
  wire  _GEN_5159 = 6'h35 == architecturalRegMap_30 ? 1'h0 : _GEN_5031; // @[decode.scala 393:{46,46}]
  wire  _GEN_5160 = 6'h36 == architecturalRegMap_30 ? 1'h0 : _GEN_5032; // @[decode.scala 393:{46,46}]
  wire  _GEN_5161 = 6'h37 == architecturalRegMap_30 ? 1'h0 : _GEN_5033; // @[decode.scala 393:{46,46}]
  wire  _GEN_5162 = 6'h38 == architecturalRegMap_30 ? 1'h0 : _GEN_5034; // @[decode.scala 393:{46,46}]
  wire  _GEN_5163 = 6'h39 == architecturalRegMap_30 ? 1'h0 : _GEN_5035; // @[decode.scala 393:{46,46}]
  wire  _GEN_5164 = 6'h3a == architecturalRegMap_30 ? 1'h0 : _GEN_5036; // @[decode.scala 393:{46,46}]
  wire  _GEN_5165 = 6'h3b == architecturalRegMap_30 ? 1'h0 : _GEN_5037; // @[decode.scala 393:{46,46}]
  wire  _GEN_5166 = 6'h3c == architecturalRegMap_30 ? 1'h0 : _GEN_5038; // @[decode.scala 393:{46,46}]
  wire  _GEN_5167 = 6'h3d == architecturalRegMap_30 ? 1'h0 : _GEN_5039; // @[decode.scala 393:{46,46}]
  wire  _GEN_5168 = 6'h3e == architecturalRegMap_30 ? 1'h0 : _GEN_5040; // @[decode.scala 393:{46,46}]
  wire  _GEN_5170 = 6'h0 == architecturalRegMap_31 | _GEN_5042; // @[decode.scala 392:{47,47}]
  wire  _GEN_5171 = 6'h1 == architecturalRegMap_31 | _GEN_5043; // @[decode.scala 392:{47,47}]
  wire  _GEN_5172 = 6'h2 == architecturalRegMap_31 | _GEN_5044; // @[decode.scala 392:{47,47}]
  wire  _GEN_5173 = 6'h3 == architecturalRegMap_31 | _GEN_5045; // @[decode.scala 392:{47,47}]
  wire  _GEN_5174 = 6'h4 == architecturalRegMap_31 | _GEN_5046; // @[decode.scala 392:{47,47}]
  wire  _GEN_5175 = 6'h5 == architecturalRegMap_31 | _GEN_5047; // @[decode.scala 392:{47,47}]
  wire  _GEN_5176 = 6'h6 == architecturalRegMap_31 | _GEN_5048; // @[decode.scala 392:{47,47}]
  wire  _GEN_5177 = 6'h7 == architecturalRegMap_31 | _GEN_5049; // @[decode.scala 392:{47,47}]
  wire  _GEN_5178 = 6'h8 == architecturalRegMap_31 | _GEN_5050; // @[decode.scala 392:{47,47}]
  wire  _GEN_5179 = 6'h9 == architecturalRegMap_31 | _GEN_5051; // @[decode.scala 392:{47,47}]
  wire  _GEN_5180 = 6'ha == architecturalRegMap_31 | _GEN_5052; // @[decode.scala 392:{47,47}]
  wire  _GEN_5181 = 6'hb == architecturalRegMap_31 | _GEN_5053; // @[decode.scala 392:{47,47}]
  wire  _GEN_5182 = 6'hc == architecturalRegMap_31 | _GEN_5054; // @[decode.scala 392:{47,47}]
  wire  _GEN_5183 = 6'hd == architecturalRegMap_31 | _GEN_5055; // @[decode.scala 392:{47,47}]
  wire  _GEN_5184 = 6'he == architecturalRegMap_31 | _GEN_5056; // @[decode.scala 392:{47,47}]
  wire  _GEN_5185 = 6'hf == architecturalRegMap_31 | _GEN_5057; // @[decode.scala 392:{47,47}]
  wire  _GEN_5186 = 6'h10 == architecturalRegMap_31 | _GEN_5058; // @[decode.scala 392:{47,47}]
  wire  _GEN_5187 = 6'h11 == architecturalRegMap_31 | _GEN_5059; // @[decode.scala 392:{47,47}]
  wire  _GEN_5188 = 6'h12 == architecturalRegMap_31 | _GEN_5060; // @[decode.scala 392:{47,47}]
  wire  _GEN_5189 = 6'h13 == architecturalRegMap_31 | _GEN_5061; // @[decode.scala 392:{47,47}]
  wire  _GEN_5190 = 6'h14 == architecturalRegMap_31 | _GEN_5062; // @[decode.scala 392:{47,47}]
  wire  _GEN_5191 = 6'h15 == architecturalRegMap_31 | _GEN_5063; // @[decode.scala 392:{47,47}]
  wire  _GEN_5192 = 6'h16 == architecturalRegMap_31 | _GEN_5064; // @[decode.scala 392:{47,47}]
  wire  _GEN_5193 = 6'h17 == architecturalRegMap_31 | _GEN_5065; // @[decode.scala 392:{47,47}]
  wire  _GEN_5194 = 6'h18 == architecturalRegMap_31 | _GEN_5066; // @[decode.scala 392:{47,47}]
  wire  _GEN_5195 = 6'h19 == architecturalRegMap_31 | _GEN_5067; // @[decode.scala 392:{47,47}]
  wire  _GEN_5196 = 6'h1a == architecturalRegMap_31 | _GEN_5068; // @[decode.scala 392:{47,47}]
  wire  _GEN_5197 = 6'h1b == architecturalRegMap_31 | _GEN_5069; // @[decode.scala 392:{47,47}]
  wire  _GEN_5198 = 6'h1c == architecturalRegMap_31 | _GEN_5070; // @[decode.scala 392:{47,47}]
  wire  _GEN_5199 = 6'h1d == architecturalRegMap_31 | _GEN_5071; // @[decode.scala 392:{47,47}]
  wire  _GEN_5200 = 6'h1e == architecturalRegMap_31 | _GEN_5072; // @[decode.scala 392:{47,47}]
  wire  _GEN_5201 = 6'h1f == architecturalRegMap_31 | _GEN_5073; // @[decode.scala 392:{47,47}]
  wire  _GEN_5202 = 6'h20 == architecturalRegMap_31 | _GEN_5074; // @[decode.scala 392:{47,47}]
  wire  _GEN_5203 = 6'h21 == architecturalRegMap_31 | _GEN_5075; // @[decode.scala 392:{47,47}]
  wire  _GEN_5204 = 6'h22 == architecturalRegMap_31 | _GEN_5076; // @[decode.scala 392:{47,47}]
  wire  _GEN_5205 = 6'h23 == architecturalRegMap_31 | _GEN_5077; // @[decode.scala 392:{47,47}]
  wire  _GEN_5206 = 6'h24 == architecturalRegMap_31 | _GEN_5078; // @[decode.scala 392:{47,47}]
  wire  _GEN_5207 = 6'h25 == architecturalRegMap_31 | _GEN_5079; // @[decode.scala 392:{47,47}]
  wire  _GEN_5208 = 6'h26 == architecturalRegMap_31 | _GEN_5080; // @[decode.scala 392:{47,47}]
  wire  _GEN_5209 = 6'h27 == architecturalRegMap_31 | _GEN_5081; // @[decode.scala 392:{47,47}]
  wire  _GEN_5210 = 6'h28 == architecturalRegMap_31 | _GEN_5082; // @[decode.scala 392:{47,47}]
  wire  _GEN_5211 = 6'h29 == architecturalRegMap_31 | _GEN_5083; // @[decode.scala 392:{47,47}]
  wire  _GEN_5212 = 6'h2a == architecturalRegMap_31 | _GEN_5084; // @[decode.scala 392:{47,47}]
  wire  _GEN_5213 = 6'h2b == architecturalRegMap_31 | _GEN_5085; // @[decode.scala 392:{47,47}]
  wire  _GEN_5214 = 6'h2c == architecturalRegMap_31 | _GEN_5086; // @[decode.scala 392:{47,47}]
  wire  _GEN_5215 = 6'h2d == architecturalRegMap_31 | _GEN_5087; // @[decode.scala 392:{47,47}]
  wire  _GEN_5216 = 6'h2e == architecturalRegMap_31 | _GEN_5088; // @[decode.scala 392:{47,47}]
  wire  _GEN_5217 = 6'h2f == architecturalRegMap_31 | _GEN_5089; // @[decode.scala 392:{47,47}]
  wire  _GEN_5218 = 6'h30 == architecturalRegMap_31 | _GEN_5090; // @[decode.scala 392:{47,47}]
  wire  _GEN_5219 = 6'h31 == architecturalRegMap_31 | _GEN_5091; // @[decode.scala 392:{47,47}]
  wire  _GEN_5220 = 6'h32 == architecturalRegMap_31 | _GEN_5092; // @[decode.scala 392:{47,47}]
  wire  _GEN_5221 = 6'h33 == architecturalRegMap_31 | _GEN_5093; // @[decode.scala 392:{47,47}]
  wire  _GEN_5222 = 6'h34 == architecturalRegMap_31 | _GEN_5094; // @[decode.scala 392:{47,47}]
  wire  _GEN_5223 = 6'h35 == architecturalRegMap_31 | _GEN_5095; // @[decode.scala 392:{47,47}]
  wire  _GEN_5224 = 6'h36 == architecturalRegMap_31 | _GEN_5096; // @[decode.scala 392:{47,47}]
  wire  _GEN_5225 = 6'h37 == architecturalRegMap_31 | _GEN_5097; // @[decode.scala 392:{47,47}]
  wire  _GEN_5226 = 6'h38 == architecturalRegMap_31 | _GEN_5098; // @[decode.scala 392:{47,47}]
  wire  _GEN_5227 = 6'h39 == architecturalRegMap_31 | _GEN_5099; // @[decode.scala 392:{47,47}]
  wire  _GEN_5228 = 6'h3a == architecturalRegMap_31 | _GEN_5100; // @[decode.scala 392:{47,47}]
  wire  _GEN_5229 = 6'h3b == architecturalRegMap_31 | _GEN_5101; // @[decode.scala 392:{47,47}]
  wire  _GEN_5230 = 6'h3c == architecturalRegMap_31 | _GEN_5102; // @[decode.scala 392:{47,47}]
  wire  _GEN_5231 = 6'h3d == architecturalRegMap_31 | _GEN_5103; // @[decode.scala 392:{47,47}]
  wire  _GEN_5232 = 6'h3e == architecturalRegMap_31 | _GEN_5104; // @[decode.scala 392:{47,47}]
  wire  _GEN_5233 = 6'h3f == architecturalRegMap_31 | _GEN_5105; // @[decode.scala 392:{47,47}]
  wire  _GEN_5234 = 6'h0 == architecturalRegMap_31 ? 1'h0 : _GEN_5106; // @[decode.scala 393:{46,46}]
  wire  _GEN_5235 = 6'h1 == architecturalRegMap_31 ? 1'h0 : _GEN_5107; // @[decode.scala 393:{46,46}]
  wire  _GEN_5236 = 6'h2 == architecturalRegMap_31 ? 1'h0 : _GEN_5108; // @[decode.scala 393:{46,46}]
  wire  _GEN_5237 = 6'h3 == architecturalRegMap_31 ? 1'h0 : _GEN_5109; // @[decode.scala 393:{46,46}]
  wire  _GEN_5238 = 6'h4 == architecturalRegMap_31 ? 1'h0 : _GEN_5110; // @[decode.scala 393:{46,46}]
  wire  _GEN_5239 = 6'h5 == architecturalRegMap_31 ? 1'h0 : _GEN_5111; // @[decode.scala 393:{46,46}]
  wire  _GEN_5240 = 6'h6 == architecturalRegMap_31 ? 1'h0 : _GEN_5112; // @[decode.scala 393:{46,46}]
  wire  _GEN_5241 = 6'h7 == architecturalRegMap_31 ? 1'h0 : _GEN_5113; // @[decode.scala 393:{46,46}]
  wire  _GEN_5242 = 6'h8 == architecturalRegMap_31 ? 1'h0 : _GEN_5114; // @[decode.scala 393:{46,46}]
  wire  _GEN_5243 = 6'h9 == architecturalRegMap_31 ? 1'h0 : _GEN_5115; // @[decode.scala 393:{46,46}]
  wire  _GEN_5244 = 6'ha == architecturalRegMap_31 ? 1'h0 : _GEN_5116; // @[decode.scala 393:{46,46}]
  wire  _GEN_5245 = 6'hb == architecturalRegMap_31 ? 1'h0 : _GEN_5117; // @[decode.scala 393:{46,46}]
  wire  _GEN_5246 = 6'hc == architecturalRegMap_31 ? 1'h0 : _GEN_5118; // @[decode.scala 393:{46,46}]
  wire  _GEN_5247 = 6'hd == architecturalRegMap_31 ? 1'h0 : _GEN_5119; // @[decode.scala 393:{46,46}]
  wire  _GEN_5248 = 6'he == architecturalRegMap_31 ? 1'h0 : _GEN_5120; // @[decode.scala 393:{46,46}]
  wire  _GEN_5249 = 6'hf == architecturalRegMap_31 ? 1'h0 : _GEN_5121; // @[decode.scala 393:{46,46}]
  wire  _GEN_5250 = 6'h10 == architecturalRegMap_31 ? 1'h0 : _GEN_5122; // @[decode.scala 393:{46,46}]
  wire  _GEN_5251 = 6'h11 == architecturalRegMap_31 ? 1'h0 : _GEN_5123; // @[decode.scala 393:{46,46}]
  wire  _GEN_5252 = 6'h12 == architecturalRegMap_31 ? 1'h0 : _GEN_5124; // @[decode.scala 393:{46,46}]
  wire  _GEN_5253 = 6'h13 == architecturalRegMap_31 ? 1'h0 : _GEN_5125; // @[decode.scala 393:{46,46}]
  wire  _GEN_5254 = 6'h14 == architecturalRegMap_31 ? 1'h0 : _GEN_5126; // @[decode.scala 393:{46,46}]
  wire  _GEN_5255 = 6'h15 == architecturalRegMap_31 ? 1'h0 : _GEN_5127; // @[decode.scala 393:{46,46}]
  wire  _GEN_5256 = 6'h16 == architecturalRegMap_31 ? 1'h0 : _GEN_5128; // @[decode.scala 393:{46,46}]
  wire  _GEN_5257 = 6'h17 == architecturalRegMap_31 ? 1'h0 : _GEN_5129; // @[decode.scala 393:{46,46}]
  wire  _GEN_5258 = 6'h18 == architecturalRegMap_31 ? 1'h0 : _GEN_5130; // @[decode.scala 393:{46,46}]
  wire  _GEN_5259 = 6'h19 == architecturalRegMap_31 ? 1'h0 : _GEN_5131; // @[decode.scala 393:{46,46}]
  wire  _GEN_5260 = 6'h1a == architecturalRegMap_31 ? 1'h0 : _GEN_5132; // @[decode.scala 393:{46,46}]
  wire  _GEN_5261 = 6'h1b == architecturalRegMap_31 ? 1'h0 : _GEN_5133; // @[decode.scala 393:{46,46}]
  wire  _GEN_5262 = 6'h1c == architecturalRegMap_31 ? 1'h0 : _GEN_5134; // @[decode.scala 393:{46,46}]
  wire  _GEN_5263 = 6'h1d == architecturalRegMap_31 ? 1'h0 : _GEN_5135; // @[decode.scala 393:{46,46}]
  wire  _GEN_5264 = 6'h1e == architecturalRegMap_31 ? 1'h0 : _GEN_5136; // @[decode.scala 393:{46,46}]
  wire  _GEN_5265 = 6'h1f == architecturalRegMap_31 ? 1'h0 : _GEN_5137; // @[decode.scala 393:{46,46}]
  wire  _GEN_5266 = 6'h20 == architecturalRegMap_31 ? 1'h0 : _GEN_5138; // @[decode.scala 393:{46,46}]
  wire  _GEN_5267 = 6'h21 == architecturalRegMap_31 ? 1'h0 : _GEN_5139; // @[decode.scala 393:{46,46}]
  wire  _GEN_5268 = 6'h22 == architecturalRegMap_31 ? 1'h0 : _GEN_5140; // @[decode.scala 393:{46,46}]
  wire  _GEN_5269 = 6'h23 == architecturalRegMap_31 ? 1'h0 : _GEN_5141; // @[decode.scala 393:{46,46}]
  wire  _GEN_5270 = 6'h24 == architecturalRegMap_31 ? 1'h0 : _GEN_5142; // @[decode.scala 393:{46,46}]
  wire  _GEN_5271 = 6'h25 == architecturalRegMap_31 ? 1'h0 : _GEN_5143; // @[decode.scala 393:{46,46}]
  wire  _GEN_5272 = 6'h26 == architecturalRegMap_31 ? 1'h0 : _GEN_5144; // @[decode.scala 393:{46,46}]
  wire  _GEN_5273 = 6'h27 == architecturalRegMap_31 ? 1'h0 : _GEN_5145; // @[decode.scala 393:{46,46}]
  wire  _GEN_5274 = 6'h28 == architecturalRegMap_31 ? 1'h0 : _GEN_5146; // @[decode.scala 393:{46,46}]
  wire  _GEN_5275 = 6'h29 == architecturalRegMap_31 ? 1'h0 : _GEN_5147; // @[decode.scala 393:{46,46}]
  wire  _GEN_5276 = 6'h2a == architecturalRegMap_31 ? 1'h0 : _GEN_5148; // @[decode.scala 393:{46,46}]
  wire  _GEN_5277 = 6'h2b == architecturalRegMap_31 ? 1'h0 : _GEN_5149; // @[decode.scala 393:{46,46}]
  wire  _GEN_5278 = 6'h2c == architecturalRegMap_31 ? 1'h0 : _GEN_5150; // @[decode.scala 393:{46,46}]
  wire  _GEN_5279 = 6'h2d == architecturalRegMap_31 ? 1'h0 : _GEN_5151; // @[decode.scala 393:{46,46}]
  wire  _GEN_5280 = 6'h2e == architecturalRegMap_31 ? 1'h0 : _GEN_5152; // @[decode.scala 393:{46,46}]
  wire  _GEN_5281 = 6'h2f == architecturalRegMap_31 ? 1'h0 : _GEN_5153; // @[decode.scala 393:{46,46}]
  wire  _GEN_5282 = 6'h30 == architecturalRegMap_31 ? 1'h0 : _GEN_5154; // @[decode.scala 393:{46,46}]
  wire  _GEN_5283 = 6'h31 == architecturalRegMap_31 ? 1'h0 : _GEN_5155; // @[decode.scala 393:{46,46}]
  wire  _GEN_5284 = 6'h32 == architecturalRegMap_31 ? 1'h0 : _GEN_5156; // @[decode.scala 393:{46,46}]
  wire  _GEN_5285 = 6'h33 == architecturalRegMap_31 ? 1'h0 : _GEN_5157; // @[decode.scala 393:{46,46}]
  wire  _GEN_5286 = 6'h34 == architecturalRegMap_31 ? 1'h0 : _GEN_5158; // @[decode.scala 393:{46,46}]
  wire  _GEN_5287 = 6'h35 == architecturalRegMap_31 ? 1'h0 : _GEN_5159; // @[decode.scala 393:{46,46}]
  wire  _GEN_5288 = 6'h36 == architecturalRegMap_31 ? 1'h0 : _GEN_5160; // @[decode.scala 393:{46,46}]
  wire  _GEN_5289 = 6'h37 == architecturalRegMap_31 ? 1'h0 : _GEN_5161; // @[decode.scala 393:{46,46}]
  wire  _GEN_5290 = 6'h38 == architecturalRegMap_31 ? 1'h0 : _GEN_5162; // @[decode.scala 393:{46,46}]
  wire  _GEN_5291 = 6'h39 == architecturalRegMap_31 ? 1'h0 : _GEN_5163; // @[decode.scala 393:{46,46}]
  wire  _GEN_5292 = 6'h3a == architecturalRegMap_31 ? 1'h0 : _GEN_5164; // @[decode.scala 393:{46,46}]
  wire  _GEN_5293 = 6'h3b == architecturalRegMap_31 ? 1'h0 : _GEN_5165; // @[decode.scala 393:{46,46}]
  wire  _GEN_5294 = 6'h3c == architecturalRegMap_31 ? 1'h0 : _GEN_5166; // @[decode.scala 393:{46,46}]
  wire  _GEN_5295 = 6'h3d == architecturalRegMap_31 ? 1'h0 : _GEN_5167; // @[decode.scala 393:{46,46}]
  wire  _GEN_5296 = 6'h3e == architecturalRegMap_31 ? 1'h0 : _GEN_5168; // @[decode.scala 393:{46,46}]
  wire  _GEN_5330 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_0 | PRFFreeList_0 : _GEN_5234; // @[decode.scala 381:45 383:22]
  wire  _GEN_5331 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_1 | PRFFreeList_1 : _GEN_5235; // @[decode.scala 381:45 383:22]
  wire  _GEN_5332 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_2 | PRFFreeList_2 : _GEN_5236; // @[decode.scala 381:45 383:22]
  wire  _GEN_5333 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_3 | PRFFreeList_3 : _GEN_5237; // @[decode.scala 381:45 383:22]
  wire  _GEN_5334 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_4 | PRFFreeList_4 : _GEN_5238; // @[decode.scala 381:45 383:22]
  wire  _GEN_5335 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_5 | PRFFreeList_5 : _GEN_5239; // @[decode.scala 381:45 383:22]
  wire  _GEN_5336 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_6 | PRFFreeList_6 : _GEN_5240; // @[decode.scala 381:45 383:22]
  wire  _GEN_5337 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_7 | PRFFreeList_7 : _GEN_5241; // @[decode.scala 381:45 383:22]
  wire  _GEN_5338 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_8 | PRFFreeList_8 : _GEN_5242; // @[decode.scala 381:45 383:22]
  wire  _GEN_5339 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_9 | PRFFreeList_9 : _GEN_5243; // @[decode.scala 381:45 383:22]
  wire  _GEN_5340 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_10 | PRFFreeList_10 : _GEN_5244; // @[decode.scala 381:45 383:22]
  wire  _GEN_5341 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_11 | PRFFreeList_11 : _GEN_5245; // @[decode.scala 381:45 383:22]
  wire  _GEN_5342 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_12 | PRFFreeList_12 : _GEN_5246; // @[decode.scala 381:45 383:22]
  wire  _GEN_5343 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_13 | PRFFreeList_13 : _GEN_5247; // @[decode.scala 381:45 383:22]
  wire  _GEN_5344 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_14 | PRFFreeList_14 : _GEN_5248; // @[decode.scala 381:45 383:22]
  wire  _GEN_5345 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_15 | PRFFreeList_15 : _GEN_5249; // @[decode.scala 381:45 383:22]
  wire  _GEN_5346 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_16 | PRFFreeList_16 : _GEN_5250; // @[decode.scala 381:45 383:22]
  wire  _GEN_5347 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_17 | PRFFreeList_17 : _GEN_5251; // @[decode.scala 381:45 383:22]
  wire  _GEN_5348 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_18 | PRFFreeList_18 : _GEN_5252; // @[decode.scala 381:45 383:22]
  wire  _GEN_5349 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_19 | PRFFreeList_19 : _GEN_5253; // @[decode.scala 381:45 383:22]
  wire  _GEN_5350 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_20 | PRFFreeList_20 : _GEN_5254; // @[decode.scala 381:45 383:22]
  wire  _GEN_5351 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_21 | PRFFreeList_21 : _GEN_5255; // @[decode.scala 381:45 383:22]
  wire  _GEN_5352 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_22 | PRFFreeList_22 : _GEN_5256; // @[decode.scala 381:45 383:22]
  wire  _GEN_5353 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_23 | PRFFreeList_23 : _GEN_5257; // @[decode.scala 381:45 383:22]
  wire  _GEN_5354 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_24 | PRFFreeList_24 : _GEN_5258; // @[decode.scala 381:45 383:22]
  wire  _GEN_5355 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_25 | PRFFreeList_25 : _GEN_5259; // @[decode.scala 381:45 383:22]
  wire  _GEN_5356 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_26 | PRFFreeList_26 : _GEN_5260; // @[decode.scala 381:45 383:22]
  wire  _GEN_5357 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_27 | PRFFreeList_27 : _GEN_5261; // @[decode.scala 381:45 383:22]
  wire  _GEN_5358 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_28 | PRFFreeList_28 : _GEN_5262; // @[decode.scala 381:45 383:22]
  wire  _GEN_5359 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_29 | PRFFreeList_29 : _GEN_5263; // @[decode.scala 381:45 383:22]
  wire  _GEN_5360 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_30 | PRFFreeList_30 : _GEN_5264; // @[decode.scala 381:45 383:22]
  wire  _GEN_5361 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_31 | PRFFreeList_31 : _GEN_5265; // @[decode.scala 381:45 383:22]
  wire  _GEN_5362 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_32 | PRFFreeList_32 : _GEN_5266; // @[decode.scala 381:45 383:22]
  wire  _GEN_5363 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_33 | PRFFreeList_33 : _GEN_5267; // @[decode.scala 381:45 383:22]
  wire  _GEN_5364 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_34 | PRFFreeList_34 : _GEN_5268; // @[decode.scala 381:45 383:22]
  wire  _GEN_5365 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_35 | PRFFreeList_35 : _GEN_5269; // @[decode.scala 381:45 383:22]
  wire  _GEN_5366 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_36 | PRFFreeList_36 : _GEN_5270; // @[decode.scala 381:45 383:22]
  wire  _GEN_5367 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_37 | PRFFreeList_37 : _GEN_5271; // @[decode.scala 381:45 383:22]
  wire  _GEN_5368 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_38 | PRFFreeList_38 : _GEN_5272; // @[decode.scala 381:45 383:22]
  wire  _GEN_5369 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_39 | PRFFreeList_39 : _GEN_5273; // @[decode.scala 381:45 383:22]
  wire  _GEN_5370 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_40 | PRFFreeList_40 : _GEN_5274; // @[decode.scala 381:45 383:22]
  wire  _GEN_5371 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_41 | PRFFreeList_41 : _GEN_5275; // @[decode.scala 381:45 383:22]
  wire  _GEN_5372 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_42 | PRFFreeList_42 : _GEN_5276; // @[decode.scala 381:45 383:22]
  wire  _GEN_5373 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_43 | PRFFreeList_43 : _GEN_5277; // @[decode.scala 381:45 383:22]
  wire  _GEN_5374 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_44 | PRFFreeList_44 : _GEN_5278; // @[decode.scala 381:45 383:22]
  wire  _GEN_5375 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_45 | PRFFreeList_45 : _GEN_5279; // @[decode.scala 381:45 383:22]
  wire  _GEN_5376 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_46 | PRFFreeList_46 : _GEN_5280; // @[decode.scala 381:45 383:22]
  wire  _GEN_5377 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_47 | PRFFreeList_47 : _GEN_5281; // @[decode.scala 381:45 383:22]
  wire  _GEN_5378 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_48 | PRFFreeList_48 : _GEN_5282; // @[decode.scala 381:45 383:22]
  wire  _GEN_5379 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_49 | PRFFreeList_49 : _GEN_5283; // @[decode.scala 381:45 383:22]
  wire  _GEN_5380 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_50 | PRFFreeList_50 : _GEN_5284; // @[decode.scala 381:45 383:22]
  wire  _GEN_5381 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_51 | PRFFreeList_51 : _GEN_5285; // @[decode.scala 381:45 383:22]
  wire  _GEN_5382 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_52 | PRFFreeList_52 : _GEN_5286; // @[decode.scala 381:45 383:22]
  wire  _GEN_5383 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_53 | PRFFreeList_53 : _GEN_5287; // @[decode.scala 381:45 383:22]
  wire  _GEN_5384 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_54 | PRFFreeList_54 : _GEN_5288; // @[decode.scala 381:45 383:22]
  wire  _GEN_5385 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_55 | PRFFreeList_55 : _GEN_5289; // @[decode.scala 381:45 383:22]
  wire  _GEN_5386 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_56 | PRFFreeList_56 : _GEN_5290; // @[decode.scala 381:45 383:22]
  wire  _GEN_5387 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_57 | PRFFreeList_57 : _GEN_5291; // @[decode.scala 381:45 383:22]
  wire  _GEN_5388 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_58 | PRFFreeList_58 : _GEN_5292; // @[decode.scala 381:45 383:22]
  wire  _GEN_5389 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_59 | PRFFreeList_59 : _GEN_5293; // @[decode.scala 381:45 383:22]
  wire  _GEN_5390 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_60 | PRFFreeList_60 : _GEN_5294; // @[decode.scala 381:45 383:22]
  wire  _GEN_5391 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_61 | PRFFreeList_61 : _GEN_5295; // @[decode.scala 381:45 383:22]
  wire  _GEN_5392 = |branchEvalIn_branchMask[3:0] ? reservedFreeList1_62 | PRFFreeList_62 : _GEN_5296; // @[decode.scala 381:45 383:22]
  wire  _GEN_5394 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_0 | PRFValidList_0 : _GEN_5170; // @[decode.scala 381:45 384:22]
  wire  _GEN_5395 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_1 | PRFValidList_1 : _GEN_5171; // @[decode.scala 381:45 384:22]
  wire  _GEN_5396 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_2 | PRFValidList_2 : _GEN_5172; // @[decode.scala 381:45 384:22]
  wire  _GEN_5397 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_3 | PRFValidList_3 : _GEN_5173; // @[decode.scala 381:45 384:22]
  wire  _GEN_5398 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_4 | PRFValidList_4 : _GEN_5174; // @[decode.scala 381:45 384:22]
  wire  _GEN_5399 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_5 | PRFValidList_5 : _GEN_5175; // @[decode.scala 381:45 384:22]
  wire  _GEN_5400 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_6 | PRFValidList_6 : _GEN_5176; // @[decode.scala 381:45 384:22]
  wire  _GEN_5401 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_7 | PRFValidList_7 : _GEN_5177; // @[decode.scala 381:45 384:22]
  wire  _GEN_5402 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_8 | PRFValidList_8 : _GEN_5178; // @[decode.scala 381:45 384:22]
  wire  _GEN_5403 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_9 | PRFValidList_9 : _GEN_5179; // @[decode.scala 381:45 384:22]
  wire  _GEN_5404 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_10 | PRFValidList_10 : _GEN_5180; // @[decode.scala 381:45 384:22]
  wire  _GEN_5405 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_11 | PRFValidList_11 : _GEN_5181; // @[decode.scala 381:45 384:22]
  wire  _GEN_5406 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_12 | PRFValidList_12 : _GEN_5182; // @[decode.scala 381:45 384:22]
  wire  _GEN_5407 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_13 | PRFValidList_13 : _GEN_5183; // @[decode.scala 381:45 384:22]
  wire  _GEN_5408 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_14 | PRFValidList_14 : _GEN_5184; // @[decode.scala 381:45 384:22]
  wire  _GEN_5409 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_15 | PRFValidList_15 : _GEN_5185; // @[decode.scala 381:45 384:22]
  wire  _GEN_5410 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_16 | PRFValidList_16 : _GEN_5186; // @[decode.scala 381:45 384:22]
  wire  _GEN_5411 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_17 | PRFValidList_17 : _GEN_5187; // @[decode.scala 381:45 384:22]
  wire  _GEN_5412 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_18 | PRFValidList_18 : _GEN_5188; // @[decode.scala 381:45 384:22]
  wire  _GEN_5413 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_19 | PRFValidList_19 : _GEN_5189; // @[decode.scala 381:45 384:22]
  wire  _GEN_5414 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_20 | PRFValidList_20 : _GEN_5190; // @[decode.scala 381:45 384:22]
  wire  _GEN_5415 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_21 | PRFValidList_21 : _GEN_5191; // @[decode.scala 381:45 384:22]
  wire  _GEN_5416 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_22 | PRFValidList_22 : _GEN_5192; // @[decode.scala 381:45 384:22]
  wire  _GEN_5417 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_23 | PRFValidList_23 : _GEN_5193; // @[decode.scala 381:45 384:22]
  wire  _GEN_5418 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_24 | PRFValidList_24 : _GEN_5194; // @[decode.scala 381:45 384:22]
  wire  _GEN_5419 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_25 | PRFValidList_25 : _GEN_5195; // @[decode.scala 381:45 384:22]
  wire  _GEN_5420 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_26 | PRFValidList_26 : _GEN_5196; // @[decode.scala 381:45 384:22]
  wire  _GEN_5421 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_27 | PRFValidList_27 : _GEN_5197; // @[decode.scala 381:45 384:22]
  wire  _GEN_5422 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_28 | PRFValidList_28 : _GEN_5198; // @[decode.scala 381:45 384:22]
  wire  _GEN_5423 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_29 | PRFValidList_29 : _GEN_5199; // @[decode.scala 381:45 384:22]
  wire  _GEN_5424 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_30 | PRFValidList_30 : _GEN_5200; // @[decode.scala 381:45 384:22]
  wire  _GEN_5425 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_31 | PRFValidList_31 : _GEN_5201; // @[decode.scala 381:45 384:22]
  wire  _GEN_5426 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_32 | PRFValidList_32 : _GEN_5202; // @[decode.scala 381:45 384:22]
  wire  _GEN_5427 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_33 | PRFValidList_33 : _GEN_5203; // @[decode.scala 381:45 384:22]
  wire  _GEN_5428 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_34 | PRFValidList_34 : _GEN_5204; // @[decode.scala 381:45 384:22]
  wire  _GEN_5429 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_35 | PRFValidList_35 : _GEN_5205; // @[decode.scala 381:45 384:22]
  wire  _GEN_5430 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_36 | PRFValidList_36 : _GEN_5206; // @[decode.scala 381:45 384:22]
  wire  _GEN_5431 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_37 | PRFValidList_37 : _GEN_5207; // @[decode.scala 381:45 384:22]
  wire  _GEN_5432 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_38 | PRFValidList_38 : _GEN_5208; // @[decode.scala 381:45 384:22]
  wire  _GEN_5433 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_39 | PRFValidList_39 : _GEN_5209; // @[decode.scala 381:45 384:22]
  wire  _GEN_5434 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_40 | PRFValidList_40 : _GEN_5210; // @[decode.scala 381:45 384:22]
  wire  _GEN_5435 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_41 | PRFValidList_41 : _GEN_5211; // @[decode.scala 381:45 384:22]
  wire  _GEN_5436 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_42 | PRFValidList_42 : _GEN_5212; // @[decode.scala 381:45 384:22]
  wire  _GEN_5437 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_43 | PRFValidList_43 : _GEN_5213; // @[decode.scala 381:45 384:22]
  wire  _GEN_5438 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_44 | PRFValidList_44 : _GEN_5214; // @[decode.scala 381:45 384:22]
  wire  _GEN_5439 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_45 | PRFValidList_45 : _GEN_5215; // @[decode.scala 381:45 384:22]
  wire  _GEN_5440 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_46 | PRFValidList_46 : _GEN_5216; // @[decode.scala 381:45 384:22]
  wire  _GEN_5441 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_47 | PRFValidList_47 : _GEN_5217; // @[decode.scala 381:45 384:22]
  wire  _GEN_5442 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_48 | PRFValidList_48 : _GEN_5218; // @[decode.scala 381:45 384:22]
  wire  _GEN_5443 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_49 | PRFValidList_49 : _GEN_5219; // @[decode.scala 381:45 384:22]
  wire  _GEN_5444 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_50 | PRFValidList_50 : _GEN_5220; // @[decode.scala 381:45 384:22]
  wire  _GEN_5445 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_51 | PRFValidList_51 : _GEN_5221; // @[decode.scala 381:45 384:22]
  wire  _GEN_5446 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_52 | PRFValidList_52 : _GEN_5222; // @[decode.scala 381:45 384:22]
  wire  _GEN_5447 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_53 | PRFValidList_53 : _GEN_5223; // @[decode.scala 381:45 384:22]
  wire  _GEN_5448 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_54 | PRFValidList_54 : _GEN_5224; // @[decode.scala 381:45 384:22]
  wire  _GEN_5449 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_55 | PRFValidList_55 : _GEN_5225; // @[decode.scala 381:45 384:22]
  wire  _GEN_5450 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_56 | PRFValidList_56 : _GEN_5226; // @[decode.scala 381:45 384:22]
  wire  _GEN_5451 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_57 | PRFValidList_57 : _GEN_5227; // @[decode.scala 381:45 384:22]
  wire  _GEN_5452 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_58 | PRFValidList_58 : _GEN_5228; // @[decode.scala 381:45 384:22]
  wire  _GEN_5453 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_59 | PRFValidList_59 : _GEN_5229; // @[decode.scala 381:45 384:22]
  wire  _GEN_5454 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_60 | PRFValidList_60 : _GEN_5230; // @[decode.scala 381:45 384:22]
  wire  _GEN_5455 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_61 | PRFValidList_61 : _GEN_5231; // @[decode.scala 381:45 384:22]
  wire  _GEN_5456 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_62 | PRFValidList_62 : _GEN_5232; // @[decode.scala 381:45 384:22]
  wire  _GEN_5457 = |branchEvalIn_branchMask[3:0] ? reservedValidList1_63 | PRFValidList_63 : _GEN_5233; // @[decode.scala 381:45 384:22]
  wire  _GEN_5458 = |branchEvalIn_branchMask[3:0] ? coherency : 1'h1; // @[decode.scala 189:26 381:45 389:19]
  wire  _GEN_5460 = _T_434 ? 1'h0 : _T_49[0]; // @[decode.scala 367:29 369:34 372:34]
  wire  _GEN_5461 = _T_434 ? 1'h0 : _T_49[1]; // @[decode.scala 367:29 369:34 373:34]
  wire  _GEN_5462 = _T_434 ? 1'h0 : _T_49[2]; // @[decode.scala 367:29 369:34 374:34]
  wire  _GEN_5463 = _T_434 ? 1'h0 : _T_49[3]; // @[decode.scala 367:29 369:34 375:34]
  wire  _GEN_5464 = _T_434 | _T_49[4]; // @[decode.scala 367:29 369:34 376:34]
  wire [63:0] _GEN_5465 = _T_434 ? branchEvalIn_targetPC : expectedPC; // @[decode.scala 369:34 378:18 188:27]
  wire  _GEN_5498 = _T_434 ? _GEN_5330 : _GEN_1042; // @[decode.scala 369:34]
  wire  _GEN_5499 = _T_434 ? _GEN_5331 : _GEN_1043; // @[decode.scala 369:34]
  wire  _GEN_5500 = _T_434 ? _GEN_5332 : _GEN_1044; // @[decode.scala 369:34]
  wire  _GEN_5501 = _T_434 ? _GEN_5333 : _GEN_1045; // @[decode.scala 369:34]
  wire  _GEN_5502 = _T_434 ? _GEN_5334 : _GEN_1046; // @[decode.scala 369:34]
  wire  _GEN_5503 = _T_434 ? _GEN_5335 : _GEN_1047; // @[decode.scala 369:34]
  wire  _GEN_5504 = _T_434 ? _GEN_5336 : _GEN_1048; // @[decode.scala 369:34]
  wire  _GEN_5505 = _T_434 ? _GEN_5337 : _GEN_1049; // @[decode.scala 369:34]
  wire  _GEN_5506 = _T_434 ? _GEN_5338 : _GEN_1050; // @[decode.scala 369:34]
  wire  _GEN_5507 = _T_434 ? _GEN_5339 : _GEN_1051; // @[decode.scala 369:34]
  wire  _GEN_5508 = _T_434 ? _GEN_5340 : _GEN_1052; // @[decode.scala 369:34]
  wire  _GEN_5509 = _T_434 ? _GEN_5341 : _GEN_1053; // @[decode.scala 369:34]
  wire  _GEN_5510 = _T_434 ? _GEN_5342 : _GEN_1054; // @[decode.scala 369:34]
  wire  _GEN_5511 = _T_434 ? _GEN_5343 : _GEN_1055; // @[decode.scala 369:34]
  wire  _GEN_5512 = _T_434 ? _GEN_5344 : _GEN_1056; // @[decode.scala 369:34]
  wire  _GEN_5513 = _T_434 ? _GEN_5345 : _GEN_1057; // @[decode.scala 369:34]
  wire  _GEN_5514 = _T_434 ? _GEN_5346 : _GEN_1058; // @[decode.scala 369:34]
  wire  _GEN_5515 = _T_434 ? _GEN_5347 : _GEN_1059; // @[decode.scala 369:34]
  wire  _GEN_5516 = _T_434 ? _GEN_5348 : _GEN_1060; // @[decode.scala 369:34]
  wire  _GEN_5517 = _T_434 ? _GEN_5349 : _GEN_1061; // @[decode.scala 369:34]
  wire  _GEN_5518 = _T_434 ? _GEN_5350 : _GEN_1062; // @[decode.scala 369:34]
  wire  _GEN_5519 = _T_434 ? _GEN_5351 : _GEN_1063; // @[decode.scala 369:34]
  wire  _GEN_5520 = _T_434 ? _GEN_5352 : _GEN_1064; // @[decode.scala 369:34]
  wire  _GEN_5521 = _T_434 ? _GEN_5353 : _GEN_1065; // @[decode.scala 369:34]
  wire  _GEN_5522 = _T_434 ? _GEN_5354 : _GEN_1066; // @[decode.scala 369:34]
  wire  _GEN_5523 = _T_434 ? _GEN_5355 : _GEN_1067; // @[decode.scala 369:34]
  wire  _GEN_5524 = _T_434 ? _GEN_5356 : _GEN_1068; // @[decode.scala 369:34]
  wire  _GEN_5525 = _T_434 ? _GEN_5357 : _GEN_1069; // @[decode.scala 369:34]
  wire  _GEN_5526 = _T_434 ? _GEN_5358 : _GEN_1070; // @[decode.scala 369:34]
  wire  _GEN_5527 = _T_434 ? _GEN_5359 : _GEN_1071; // @[decode.scala 369:34]
  wire  _GEN_5528 = _T_434 ? _GEN_5360 : _GEN_1072; // @[decode.scala 369:34]
  wire  _GEN_5529 = _T_434 ? _GEN_5361 : _GEN_1073; // @[decode.scala 369:34]
  wire  _GEN_5530 = _T_434 ? _GEN_5362 : _GEN_1074; // @[decode.scala 369:34]
  wire  _GEN_5531 = _T_434 ? _GEN_5363 : _GEN_1075; // @[decode.scala 369:34]
  wire  _GEN_5532 = _T_434 ? _GEN_5364 : _GEN_1076; // @[decode.scala 369:34]
  wire  _GEN_5533 = _T_434 ? _GEN_5365 : _GEN_1077; // @[decode.scala 369:34]
  wire  _GEN_5534 = _T_434 ? _GEN_5366 : _GEN_1078; // @[decode.scala 369:34]
  wire  _GEN_5535 = _T_434 ? _GEN_5367 : _GEN_1079; // @[decode.scala 369:34]
  wire  _GEN_5536 = _T_434 ? _GEN_5368 : _GEN_1080; // @[decode.scala 369:34]
  wire  _GEN_5537 = _T_434 ? _GEN_5369 : _GEN_1081; // @[decode.scala 369:34]
  wire  _GEN_5538 = _T_434 ? _GEN_5370 : _GEN_1082; // @[decode.scala 369:34]
  wire  _GEN_5539 = _T_434 ? _GEN_5371 : _GEN_1083; // @[decode.scala 369:34]
  wire  _GEN_5540 = _T_434 ? _GEN_5372 : _GEN_1084; // @[decode.scala 369:34]
  wire  _GEN_5541 = _T_434 ? _GEN_5373 : _GEN_1085; // @[decode.scala 369:34]
  wire  _GEN_5542 = _T_434 ? _GEN_5374 : _GEN_1086; // @[decode.scala 369:34]
  wire  _GEN_5543 = _T_434 ? _GEN_5375 : _GEN_1087; // @[decode.scala 369:34]
  wire  _GEN_5544 = _T_434 ? _GEN_5376 : _GEN_1088; // @[decode.scala 369:34]
  wire  _GEN_5545 = _T_434 ? _GEN_5377 : _GEN_1089; // @[decode.scala 369:34]
  wire  _GEN_5546 = _T_434 ? _GEN_5378 : _GEN_1090; // @[decode.scala 369:34]
  wire  _GEN_5547 = _T_434 ? _GEN_5379 : _GEN_1091; // @[decode.scala 369:34]
  wire  _GEN_5548 = _T_434 ? _GEN_5380 : _GEN_1092; // @[decode.scala 369:34]
  wire  _GEN_5549 = _T_434 ? _GEN_5381 : _GEN_1093; // @[decode.scala 369:34]
  wire  _GEN_5550 = _T_434 ? _GEN_5382 : _GEN_1094; // @[decode.scala 369:34]
  wire  _GEN_5551 = _T_434 ? _GEN_5383 : _GEN_1095; // @[decode.scala 369:34]
  wire  _GEN_5552 = _T_434 ? _GEN_5384 : _GEN_1096; // @[decode.scala 369:34]
  wire  _GEN_5553 = _T_434 ? _GEN_5385 : _GEN_1097; // @[decode.scala 369:34]
  wire  _GEN_5554 = _T_434 ? _GEN_5386 : _GEN_1098; // @[decode.scala 369:34]
  wire  _GEN_5555 = _T_434 ? _GEN_5387 : _GEN_1099; // @[decode.scala 369:34]
  wire  _GEN_5556 = _T_434 ? _GEN_5388 : _GEN_1100; // @[decode.scala 369:34]
  wire  _GEN_5557 = _T_434 ? _GEN_5389 : _GEN_1101; // @[decode.scala 369:34]
  wire  _GEN_5558 = _T_434 ? _GEN_5390 : _GEN_1102; // @[decode.scala 369:34]
  wire  _GEN_5559 = _T_434 ? _GEN_5391 : _GEN_1103; // @[decode.scala 369:34]
  wire  _GEN_5560 = _T_434 ? _GEN_5392 : _GEN_1104; // @[decode.scala 369:34]
  wire  _GEN_5562 = _T_434 ? _GEN_5394 : _GEN_1106; // @[decode.scala 369:34]
  wire  _GEN_5563 = _T_434 ? _GEN_5395 : _GEN_1107; // @[decode.scala 369:34]
  wire  _GEN_5564 = _T_434 ? _GEN_5396 : _GEN_1108; // @[decode.scala 369:34]
  wire  _GEN_5565 = _T_434 ? _GEN_5397 : _GEN_1109; // @[decode.scala 369:34]
  wire  _GEN_5566 = _T_434 ? _GEN_5398 : _GEN_1110; // @[decode.scala 369:34]
  wire  _GEN_5567 = _T_434 ? _GEN_5399 : _GEN_1111; // @[decode.scala 369:34]
  wire  _GEN_5568 = _T_434 ? _GEN_5400 : _GEN_1112; // @[decode.scala 369:34]
  wire  _GEN_5569 = _T_434 ? _GEN_5401 : _GEN_1113; // @[decode.scala 369:34]
  wire  _GEN_5570 = _T_434 ? _GEN_5402 : _GEN_1114; // @[decode.scala 369:34]
  wire  _GEN_5571 = _T_434 ? _GEN_5403 : _GEN_1115; // @[decode.scala 369:34]
  wire  _GEN_5572 = _T_434 ? _GEN_5404 : _GEN_1116; // @[decode.scala 369:34]
  wire  _GEN_5573 = _T_434 ? _GEN_5405 : _GEN_1117; // @[decode.scala 369:34]
  wire  _GEN_5574 = _T_434 ? _GEN_5406 : _GEN_1118; // @[decode.scala 369:34]
  wire  _GEN_5575 = _T_434 ? _GEN_5407 : _GEN_1119; // @[decode.scala 369:34]
  wire  _GEN_5576 = _T_434 ? _GEN_5408 : _GEN_1120; // @[decode.scala 369:34]
  wire  _GEN_5577 = _T_434 ? _GEN_5409 : _GEN_1121; // @[decode.scala 369:34]
  wire  _GEN_5578 = _T_434 ? _GEN_5410 : _GEN_1122; // @[decode.scala 369:34]
  wire  _GEN_5579 = _T_434 ? _GEN_5411 : _GEN_1123; // @[decode.scala 369:34]
  wire  _GEN_5580 = _T_434 ? _GEN_5412 : _GEN_1124; // @[decode.scala 369:34]
  wire  _GEN_5581 = _T_434 ? _GEN_5413 : _GEN_1125; // @[decode.scala 369:34]
  wire  _GEN_5582 = _T_434 ? _GEN_5414 : _GEN_1126; // @[decode.scala 369:34]
  wire  _GEN_5583 = _T_434 ? _GEN_5415 : _GEN_1127; // @[decode.scala 369:34]
  wire  _GEN_5584 = _T_434 ? _GEN_5416 : _GEN_1128; // @[decode.scala 369:34]
  wire  _GEN_5585 = _T_434 ? _GEN_5417 : _GEN_1129; // @[decode.scala 369:34]
  wire  _GEN_5586 = _T_434 ? _GEN_5418 : _GEN_1130; // @[decode.scala 369:34]
  wire  _GEN_5587 = _T_434 ? _GEN_5419 : _GEN_1131; // @[decode.scala 369:34]
  wire  _GEN_5588 = _T_434 ? _GEN_5420 : _GEN_1132; // @[decode.scala 369:34]
  wire  _GEN_5589 = _T_434 ? _GEN_5421 : _GEN_1133; // @[decode.scala 369:34]
  wire  _GEN_5590 = _T_434 ? _GEN_5422 : _GEN_1134; // @[decode.scala 369:34]
  wire  _GEN_5591 = _T_434 ? _GEN_5423 : _GEN_1135; // @[decode.scala 369:34]
  wire  _GEN_5592 = _T_434 ? _GEN_5424 : _GEN_1136; // @[decode.scala 369:34]
  wire  _GEN_5593 = _T_434 ? _GEN_5425 : _GEN_1137; // @[decode.scala 369:34]
  wire  _GEN_5594 = _T_434 ? _GEN_5426 : _GEN_1138; // @[decode.scala 369:34]
  wire  _GEN_5595 = _T_434 ? _GEN_5427 : _GEN_1139; // @[decode.scala 369:34]
  wire  _GEN_5596 = _T_434 ? _GEN_5428 : _GEN_1140; // @[decode.scala 369:34]
  wire  _GEN_5597 = _T_434 ? _GEN_5429 : _GEN_1141; // @[decode.scala 369:34]
  wire  _GEN_5598 = _T_434 ? _GEN_5430 : _GEN_1142; // @[decode.scala 369:34]
  wire  _GEN_5599 = _T_434 ? _GEN_5431 : _GEN_1143; // @[decode.scala 369:34]
  wire  _GEN_5600 = _T_434 ? _GEN_5432 : _GEN_1144; // @[decode.scala 369:34]
  wire  _GEN_5601 = _T_434 ? _GEN_5433 : _GEN_1145; // @[decode.scala 369:34]
  wire  _GEN_5602 = _T_434 ? _GEN_5434 : _GEN_1146; // @[decode.scala 369:34]
  wire  _GEN_5603 = _T_434 ? _GEN_5435 : _GEN_1147; // @[decode.scala 369:34]
  wire  _GEN_5604 = _T_434 ? _GEN_5436 : _GEN_1148; // @[decode.scala 369:34]
  wire  _GEN_5605 = _T_434 ? _GEN_5437 : _GEN_1149; // @[decode.scala 369:34]
  wire  _GEN_5606 = _T_434 ? _GEN_5438 : _GEN_1150; // @[decode.scala 369:34]
  wire  _GEN_5607 = _T_434 ? _GEN_5439 : _GEN_1151; // @[decode.scala 369:34]
  wire  _GEN_5608 = _T_434 ? _GEN_5440 : _GEN_1152; // @[decode.scala 369:34]
  wire  _GEN_5609 = _T_434 ? _GEN_5441 : _GEN_1153; // @[decode.scala 369:34]
  wire  _GEN_5610 = _T_434 ? _GEN_5442 : _GEN_1154; // @[decode.scala 369:34]
  wire  _GEN_5611 = _T_434 ? _GEN_5443 : _GEN_1155; // @[decode.scala 369:34]
  wire  _GEN_5612 = _T_434 ? _GEN_5444 : _GEN_1156; // @[decode.scala 369:34]
  wire  _GEN_5613 = _T_434 ? _GEN_5445 : _GEN_1157; // @[decode.scala 369:34]
  wire  _GEN_5614 = _T_434 ? _GEN_5446 : _GEN_1158; // @[decode.scala 369:34]
  wire  _GEN_5615 = _T_434 ? _GEN_5447 : _GEN_1159; // @[decode.scala 369:34]
  wire  _GEN_5616 = _T_434 ? _GEN_5448 : _GEN_1160; // @[decode.scala 369:34]
  wire  _GEN_5617 = _T_434 ? _GEN_5449 : _GEN_1161; // @[decode.scala 369:34]
  wire  _GEN_5618 = _T_434 ? _GEN_5450 : _GEN_1162; // @[decode.scala 369:34]
  wire  _GEN_5619 = _T_434 ? _GEN_5451 : _GEN_1163; // @[decode.scala 369:34]
  wire  _GEN_5620 = _T_434 ? _GEN_5452 : _GEN_1164; // @[decode.scala 369:34]
  wire  _GEN_5621 = _T_434 ? _GEN_5453 : _GEN_1165; // @[decode.scala 369:34]
  wire  _GEN_5622 = _T_434 ? _GEN_5454 : _GEN_1166; // @[decode.scala 369:34]
  wire  _GEN_5623 = _T_434 ? _GEN_5455 : _GEN_1167; // @[decode.scala 369:34]
  wire  _GEN_5624 = _T_434 ? _GEN_5456 : _GEN_1168; // @[decode.scala 369:34]
  wire  _GEN_5625 = _T_434 ? _GEN_5457 : _GEN_1169; // @[decode.scala 369:34]
  wire [2:0] _GEN_5627 = _T_434 ? 3'h0 : _branchTracker_T_1; // @[decode.scala 364:19 369:34 398:21]
  wire [5:0] _GEN_5628 = _T_434 ? reservedRegMap1_0 : reservedRegMap2_0; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5629 = _T_434 ? reservedRegMap1_1 : reservedRegMap2_1; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5630 = _T_434 ? reservedRegMap1_2 : reservedRegMap2_2; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5631 = _T_434 ? reservedRegMap1_3 : reservedRegMap2_3; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5632 = _T_434 ? reservedRegMap1_4 : reservedRegMap2_4; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5633 = _T_434 ? reservedRegMap1_5 : reservedRegMap2_5; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5634 = _T_434 ? reservedRegMap1_6 : reservedRegMap2_6; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5635 = _T_434 ? reservedRegMap1_7 : reservedRegMap2_7; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5636 = _T_434 ? reservedRegMap1_8 : reservedRegMap2_8; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5637 = _T_434 ? reservedRegMap1_9 : reservedRegMap2_9; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5638 = _T_434 ? reservedRegMap1_10 : reservedRegMap2_10; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5639 = _T_434 ? reservedRegMap1_11 : reservedRegMap2_11; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5640 = _T_434 ? reservedRegMap1_12 : reservedRegMap2_12; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5641 = _T_434 ? reservedRegMap1_13 : reservedRegMap2_13; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5642 = _T_434 ? reservedRegMap1_14 : reservedRegMap2_14; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5643 = _T_434 ? reservedRegMap1_15 : reservedRegMap2_15; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5644 = _T_434 ? reservedRegMap1_16 : reservedRegMap2_16; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5645 = _T_434 ? reservedRegMap1_17 : reservedRegMap2_17; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5646 = _T_434 ? reservedRegMap1_18 : reservedRegMap2_18; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5647 = _T_434 ? reservedRegMap1_19 : reservedRegMap2_19; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5648 = _T_434 ? reservedRegMap1_20 : reservedRegMap2_20; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5649 = _T_434 ? reservedRegMap1_21 : reservedRegMap2_21; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5650 = _T_434 ? reservedRegMap1_22 : reservedRegMap2_22; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5651 = _T_434 ? reservedRegMap1_23 : reservedRegMap2_23; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5652 = _T_434 ? reservedRegMap1_24 : reservedRegMap2_24; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5653 = _T_434 ? reservedRegMap1_25 : reservedRegMap2_25; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5654 = _T_434 ? reservedRegMap1_26 : reservedRegMap2_26; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5655 = _T_434 ? reservedRegMap1_27 : reservedRegMap2_27; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5656 = _T_434 ? reservedRegMap1_28 : reservedRegMap2_28; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5657 = _T_434 ? reservedRegMap1_29 : reservedRegMap2_29; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5658 = _T_434 ? reservedRegMap1_30 : reservedRegMap2_30; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5659 = _T_434 ? reservedRegMap1_31 : reservedRegMap2_31; // @[decode.scala 317:28 369:34 400:23]
  wire [5:0] _GEN_5660 = _T_434 ? reservedRegMap2_0 : reservedRegMap3_0; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5661 = _T_434 ? reservedRegMap2_1 : reservedRegMap3_1; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5662 = _T_434 ? reservedRegMap2_2 : reservedRegMap3_2; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5663 = _T_434 ? reservedRegMap2_3 : reservedRegMap3_3; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5664 = _T_434 ? reservedRegMap2_4 : reservedRegMap3_4; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5665 = _T_434 ? reservedRegMap2_5 : reservedRegMap3_5; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5666 = _T_434 ? reservedRegMap2_6 : reservedRegMap3_6; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5667 = _T_434 ? reservedRegMap2_7 : reservedRegMap3_7; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5668 = _T_434 ? reservedRegMap2_8 : reservedRegMap3_8; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5669 = _T_434 ? reservedRegMap2_9 : reservedRegMap3_9; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5670 = _T_434 ? reservedRegMap2_10 : reservedRegMap3_10; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5671 = _T_434 ? reservedRegMap2_11 : reservedRegMap3_11; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5672 = _T_434 ? reservedRegMap2_12 : reservedRegMap3_12; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5673 = _T_434 ? reservedRegMap2_13 : reservedRegMap3_13; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5674 = _T_434 ? reservedRegMap2_14 : reservedRegMap3_14; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5675 = _T_434 ? reservedRegMap2_15 : reservedRegMap3_15; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5676 = _T_434 ? reservedRegMap2_16 : reservedRegMap3_16; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5677 = _T_434 ? reservedRegMap2_17 : reservedRegMap3_17; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5678 = _T_434 ? reservedRegMap2_18 : reservedRegMap3_18; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5679 = _T_434 ? reservedRegMap2_19 : reservedRegMap3_19; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5680 = _T_434 ? reservedRegMap2_20 : reservedRegMap3_20; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5681 = _T_434 ? reservedRegMap2_21 : reservedRegMap3_21; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5682 = _T_434 ? reservedRegMap2_22 : reservedRegMap3_22; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5683 = _T_434 ? reservedRegMap2_23 : reservedRegMap3_23; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5684 = _T_434 ? reservedRegMap2_24 : reservedRegMap3_24; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5685 = _T_434 ? reservedRegMap2_25 : reservedRegMap3_25; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5686 = _T_434 ? reservedRegMap2_26 : reservedRegMap3_26; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5687 = _T_434 ? reservedRegMap2_27 : reservedRegMap3_27; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5688 = _T_434 ? reservedRegMap2_28 : reservedRegMap3_28; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5689 = _T_434 ? reservedRegMap2_29 : reservedRegMap3_29; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5690 = _T_434 ? reservedRegMap2_30 : reservedRegMap3_30; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5691 = _T_434 ? reservedRegMap2_31 : reservedRegMap3_31; // @[decode.scala 318:28 369:34 401:23]
  wire [5:0] _GEN_5692 = _T_434 ? reservedRegMap3_0 : reservedRegMap4_0; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5693 = _T_434 ? reservedRegMap3_1 : reservedRegMap4_1; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5694 = _T_434 ? reservedRegMap3_2 : reservedRegMap4_2; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5695 = _T_434 ? reservedRegMap3_3 : reservedRegMap4_3; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5696 = _T_434 ? reservedRegMap3_4 : reservedRegMap4_4; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5697 = _T_434 ? reservedRegMap3_5 : reservedRegMap4_5; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5698 = _T_434 ? reservedRegMap3_6 : reservedRegMap4_6; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5699 = _T_434 ? reservedRegMap3_7 : reservedRegMap4_7; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5700 = _T_434 ? reservedRegMap3_8 : reservedRegMap4_8; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5701 = _T_434 ? reservedRegMap3_9 : reservedRegMap4_9; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5702 = _T_434 ? reservedRegMap3_10 : reservedRegMap4_10; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5703 = _T_434 ? reservedRegMap3_11 : reservedRegMap4_11; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5704 = _T_434 ? reservedRegMap3_12 : reservedRegMap4_12; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5705 = _T_434 ? reservedRegMap3_13 : reservedRegMap4_13; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5706 = _T_434 ? reservedRegMap3_14 : reservedRegMap4_14; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5707 = _T_434 ? reservedRegMap3_15 : reservedRegMap4_15; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5708 = _T_434 ? reservedRegMap3_16 : reservedRegMap4_16; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5709 = _T_434 ? reservedRegMap3_17 : reservedRegMap4_17; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5710 = _T_434 ? reservedRegMap3_18 : reservedRegMap4_18; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5711 = _T_434 ? reservedRegMap3_19 : reservedRegMap4_19; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5712 = _T_434 ? reservedRegMap3_20 : reservedRegMap4_20; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5713 = _T_434 ? reservedRegMap3_21 : reservedRegMap4_21; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5714 = _T_434 ? reservedRegMap3_22 : reservedRegMap4_22; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5715 = _T_434 ? reservedRegMap3_23 : reservedRegMap4_23; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5716 = _T_434 ? reservedRegMap3_24 : reservedRegMap4_24; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5717 = _T_434 ? reservedRegMap3_25 : reservedRegMap4_25; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5718 = _T_434 ? reservedRegMap3_26 : reservedRegMap4_26; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5719 = _T_434 ? reservedRegMap3_27 : reservedRegMap4_27; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5720 = _T_434 ? reservedRegMap3_28 : reservedRegMap4_28; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5721 = _T_434 ? reservedRegMap3_29 : reservedRegMap4_29; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5722 = _T_434 ? reservedRegMap3_30 : reservedRegMap4_30; // @[decode.scala 319:28 369:34 402:23]
  wire [5:0] _GEN_5723 = _T_434 ? reservedRegMap3_31 : reservedRegMap4_31; // @[decode.scala 319:28 369:34 402:23]
  wire  _GEN_5724 = _T_434 ? reservedFreeList1_0 : reservedFreeList2_0; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5725 = _T_434 ? reservedFreeList1_1 : reservedFreeList2_1; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5726 = _T_434 ? reservedFreeList1_2 : reservedFreeList2_2; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5727 = _T_434 ? reservedFreeList1_3 : reservedFreeList2_3; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5728 = _T_434 ? reservedFreeList1_4 : reservedFreeList2_4; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5729 = _T_434 ? reservedFreeList1_5 : reservedFreeList2_5; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5730 = _T_434 ? reservedFreeList1_6 : reservedFreeList2_6; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5731 = _T_434 ? reservedFreeList1_7 : reservedFreeList2_7; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5732 = _T_434 ? reservedFreeList1_8 : reservedFreeList2_8; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5733 = _T_434 ? reservedFreeList1_9 : reservedFreeList2_9; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5734 = _T_434 ? reservedFreeList1_10 : reservedFreeList2_10; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5735 = _T_434 ? reservedFreeList1_11 : reservedFreeList2_11; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5736 = _T_434 ? reservedFreeList1_12 : reservedFreeList2_12; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5737 = _T_434 ? reservedFreeList1_13 : reservedFreeList2_13; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5738 = _T_434 ? reservedFreeList1_14 : reservedFreeList2_14; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5739 = _T_434 ? reservedFreeList1_15 : reservedFreeList2_15; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5740 = _T_434 ? reservedFreeList1_16 : reservedFreeList2_16; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5741 = _T_434 ? reservedFreeList1_17 : reservedFreeList2_17; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5742 = _T_434 ? reservedFreeList1_18 : reservedFreeList2_18; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5743 = _T_434 ? reservedFreeList1_19 : reservedFreeList2_19; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5744 = _T_434 ? reservedFreeList1_20 : reservedFreeList2_20; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5745 = _T_434 ? reservedFreeList1_21 : reservedFreeList2_21; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5746 = _T_434 ? reservedFreeList1_22 : reservedFreeList2_22; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5747 = _T_434 ? reservedFreeList1_23 : reservedFreeList2_23; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5748 = _T_434 ? reservedFreeList1_24 : reservedFreeList2_24; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5749 = _T_434 ? reservedFreeList1_25 : reservedFreeList2_25; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5750 = _T_434 ? reservedFreeList1_26 : reservedFreeList2_26; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5751 = _T_434 ? reservedFreeList1_27 : reservedFreeList2_27; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5752 = _T_434 ? reservedFreeList1_28 : reservedFreeList2_28; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5753 = _T_434 ? reservedFreeList1_29 : reservedFreeList2_29; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5754 = _T_434 ? reservedFreeList1_30 : reservedFreeList2_30; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5755 = _T_434 ? reservedFreeList1_31 : reservedFreeList2_31; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5756 = _T_434 ? reservedFreeList1_32 : reservedFreeList2_32; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5757 = _T_434 ? reservedFreeList1_33 : reservedFreeList2_33; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5758 = _T_434 ? reservedFreeList1_34 : reservedFreeList2_34; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5759 = _T_434 ? reservedFreeList1_35 : reservedFreeList2_35; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5760 = _T_434 ? reservedFreeList1_36 : reservedFreeList2_36; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5761 = _T_434 ? reservedFreeList1_37 : reservedFreeList2_37; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5762 = _T_434 ? reservedFreeList1_38 : reservedFreeList2_38; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5763 = _T_434 ? reservedFreeList1_39 : reservedFreeList2_39; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5764 = _T_434 ? reservedFreeList1_40 : reservedFreeList2_40; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5765 = _T_434 ? reservedFreeList1_41 : reservedFreeList2_41; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5766 = _T_434 ? reservedFreeList1_42 : reservedFreeList2_42; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5767 = _T_434 ? reservedFreeList1_43 : reservedFreeList2_43; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5768 = _T_434 ? reservedFreeList1_44 : reservedFreeList2_44; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5769 = _T_434 ? reservedFreeList1_45 : reservedFreeList2_45; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5770 = _T_434 ? reservedFreeList1_46 : reservedFreeList2_46; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5771 = _T_434 ? reservedFreeList1_47 : reservedFreeList2_47; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5772 = _T_434 ? reservedFreeList1_48 : reservedFreeList2_48; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5773 = _T_434 ? reservedFreeList1_49 : reservedFreeList2_49; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5774 = _T_434 ? reservedFreeList1_50 : reservedFreeList2_50; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5775 = _T_434 ? reservedFreeList1_51 : reservedFreeList2_51; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5776 = _T_434 ? reservedFreeList1_52 : reservedFreeList2_52; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5777 = _T_434 ? reservedFreeList1_53 : reservedFreeList2_53; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5778 = _T_434 ? reservedFreeList1_54 : reservedFreeList2_54; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5779 = _T_434 ? reservedFreeList1_55 : reservedFreeList2_55; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5780 = _T_434 ? reservedFreeList1_56 : reservedFreeList2_56; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5781 = _T_434 ? reservedFreeList1_57 : reservedFreeList2_57; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5782 = _T_434 ? reservedFreeList1_58 : reservedFreeList2_58; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5783 = _T_434 ? reservedFreeList1_59 : reservedFreeList2_59; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5784 = _T_434 ? reservedFreeList1_60 : reservedFreeList2_60; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5785 = _T_434 ? reservedFreeList1_61 : reservedFreeList2_61; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5786 = _T_434 ? reservedFreeList1_62 : reservedFreeList2_62; // @[decode.scala 322:30 369:34 404:25]
  wire  _GEN_5788 = _T_434 ? reservedFreeList2_0 : reservedFreeList3_0; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5789 = _T_434 ? reservedFreeList2_1 : reservedFreeList3_1; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5790 = _T_434 ? reservedFreeList2_2 : reservedFreeList3_2; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5791 = _T_434 ? reservedFreeList2_3 : reservedFreeList3_3; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5792 = _T_434 ? reservedFreeList2_4 : reservedFreeList3_4; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5793 = _T_434 ? reservedFreeList2_5 : reservedFreeList3_5; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5794 = _T_434 ? reservedFreeList2_6 : reservedFreeList3_6; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5795 = _T_434 ? reservedFreeList2_7 : reservedFreeList3_7; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5796 = _T_434 ? reservedFreeList2_8 : reservedFreeList3_8; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5797 = _T_434 ? reservedFreeList2_9 : reservedFreeList3_9; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5798 = _T_434 ? reservedFreeList2_10 : reservedFreeList3_10; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5799 = _T_434 ? reservedFreeList2_11 : reservedFreeList3_11; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5800 = _T_434 ? reservedFreeList2_12 : reservedFreeList3_12; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5801 = _T_434 ? reservedFreeList2_13 : reservedFreeList3_13; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5802 = _T_434 ? reservedFreeList2_14 : reservedFreeList3_14; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5803 = _T_434 ? reservedFreeList2_15 : reservedFreeList3_15; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5804 = _T_434 ? reservedFreeList2_16 : reservedFreeList3_16; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5805 = _T_434 ? reservedFreeList2_17 : reservedFreeList3_17; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5806 = _T_434 ? reservedFreeList2_18 : reservedFreeList3_18; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5807 = _T_434 ? reservedFreeList2_19 : reservedFreeList3_19; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5808 = _T_434 ? reservedFreeList2_20 : reservedFreeList3_20; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5809 = _T_434 ? reservedFreeList2_21 : reservedFreeList3_21; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5810 = _T_434 ? reservedFreeList2_22 : reservedFreeList3_22; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5811 = _T_434 ? reservedFreeList2_23 : reservedFreeList3_23; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5812 = _T_434 ? reservedFreeList2_24 : reservedFreeList3_24; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5813 = _T_434 ? reservedFreeList2_25 : reservedFreeList3_25; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5814 = _T_434 ? reservedFreeList2_26 : reservedFreeList3_26; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5815 = _T_434 ? reservedFreeList2_27 : reservedFreeList3_27; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5816 = _T_434 ? reservedFreeList2_28 : reservedFreeList3_28; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5817 = _T_434 ? reservedFreeList2_29 : reservedFreeList3_29; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5818 = _T_434 ? reservedFreeList2_30 : reservedFreeList3_30; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5819 = _T_434 ? reservedFreeList2_31 : reservedFreeList3_31; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5820 = _T_434 ? reservedFreeList2_32 : reservedFreeList3_32; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5821 = _T_434 ? reservedFreeList2_33 : reservedFreeList3_33; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5822 = _T_434 ? reservedFreeList2_34 : reservedFreeList3_34; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5823 = _T_434 ? reservedFreeList2_35 : reservedFreeList3_35; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5824 = _T_434 ? reservedFreeList2_36 : reservedFreeList3_36; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5825 = _T_434 ? reservedFreeList2_37 : reservedFreeList3_37; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5826 = _T_434 ? reservedFreeList2_38 : reservedFreeList3_38; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5827 = _T_434 ? reservedFreeList2_39 : reservedFreeList3_39; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5828 = _T_434 ? reservedFreeList2_40 : reservedFreeList3_40; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5829 = _T_434 ? reservedFreeList2_41 : reservedFreeList3_41; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5830 = _T_434 ? reservedFreeList2_42 : reservedFreeList3_42; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5831 = _T_434 ? reservedFreeList2_43 : reservedFreeList3_43; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5832 = _T_434 ? reservedFreeList2_44 : reservedFreeList3_44; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5833 = _T_434 ? reservedFreeList2_45 : reservedFreeList3_45; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5834 = _T_434 ? reservedFreeList2_46 : reservedFreeList3_46; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5835 = _T_434 ? reservedFreeList2_47 : reservedFreeList3_47; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5836 = _T_434 ? reservedFreeList2_48 : reservedFreeList3_48; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5837 = _T_434 ? reservedFreeList2_49 : reservedFreeList3_49; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5838 = _T_434 ? reservedFreeList2_50 : reservedFreeList3_50; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5839 = _T_434 ? reservedFreeList2_51 : reservedFreeList3_51; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5840 = _T_434 ? reservedFreeList2_52 : reservedFreeList3_52; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5841 = _T_434 ? reservedFreeList2_53 : reservedFreeList3_53; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5842 = _T_434 ? reservedFreeList2_54 : reservedFreeList3_54; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5843 = _T_434 ? reservedFreeList2_55 : reservedFreeList3_55; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5844 = _T_434 ? reservedFreeList2_56 : reservedFreeList3_56; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5845 = _T_434 ? reservedFreeList2_57 : reservedFreeList3_57; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5846 = _T_434 ? reservedFreeList2_58 : reservedFreeList3_58; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5847 = _T_434 ? reservedFreeList2_59 : reservedFreeList3_59; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5848 = _T_434 ? reservedFreeList2_60 : reservedFreeList3_60; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5849 = _T_434 ? reservedFreeList2_61 : reservedFreeList3_61; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5850 = _T_434 ? reservedFreeList2_62 : reservedFreeList3_62; // @[decode.scala 323:30 369:34 405:25]
  wire  _GEN_5852 = _T_434 ? reservedFreeList3_0 : reservedFreeList4_0; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5853 = _T_434 ? reservedFreeList3_1 : reservedFreeList4_1; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5854 = _T_434 ? reservedFreeList3_2 : reservedFreeList4_2; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5855 = _T_434 ? reservedFreeList3_3 : reservedFreeList4_3; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5856 = _T_434 ? reservedFreeList3_4 : reservedFreeList4_4; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5857 = _T_434 ? reservedFreeList3_5 : reservedFreeList4_5; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5858 = _T_434 ? reservedFreeList3_6 : reservedFreeList4_6; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5859 = _T_434 ? reservedFreeList3_7 : reservedFreeList4_7; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5860 = _T_434 ? reservedFreeList3_8 : reservedFreeList4_8; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5861 = _T_434 ? reservedFreeList3_9 : reservedFreeList4_9; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5862 = _T_434 ? reservedFreeList3_10 : reservedFreeList4_10; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5863 = _T_434 ? reservedFreeList3_11 : reservedFreeList4_11; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5864 = _T_434 ? reservedFreeList3_12 : reservedFreeList4_12; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5865 = _T_434 ? reservedFreeList3_13 : reservedFreeList4_13; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5866 = _T_434 ? reservedFreeList3_14 : reservedFreeList4_14; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5867 = _T_434 ? reservedFreeList3_15 : reservedFreeList4_15; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5868 = _T_434 ? reservedFreeList3_16 : reservedFreeList4_16; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5869 = _T_434 ? reservedFreeList3_17 : reservedFreeList4_17; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5870 = _T_434 ? reservedFreeList3_18 : reservedFreeList4_18; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5871 = _T_434 ? reservedFreeList3_19 : reservedFreeList4_19; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5872 = _T_434 ? reservedFreeList3_20 : reservedFreeList4_20; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5873 = _T_434 ? reservedFreeList3_21 : reservedFreeList4_21; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5874 = _T_434 ? reservedFreeList3_22 : reservedFreeList4_22; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5875 = _T_434 ? reservedFreeList3_23 : reservedFreeList4_23; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5876 = _T_434 ? reservedFreeList3_24 : reservedFreeList4_24; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5877 = _T_434 ? reservedFreeList3_25 : reservedFreeList4_25; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5878 = _T_434 ? reservedFreeList3_26 : reservedFreeList4_26; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5879 = _T_434 ? reservedFreeList3_27 : reservedFreeList4_27; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5880 = _T_434 ? reservedFreeList3_28 : reservedFreeList4_28; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5881 = _T_434 ? reservedFreeList3_29 : reservedFreeList4_29; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5882 = _T_434 ? reservedFreeList3_30 : reservedFreeList4_30; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5883 = _T_434 ? reservedFreeList3_31 : reservedFreeList4_31; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5884 = _T_434 ? reservedFreeList3_32 : reservedFreeList4_32; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5885 = _T_434 ? reservedFreeList3_33 : reservedFreeList4_33; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5886 = _T_434 ? reservedFreeList3_34 : reservedFreeList4_34; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5887 = _T_434 ? reservedFreeList3_35 : reservedFreeList4_35; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5888 = _T_434 ? reservedFreeList3_36 : reservedFreeList4_36; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5889 = _T_434 ? reservedFreeList3_37 : reservedFreeList4_37; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5890 = _T_434 ? reservedFreeList3_38 : reservedFreeList4_38; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5891 = _T_434 ? reservedFreeList3_39 : reservedFreeList4_39; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5892 = _T_434 ? reservedFreeList3_40 : reservedFreeList4_40; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5893 = _T_434 ? reservedFreeList3_41 : reservedFreeList4_41; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5894 = _T_434 ? reservedFreeList3_42 : reservedFreeList4_42; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5895 = _T_434 ? reservedFreeList3_43 : reservedFreeList4_43; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5896 = _T_434 ? reservedFreeList3_44 : reservedFreeList4_44; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5897 = _T_434 ? reservedFreeList3_45 : reservedFreeList4_45; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5898 = _T_434 ? reservedFreeList3_46 : reservedFreeList4_46; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5899 = _T_434 ? reservedFreeList3_47 : reservedFreeList4_47; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5900 = _T_434 ? reservedFreeList3_48 : reservedFreeList4_48; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5901 = _T_434 ? reservedFreeList3_49 : reservedFreeList4_49; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5902 = _T_434 ? reservedFreeList3_50 : reservedFreeList4_50; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5903 = _T_434 ? reservedFreeList3_51 : reservedFreeList4_51; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5904 = _T_434 ? reservedFreeList3_52 : reservedFreeList4_52; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5905 = _T_434 ? reservedFreeList3_53 : reservedFreeList4_53; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5906 = _T_434 ? reservedFreeList3_54 : reservedFreeList4_54; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5907 = _T_434 ? reservedFreeList3_55 : reservedFreeList4_55; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5908 = _T_434 ? reservedFreeList3_56 : reservedFreeList4_56; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5909 = _T_434 ? reservedFreeList3_57 : reservedFreeList4_57; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5910 = _T_434 ? reservedFreeList3_58 : reservedFreeList4_58; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5911 = _T_434 ? reservedFreeList3_59 : reservedFreeList4_59; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5912 = _T_434 ? reservedFreeList3_60 : reservedFreeList4_60; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5913 = _T_434 ? reservedFreeList3_61 : reservedFreeList4_61; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5914 = _T_434 ? reservedFreeList3_62 : reservedFreeList4_62; // @[decode.scala 324:30 369:34 406:25]
  wire  _GEN_5916 = _T_434 ? reservedValidList1_0 : reservedValidList2_0; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5917 = _T_434 ? reservedValidList1_1 : reservedValidList2_1; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5918 = _T_434 ? reservedValidList1_2 : reservedValidList2_2; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5919 = _T_434 ? reservedValidList1_3 : reservedValidList2_3; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5920 = _T_434 ? reservedValidList1_4 : reservedValidList2_4; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5921 = _T_434 ? reservedValidList1_5 : reservedValidList2_5; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5922 = _T_434 ? reservedValidList1_6 : reservedValidList2_6; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5923 = _T_434 ? reservedValidList1_7 : reservedValidList2_7; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5924 = _T_434 ? reservedValidList1_8 : reservedValidList2_8; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5925 = _T_434 ? reservedValidList1_9 : reservedValidList2_9; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5926 = _T_434 ? reservedValidList1_10 : reservedValidList2_10; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5927 = _T_434 ? reservedValidList1_11 : reservedValidList2_11; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5928 = _T_434 ? reservedValidList1_12 : reservedValidList2_12; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5929 = _T_434 ? reservedValidList1_13 : reservedValidList2_13; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5930 = _T_434 ? reservedValidList1_14 : reservedValidList2_14; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5931 = _T_434 ? reservedValidList1_15 : reservedValidList2_15; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5932 = _T_434 ? reservedValidList1_16 : reservedValidList2_16; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5933 = _T_434 ? reservedValidList1_17 : reservedValidList2_17; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5934 = _T_434 ? reservedValidList1_18 : reservedValidList2_18; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5935 = _T_434 ? reservedValidList1_19 : reservedValidList2_19; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5936 = _T_434 ? reservedValidList1_20 : reservedValidList2_20; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5937 = _T_434 ? reservedValidList1_21 : reservedValidList2_21; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5938 = _T_434 ? reservedValidList1_22 : reservedValidList2_22; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5939 = _T_434 ? reservedValidList1_23 : reservedValidList2_23; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5940 = _T_434 ? reservedValidList1_24 : reservedValidList2_24; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5941 = _T_434 ? reservedValidList1_25 : reservedValidList2_25; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5942 = _T_434 ? reservedValidList1_26 : reservedValidList2_26; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5943 = _T_434 ? reservedValidList1_27 : reservedValidList2_27; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5944 = _T_434 ? reservedValidList1_28 : reservedValidList2_28; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5945 = _T_434 ? reservedValidList1_29 : reservedValidList2_29; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5946 = _T_434 ? reservedValidList1_30 : reservedValidList2_30; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5947 = _T_434 ? reservedValidList1_31 : reservedValidList2_31; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5948 = _T_434 ? reservedValidList1_32 : reservedValidList2_32; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5949 = _T_434 ? reservedValidList1_33 : reservedValidList2_33; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5950 = _T_434 ? reservedValidList1_34 : reservedValidList2_34; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5951 = _T_434 ? reservedValidList1_35 : reservedValidList2_35; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5952 = _T_434 ? reservedValidList1_36 : reservedValidList2_36; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5953 = _T_434 ? reservedValidList1_37 : reservedValidList2_37; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5954 = _T_434 ? reservedValidList1_38 : reservedValidList2_38; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5955 = _T_434 ? reservedValidList1_39 : reservedValidList2_39; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5956 = _T_434 ? reservedValidList1_40 : reservedValidList2_40; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5957 = _T_434 ? reservedValidList1_41 : reservedValidList2_41; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5958 = _T_434 ? reservedValidList1_42 : reservedValidList2_42; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5959 = _T_434 ? reservedValidList1_43 : reservedValidList2_43; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5960 = _T_434 ? reservedValidList1_44 : reservedValidList2_44; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5961 = _T_434 ? reservedValidList1_45 : reservedValidList2_45; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5962 = _T_434 ? reservedValidList1_46 : reservedValidList2_46; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5963 = _T_434 ? reservedValidList1_47 : reservedValidList2_47; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5964 = _T_434 ? reservedValidList1_48 : reservedValidList2_48; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5965 = _T_434 ? reservedValidList1_49 : reservedValidList2_49; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5966 = _T_434 ? reservedValidList1_50 : reservedValidList2_50; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5967 = _T_434 ? reservedValidList1_51 : reservedValidList2_51; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5968 = _T_434 ? reservedValidList1_52 : reservedValidList2_52; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5969 = _T_434 ? reservedValidList1_53 : reservedValidList2_53; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5970 = _T_434 ? reservedValidList1_54 : reservedValidList2_54; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5971 = _T_434 ? reservedValidList1_55 : reservedValidList2_55; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5972 = _T_434 ? reservedValidList1_56 : reservedValidList2_56; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5973 = _T_434 ? reservedValidList1_57 : reservedValidList2_57; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5974 = _T_434 ? reservedValidList1_58 : reservedValidList2_58; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5975 = _T_434 ? reservedValidList1_59 : reservedValidList2_59; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5976 = _T_434 ? reservedValidList1_60 : reservedValidList2_60; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5977 = _T_434 ? reservedValidList1_61 : reservedValidList2_61; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5978 = _T_434 ? reservedValidList1_62 : reservedValidList2_62; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5979 = _T_434 ? reservedValidList1_63 : reservedValidList2_63; // @[decode.scala 327:31 369:34 408:26]
  wire  _GEN_5980 = _T_434 ? reservedValidList2_0 : reservedValidList3_0; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_5981 = _T_434 ? reservedValidList2_1 : reservedValidList3_1; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_5982 = _T_434 ? reservedValidList2_2 : reservedValidList3_2; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_5983 = _T_434 ? reservedValidList2_3 : reservedValidList3_3; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_5984 = _T_434 ? reservedValidList2_4 : reservedValidList3_4; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_5985 = _T_434 ? reservedValidList2_5 : reservedValidList3_5; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_5986 = _T_434 ? reservedValidList2_6 : reservedValidList3_6; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_5987 = _T_434 ? reservedValidList2_7 : reservedValidList3_7; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_5988 = _T_434 ? reservedValidList2_8 : reservedValidList3_8; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_5989 = _T_434 ? reservedValidList2_9 : reservedValidList3_9; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_5990 = _T_434 ? reservedValidList2_10 : reservedValidList3_10; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_5991 = _T_434 ? reservedValidList2_11 : reservedValidList3_11; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_5992 = _T_434 ? reservedValidList2_12 : reservedValidList3_12; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_5993 = _T_434 ? reservedValidList2_13 : reservedValidList3_13; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_5994 = _T_434 ? reservedValidList2_14 : reservedValidList3_14; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_5995 = _T_434 ? reservedValidList2_15 : reservedValidList3_15; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_5996 = _T_434 ? reservedValidList2_16 : reservedValidList3_16; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_5997 = _T_434 ? reservedValidList2_17 : reservedValidList3_17; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_5998 = _T_434 ? reservedValidList2_18 : reservedValidList3_18; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_5999 = _T_434 ? reservedValidList2_19 : reservedValidList3_19; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6000 = _T_434 ? reservedValidList2_20 : reservedValidList3_20; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6001 = _T_434 ? reservedValidList2_21 : reservedValidList3_21; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6002 = _T_434 ? reservedValidList2_22 : reservedValidList3_22; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6003 = _T_434 ? reservedValidList2_23 : reservedValidList3_23; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6004 = _T_434 ? reservedValidList2_24 : reservedValidList3_24; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6005 = _T_434 ? reservedValidList2_25 : reservedValidList3_25; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6006 = _T_434 ? reservedValidList2_26 : reservedValidList3_26; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6007 = _T_434 ? reservedValidList2_27 : reservedValidList3_27; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6008 = _T_434 ? reservedValidList2_28 : reservedValidList3_28; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6009 = _T_434 ? reservedValidList2_29 : reservedValidList3_29; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6010 = _T_434 ? reservedValidList2_30 : reservedValidList3_30; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6011 = _T_434 ? reservedValidList2_31 : reservedValidList3_31; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6012 = _T_434 ? reservedValidList2_32 : reservedValidList3_32; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6013 = _T_434 ? reservedValidList2_33 : reservedValidList3_33; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6014 = _T_434 ? reservedValidList2_34 : reservedValidList3_34; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6015 = _T_434 ? reservedValidList2_35 : reservedValidList3_35; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6016 = _T_434 ? reservedValidList2_36 : reservedValidList3_36; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6017 = _T_434 ? reservedValidList2_37 : reservedValidList3_37; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6018 = _T_434 ? reservedValidList2_38 : reservedValidList3_38; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6019 = _T_434 ? reservedValidList2_39 : reservedValidList3_39; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6020 = _T_434 ? reservedValidList2_40 : reservedValidList3_40; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6021 = _T_434 ? reservedValidList2_41 : reservedValidList3_41; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6022 = _T_434 ? reservedValidList2_42 : reservedValidList3_42; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6023 = _T_434 ? reservedValidList2_43 : reservedValidList3_43; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6024 = _T_434 ? reservedValidList2_44 : reservedValidList3_44; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6025 = _T_434 ? reservedValidList2_45 : reservedValidList3_45; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6026 = _T_434 ? reservedValidList2_46 : reservedValidList3_46; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6027 = _T_434 ? reservedValidList2_47 : reservedValidList3_47; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6028 = _T_434 ? reservedValidList2_48 : reservedValidList3_48; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6029 = _T_434 ? reservedValidList2_49 : reservedValidList3_49; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6030 = _T_434 ? reservedValidList2_50 : reservedValidList3_50; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6031 = _T_434 ? reservedValidList2_51 : reservedValidList3_51; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6032 = _T_434 ? reservedValidList2_52 : reservedValidList3_52; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6033 = _T_434 ? reservedValidList2_53 : reservedValidList3_53; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6034 = _T_434 ? reservedValidList2_54 : reservedValidList3_54; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6035 = _T_434 ? reservedValidList2_55 : reservedValidList3_55; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6036 = _T_434 ? reservedValidList2_56 : reservedValidList3_56; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6037 = _T_434 ? reservedValidList2_57 : reservedValidList3_57; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6038 = _T_434 ? reservedValidList2_58 : reservedValidList3_58; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6039 = _T_434 ? reservedValidList2_59 : reservedValidList3_59; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6040 = _T_434 ? reservedValidList2_60 : reservedValidList3_60; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6041 = _T_434 ? reservedValidList2_61 : reservedValidList3_61; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6042 = _T_434 ? reservedValidList2_62 : reservedValidList3_62; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6043 = _T_434 ? reservedValidList2_63 : reservedValidList3_63; // @[decode.scala 328:31 369:34 409:26]
  wire  _GEN_6044 = _T_434 ? reservedValidList3_0 : reservedValidList4_0; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6045 = _T_434 ? reservedValidList3_1 : reservedValidList4_1; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6046 = _T_434 ? reservedValidList3_2 : reservedValidList4_2; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6047 = _T_434 ? reservedValidList3_3 : reservedValidList4_3; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6048 = _T_434 ? reservedValidList3_4 : reservedValidList4_4; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6049 = _T_434 ? reservedValidList3_5 : reservedValidList4_5; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6050 = _T_434 ? reservedValidList3_6 : reservedValidList4_6; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6051 = _T_434 ? reservedValidList3_7 : reservedValidList4_7; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6052 = _T_434 ? reservedValidList3_8 : reservedValidList4_8; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6053 = _T_434 ? reservedValidList3_9 : reservedValidList4_9; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6054 = _T_434 ? reservedValidList3_10 : reservedValidList4_10; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6055 = _T_434 ? reservedValidList3_11 : reservedValidList4_11; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6056 = _T_434 ? reservedValidList3_12 : reservedValidList4_12; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6057 = _T_434 ? reservedValidList3_13 : reservedValidList4_13; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6058 = _T_434 ? reservedValidList3_14 : reservedValidList4_14; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6059 = _T_434 ? reservedValidList3_15 : reservedValidList4_15; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6060 = _T_434 ? reservedValidList3_16 : reservedValidList4_16; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6061 = _T_434 ? reservedValidList3_17 : reservedValidList4_17; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6062 = _T_434 ? reservedValidList3_18 : reservedValidList4_18; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6063 = _T_434 ? reservedValidList3_19 : reservedValidList4_19; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6064 = _T_434 ? reservedValidList3_20 : reservedValidList4_20; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6065 = _T_434 ? reservedValidList3_21 : reservedValidList4_21; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6066 = _T_434 ? reservedValidList3_22 : reservedValidList4_22; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6067 = _T_434 ? reservedValidList3_23 : reservedValidList4_23; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6068 = _T_434 ? reservedValidList3_24 : reservedValidList4_24; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6069 = _T_434 ? reservedValidList3_25 : reservedValidList4_25; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6070 = _T_434 ? reservedValidList3_26 : reservedValidList4_26; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6071 = _T_434 ? reservedValidList3_27 : reservedValidList4_27; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6072 = _T_434 ? reservedValidList3_28 : reservedValidList4_28; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6073 = _T_434 ? reservedValidList3_29 : reservedValidList4_29; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6074 = _T_434 ? reservedValidList3_30 : reservedValidList4_30; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6075 = _T_434 ? reservedValidList3_31 : reservedValidList4_31; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6076 = _T_434 ? reservedValidList3_32 : reservedValidList4_32; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6077 = _T_434 ? reservedValidList3_33 : reservedValidList4_33; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6078 = _T_434 ? reservedValidList3_34 : reservedValidList4_34; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6079 = _T_434 ? reservedValidList3_35 : reservedValidList4_35; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6080 = _T_434 ? reservedValidList3_36 : reservedValidList4_36; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6081 = _T_434 ? reservedValidList3_37 : reservedValidList4_37; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6082 = _T_434 ? reservedValidList3_38 : reservedValidList4_38; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6083 = _T_434 ? reservedValidList3_39 : reservedValidList4_39; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6084 = _T_434 ? reservedValidList3_40 : reservedValidList4_40; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6085 = _T_434 ? reservedValidList3_41 : reservedValidList4_41; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6086 = _T_434 ? reservedValidList3_42 : reservedValidList4_42; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6087 = _T_434 ? reservedValidList3_43 : reservedValidList4_43; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6088 = _T_434 ? reservedValidList3_44 : reservedValidList4_44; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6089 = _T_434 ? reservedValidList3_45 : reservedValidList4_45; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6090 = _T_434 ? reservedValidList3_46 : reservedValidList4_46; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6091 = _T_434 ? reservedValidList3_47 : reservedValidList4_47; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6092 = _T_434 ? reservedValidList3_48 : reservedValidList4_48; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6093 = _T_434 ? reservedValidList3_49 : reservedValidList4_49; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6094 = _T_434 ? reservedValidList3_50 : reservedValidList4_50; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6095 = _T_434 ? reservedValidList3_51 : reservedValidList4_51; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6096 = _T_434 ? reservedValidList3_52 : reservedValidList4_52; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6097 = _T_434 ? reservedValidList3_53 : reservedValidList4_53; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6098 = _T_434 ? reservedValidList3_54 : reservedValidList4_54; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6099 = _T_434 ? reservedValidList3_55 : reservedValidList4_55; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6100 = _T_434 ? reservedValidList3_56 : reservedValidList4_56; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6101 = _T_434 ? reservedValidList3_57 : reservedValidList4_57; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6102 = _T_434 ? reservedValidList3_58 : reservedValidList4_58; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6103 = _T_434 ? reservedValidList3_59 : reservedValidList4_59; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6104 = _T_434 ? reservedValidList3_60 : reservedValidList4_60; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6105 = _T_434 ? reservedValidList3_61 : reservedValidList4_61; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6106 = _T_434 ? reservedValidList3_62 : reservedValidList4_62; // @[decode.scala 329:31 369:34 410:26]
  wire  _GEN_6107 = _T_434 ? reservedValidList3_63 : reservedValidList4_63; // @[decode.scala 329:31 369:34 410:26]
  wire [2:0] _GEN_6108 = branchEvalIn_fired ? _GEN_5627 : branchTracker; // @[decode.scala 363:28 178:30]
  wire  _GEN_6109 = branchEvalIn_fired ? _GEN_5460 : branchBuffer_branchMask_0; // @[decode.scala 363:28 142:29]
  wire  _GEN_6110 = branchEvalIn_fired ? _GEN_5461 : branchBuffer_branchMask_1; // @[decode.scala 363:28 142:29]
  wire  _GEN_6111 = branchEvalIn_fired ? _GEN_5462 : branchBuffer_branchMask_2; // @[decode.scala 363:28 142:29]
  wire  _GEN_6112 = branchEvalIn_fired ? _GEN_5463 : branchBuffer_branchMask_3; // @[decode.scala 363:28 142:29]
  wire  _GEN_6113 = branchEvalIn_fired ? _GEN_5464 : branchBuffer_branchMask_4; // @[decode.scala 363:28 142:29]
  wire [63:0] _GEN_6115 = branchEvalIn_fired ? _GEN_5465 : expectedPC; // @[decode.scala 188:27 363:28]
  wire  _GEN_6148 = branchEvalIn_fired ? _GEN_5498 : _GEN_1042; // @[decode.scala 363:28]
  wire  _GEN_6149 = branchEvalIn_fired ? _GEN_5499 : _GEN_1043; // @[decode.scala 363:28]
  wire  _GEN_6150 = branchEvalIn_fired ? _GEN_5500 : _GEN_1044; // @[decode.scala 363:28]
  wire  _GEN_6151 = branchEvalIn_fired ? _GEN_5501 : _GEN_1045; // @[decode.scala 363:28]
  wire  _GEN_6152 = branchEvalIn_fired ? _GEN_5502 : _GEN_1046; // @[decode.scala 363:28]
  wire  _GEN_6153 = branchEvalIn_fired ? _GEN_5503 : _GEN_1047; // @[decode.scala 363:28]
  wire  _GEN_6154 = branchEvalIn_fired ? _GEN_5504 : _GEN_1048; // @[decode.scala 363:28]
  wire  _GEN_6155 = branchEvalIn_fired ? _GEN_5505 : _GEN_1049; // @[decode.scala 363:28]
  wire  _GEN_6156 = branchEvalIn_fired ? _GEN_5506 : _GEN_1050; // @[decode.scala 363:28]
  wire  _GEN_6157 = branchEvalIn_fired ? _GEN_5507 : _GEN_1051; // @[decode.scala 363:28]
  wire  _GEN_6158 = branchEvalIn_fired ? _GEN_5508 : _GEN_1052; // @[decode.scala 363:28]
  wire  _GEN_6159 = branchEvalIn_fired ? _GEN_5509 : _GEN_1053; // @[decode.scala 363:28]
  wire  _GEN_6160 = branchEvalIn_fired ? _GEN_5510 : _GEN_1054; // @[decode.scala 363:28]
  wire  _GEN_6161 = branchEvalIn_fired ? _GEN_5511 : _GEN_1055; // @[decode.scala 363:28]
  wire  _GEN_6162 = branchEvalIn_fired ? _GEN_5512 : _GEN_1056; // @[decode.scala 363:28]
  wire  _GEN_6163 = branchEvalIn_fired ? _GEN_5513 : _GEN_1057; // @[decode.scala 363:28]
  wire  _GEN_6164 = branchEvalIn_fired ? _GEN_5514 : _GEN_1058; // @[decode.scala 363:28]
  wire  _GEN_6165 = branchEvalIn_fired ? _GEN_5515 : _GEN_1059; // @[decode.scala 363:28]
  wire  _GEN_6166 = branchEvalIn_fired ? _GEN_5516 : _GEN_1060; // @[decode.scala 363:28]
  wire  _GEN_6167 = branchEvalIn_fired ? _GEN_5517 : _GEN_1061; // @[decode.scala 363:28]
  wire  _GEN_6168 = branchEvalIn_fired ? _GEN_5518 : _GEN_1062; // @[decode.scala 363:28]
  wire  _GEN_6169 = branchEvalIn_fired ? _GEN_5519 : _GEN_1063; // @[decode.scala 363:28]
  wire  _GEN_6170 = branchEvalIn_fired ? _GEN_5520 : _GEN_1064; // @[decode.scala 363:28]
  wire  _GEN_6171 = branchEvalIn_fired ? _GEN_5521 : _GEN_1065; // @[decode.scala 363:28]
  wire  _GEN_6172 = branchEvalIn_fired ? _GEN_5522 : _GEN_1066; // @[decode.scala 363:28]
  wire  _GEN_6173 = branchEvalIn_fired ? _GEN_5523 : _GEN_1067; // @[decode.scala 363:28]
  wire  _GEN_6174 = branchEvalIn_fired ? _GEN_5524 : _GEN_1068; // @[decode.scala 363:28]
  wire  _GEN_6175 = branchEvalIn_fired ? _GEN_5525 : _GEN_1069; // @[decode.scala 363:28]
  wire  _GEN_6176 = branchEvalIn_fired ? _GEN_5526 : _GEN_1070; // @[decode.scala 363:28]
  wire  _GEN_6177 = branchEvalIn_fired ? _GEN_5527 : _GEN_1071; // @[decode.scala 363:28]
  wire  _GEN_6178 = branchEvalIn_fired ? _GEN_5528 : _GEN_1072; // @[decode.scala 363:28]
  wire  _GEN_6179 = branchEvalIn_fired ? _GEN_5529 : _GEN_1073; // @[decode.scala 363:28]
  wire  _GEN_6180 = branchEvalIn_fired ? _GEN_5530 : _GEN_1074; // @[decode.scala 363:28]
  wire  _GEN_6181 = branchEvalIn_fired ? _GEN_5531 : _GEN_1075; // @[decode.scala 363:28]
  wire  _GEN_6182 = branchEvalIn_fired ? _GEN_5532 : _GEN_1076; // @[decode.scala 363:28]
  wire  _GEN_6183 = branchEvalIn_fired ? _GEN_5533 : _GEN_1077; // @[decode.scala 363:28]
  wire  _GEN_6184 = branchEvalIn_fired ? _GEN_5534 : _GEN_1078; // @[decode.scala 363:28]
  wire  _GEN_6185 = branchEvalIn_fired ? _GEN_5535 : _GEN_1079; // @[decode.scala 363:28]
  wire  _GEN_6186 = branchEvalIn_fired ? _GEN_5536 : _GEN_1080; // @[decode.scala 363:28]
  wire  _GEN_6187 = branchEvalIn_fired ? _GEN_5537 : _GEN_1081; // @[decode.scala 363:28]
  wire  _GEN_6188 = branchEvalIn_fired ? _GEN_5538 : _GEN_1082; // @[decode.scala 363:28]
  wire  _GEN_6189 = branchEvalIn_fired ? _GEN_5539 : _GEN_1083; // @[decode.scala 363:28]
  wire  _GEN_6190 = branchEvalIn_fired ? _GEN_5540 : _GEN_1084; // @[decode.scala 363:28]
  wire  _GEN_6191 = branchEvalIn_fired ? _GEN_5541 : _GEN_1085; // @[decode.scala 363:28]
  wire  _GEN_6192 = branchEvalIn_fired ? _GEN_5542 : _GEN_1086; // @[decode.scala 363:28]
  wire  _GEN_6193 = branchEvalIn_fired ? _GEN_5543 : _GEN_1087; // @[decode.scala 363:28]
  wire  _GEN_6194 = branchEvalIn_fired ? _GEN_5544 : _GEN_1088; // @[decode.scala 363:28]
  wire  _GEN_6195 = branchEvalIn_fired ? _GEN_5545 : _GEN_1089; // @[decode.scala 363:28]
  wire  _GEN_6196 = branchEvalIn_fired ? _GEN_5546 : _GEN_1090; // @[decode.scala 363:28]
  wire  _GEN_6197 = branchEvalIn_fired ? _GEN_5547 : _GEN_1091; // @[decode.scala 363:28]
  wire  _GEN_6198 = branchEvalIn_fired ? _GEN_5548 : _GEN_1092; // @[decode.scala 363:28]
  wire  _GEN_6199 = branchEvalIn_fired ? _GEN_5549 : _GEN_1093; // @[decode.scala 363:28]
  wire  _GEN_6200 = branchEvalIn_fired ? _GEN_5550 : _GEN_1094; // @[decode.scala 363:28]
  wire  _GEN_6201 = branchEvalIn_fired ? _GEN_5551 : _GEN_1095; // @[decode.scala 363:28]
  wire  _GEN_6202 = branchEvalIn_fired ? _GEN_5552 : _GEN_1096; // @[decode.scala 363:28]
  wire  _GEN_6203 = branchEvalIn_fired ? _GEN_5553 : _GEN_1097; // @[decode.scala 363:28]
  wire  _GEN_6204 = branchEvalIn_fired ? _GEN_5554 : _GEN_1098; // @[decode.scala 363:28]
  wire  _GEN_6205 = branchEvalIn_fired ? _GEN_5555 : _GEN_1099; // @[decode.scala 363:28]
  wire  _GEN_6206 = branchEvalIn_fired ? _GEN_5556 : _GEN_1100; // @[decode.scala 363:28]
  wire  _GEN_6207 = branchEvalIn_fired ? _GEN_5557 : _GEN_1101; // @[decode.scala 363:28]
  wire  _GEN_6208 = branchEvalIn_fired ? _GEN_5558 : _GEN_1102; // @[decode.scala 363:28]
  wire  _GEN_6209 = branchEvalIn_fired ? _GEN_5559 : _GEN_1103; // @[decode.scala 363:28]
  wire  _GEN_6210 = branchEvalIn_fired ? _GEN_5560 : _GEN_1104; // @[decode.scala 363:28]
  wire  _GEN_6212 = branchEvalIn_fired ? _GEN_5562 : _GEN_1106; // @[decode.scala 363:28]
  wire  _GEN_6213 = branchEvalIn_fired ? _GEN_5563 : _GEN_1107; // @[decode.scala 363:28]
  wire  _GEN_6214 = branchEvalIn_fired ? _GEN_5564 : _GEN_1108; // @[decode.scala 363:28]
  wire  _GEN_6215 = branchEvalIn_fired ? _GEN_5565 : _GEN_1109; // @[decode.scala 363:28]
  wire  _GEN_6216 = branchEvalIn_fired ? _GEN_5566 : _GEN_1110; // @[decode.scala 363:28]
  wire  _GEN_6217 = branchEvalIn_fired ? _GEN_5567 : _GEN_1111; // @[decode.scala 363:28]
  wire  _GEN_6218 = branchEvalIn_fired ? _GEN_5568 : _GEN_1112; // @[decode.scala 363:28]
  wire  _GEN_6219 = branchEvalIn_fired ? _GEN_5569 : _GEN_1113; // @[decode.scala 363:28]
  wire  _GEN_6220 = branchEvalIn_fired ? _GEN_5570 : _GEN_1114; // @[decode.scala 363:28]
  wire  _GEN_6221 = branchEvalIn_fired ? _GEN_5571 : _GEN_1115; // @[decode.scala 363:28]
  wire  _GEN_6222 = branchEvalIn_fired ? _GEN_5572 : _GEN_1116; // @[decode.scala 363:28]
  wire  _GEN_6223 = branchEvalIn_fired ? _GEN_5573 : _GEN_1117; // @[decode.scala 363:28]
  wire  _GEN_6224 = branchEvalIn_fired ? _GEN_5574 : _GEN_1118; // @[decode.scala 363:28]
  wire  _GEN_6225 = branchEvalIn_fired ? _GEN_5575 : _GEN_1119; // @[decode.scala 363:28]
  wire  _GEN_6226 = branchEvalIn_fired ? _GEN_5576 : _GEN_1120; // @[decode.scala 363:28]
  wire  _GEN_6227 = branchEvalIn_fired ? _GEN_5577 : _GEN_1121; // @[decode.scala 363:28]
  wire  _GEN_6228 = branchEvalIn_fired ? _GEN_5578 : _GEN_1122; // @[decode.scala 363:28]
  wire  _GEN_6229 = branchEvalIn_fired ? _GEN_5579 : _GEN_1123; // @[decode.scala 363:28]
  wire  _GEN_6230 = branchEvalIn_fired ? _GEN_5580 : _GEN_1124; // @[decode.scala 363:28]
  wire  _GEN_6231 = branchEvalIn_fired ? _GEN_5581 : _GEN_1125; // @[decode.scala 363:28]
  wire  _GEN_6232 = branchEvalIn_fired ? _GEN_5582 : _GEN_1126; // @[decode.scala 363:28]
  wire  _GEN_6233 = branchEvalIn_fired ? _GEN_5583 : _GEN_1127; // @[decode.scala 363:28]
  wire  _GEN_6234 = branchEvalIn_fired ? _GEN_5584 : _GEN_1128; // @[decode.scala 363:28]
  wire  _GEN_6235 = branchEvalIn_fired ? _GEN_5585 : _GEN_1129; // @[decode.scala 363:28]
  wire  _GEN_6236 = branchEvalIn_fired ? _GEN_5586 : _GEN_1130; // @[decode.scala 363:28]
  wire  _GEN_6237 = branchEvalIn_fired ? _GEN_5587 : _GEN_1131; // @[decode.scala 363:28]
  wire  _GEN_6238 = branchEvalIn_fired ? _GEN_5588 : _GEN_1132; // @[decode.scala 363:28]
  wire  _GEN_6239 = branchEvalIn_fired ? _GEN_5589 : _GEN_1133; // @[decode.scala 363:28]
  wire  _GEN_6240 = branchEvalIn_fired ? _GEN_5590 : _GEN_1134; // @[decode.scala 363:28]
  wire  _GEN_6241 = branchEvalIn_fired ? _GEN_5591 : _GEN_1135; // @[decode.scala 363:28]
  wire  _GEN_6242 = branchEvalIn_fired ? _GEN_5592 : _GEN_1136; // @[decode.scala 363:28]
  wire  _GEN_6243 = branchEvalIn_fired ? _GEN_5593 : _GEN_1137; // @[decode.scala 363:28]
  wire  _GEN_6244 = branchEvalIn_fired ? _GEN_5594 : _GEN_1138; // @[decode.scala 363:28]
  wire  _GEN_6245 = branchEvalIn_fired ? _GEN_5595 : _GEN_1139; // @[decode.scala 363:28]
  wire  _GEN_6246 = branchEvalIn_fired ? _GEN_5596 : _GEN_1140; // @[decode.scala 363:28]
  wire  _GEN_6247 = branchEvalIn_fired ? _GEN_5597 : _GEN_1141; // @[decode.scala 363:28]
  wire  _GEN_6248 = branchEvalIn_fired ? _GEN_5598 : _GEN_1142; // @[decode.scala 363:28]
  wire  _GEN_6249 = branchEvalIn_fired ? _GEN_5599 : _GEN_1143; // @[decode.scala 363:28]
  wire  _GEN_6250 = branchEvalIn_fired ? _GEN_5600 : _GEN_1144; // @[decode.scala 363:28]
  wire  _GEN_6251 = branchEvalIn_fired ? _GEN_5601 : _GEN_1145; // @[decode.scala 363:28]
  wire  _GEN_6252 = branchEvalIn_fired ? _GEN_5602 : _GEN_1146; // @[decode.scala 363:28]
  wire  _GEN_6253 = branchEvalIn_fired ? _GEN_5603 : _GEN_1147; // @[decode.scala 363:28]
  wire  _GEN_6254 = branchEvalIn_fired ? _GEN_5604 : _GEN_1148; // @[decode.scala 363:28]
  wire  _GEN_6255 = branchEvalIn_fired ? _GEN_5605 : _GEN_1149; // @[decode.scala 363:28]
  wire  _GEN_6256 = branchEvalIn_fired ? _GEN_5606 : _GEN_1150; // @[decode.scala 363:28]
  wire  _GEN_6257 = branchEvalIn_fired ? _GEN_5607 : _GEN_1151; // @[decode.scala 363:28]
  wire  _GEN_6258 = branchEvalIn_fired ? _GEN_5608 : _GEN_1152; // @[decode.scala 363:28]
  wire  _GEN_6259 = branchEvalIn_fired ? _GEN_5609 : _GEN_1153; // @[decode.scala 363:28]
  wire  _GEN_6260 = branchEvalIn_fired ? _GEN_5610 : _GEN_1154; // @[decode.scala 363:28]
  wire  _GEN_6261 = branchEvalIn_fired ? _GEN_5611 : _GEN_1155; // @[decode.scala 363:28]
  wire  _GEN_6262 = branchEvalIn_fired ? _GEN_5612 : _GEN_1156; // @[decode.scala 363:28]
  wire  _GEN_6263 = branchEvalIn_fired ? _GEN_5613 : _GEN_1157; // @[decode.scala 363:28]
  wire  _GEN_6264 = branchEvalIn_fired ? _GEN_5614 : _GEN_1158; // @[decode.scala 363:28]
  wire  _GEN_6265 = branchEvalIn_fired ? _GEN_5615 : _GEN_1159; // @[decode.scala 363:28]
  wire  _GEN_6266 = branchEvalIn_fired ? _GEN_5616 : _GEN_1160; // @[decode.scala 363:28]
  wire  _GEN_6267 = branchEvalIn_fired ? _GEN_5617 : _GEN_1161; // @[decode.scala 363:28]
  wire  _GEN_6268 = branchEvalIn_fired ? _GEN_5618 : _GEN_1162; // @[decode.scala 363:28]
  wire  _GEN_6269 = branchEvalIn_fired ? _GEN_5619 : _GEN_1163; // @[decode.scala 363:28]
  wire  _GEN_6270 = branchEvalIn_fired ? _GEN_5620 : _GEN_1164; // @[decode.scala 363:28]
  wire  _GEN_6271 = branchEvalIn_fired ? _GEN_5621 : _GEN_1165; // @[decode.scala 363:28]
  wire  _GEN_6272 = branchEvalIn_fired ? _GEN_5622 : _GEN_1166; // @[decode.scala 363:28]
  wire  _GEN_6273 = branchEvalIn_fired ? _GEN_5623 : _GEN_1167; // @[decode.scala 363:28]
  wire  _GEN_6274 = branchEvalIn_fired ? _GEN_5624 : _GEN_1168; // @[decode.scala 363:28]
  wire  _GEN_6275 = branchEvalIn_fired ? _GEN_5625 : _GEN_1169; // @[decode.scala 363:28]
  wire [5:0] _GEN_6277 = branchEvalIn_fired ? _GEN_5628 : reservedRegMap1_0; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6278 = branchEvalIn_fired ? _GEN_5629 : reservedRegMap1_1; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6279 = branchEvalIn_fired ? _GEN_5630 : reservedRegMap1_2; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6280 = branchEvalIn_fired ? _GEN_5631 : reservedRegMap1_3; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6281 = branchEvalIn_fired ? _GEN_5632 : reservedRegMap1_4; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6282 = branchEvalIn_fired ? _GEN_5633 : reservedRegMap1_5; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6283 = branchEvalIn_fired ? _GEN_5634 : reservedRegMap1_6; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6284 = branchEvalIn_fired ? _GEN_5635 : reservedRegMap1_7; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6285 = branchEvalIn_fired ? _GEN_5636 : reservedRegMap1_8; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6286 = branchEvalIn_fired ? _GEN_5637 : reservedRegMap1_9; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6287 = branchEvalIn_fired ? _GEN_5638 : reservedRegMap1_10; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6288 = branchEvalIn_fired ? _GEN_5639 : reservedRegMap1_11; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6289 = branchEvalIn_fired ? _GEN_5640 : reservedRegMap1_12; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6290 = branchEvalIn_fired ? _GEN_5641 : reservedRegMap1_13; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6291 = branchEvalIn_fired ? _GEN_5642 : reservedRegMap1_14; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6292 = branchEvalIn_fired ? _GEN_5643 : reservedRegMap1_15; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6293 = branchEvalIn_fired ? _GEN_5644 : reservedRegMap1_16; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6294 = branchEvalIn_fired ? _GEN_5645 : reservedRegMap1_17; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6295 = branchEvalIn_fired ? _GEN_5646 : reservedRegMap1_18; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6296 = branchEvalIn_fired ? _GEN_5647 : reservedRegMap1_19; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6297 = branchEvalIn_fired ? _GEN_5648 : reservedRegMap1_20; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6298 = branchEvalIn_fired ? _GEN_5649 : reservedRegMap1_21; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6299 = branchEvalIn_fired ? _GEN_5650 : reservedRegMap1_22; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6300 = branchEvalIn_fired ? _GEN_5651 : reservedRegMap1_23; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6301 = branchEvalIn_fired ? _GEN_5652 : reservedRegMap1_24; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6302 = branchEvalIn_fired ? _GEN_5653 : reservedRegMap1_25; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6303 = branchEvalIn_fired ? _GEN_5654 : reservedRegMap1_26; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6304 = branchEvalIn_fired ? _GEN_5655 : reservedRegMap1_27; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6305 = branchEvalIn_fired ? _GEN_5656 : reservedRegMap1_28; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6306 = branchEvalIn_fired ? _GEN_5657 : reservedRegMap1_29; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6307 = branchEvalIn_fired ? _GEN_5658 : reservedRegMap1_30; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6308 = branchEvalIn_fired ? _GEN_5659 : reservedRegMap1_31; // @[decode.scala 317:28 363:28]
  wire [5:0] _GEN_6309 = branchEvalIn_fired ? _GEN_5660 : reservedRegMap2_0; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6310 = branchEvalIn_fired ? _GEN_5661 : reservedRegMap2_1; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6311 = branchEvalIn_fired ? _GEN_5662 : reservedRegMap2_2; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6312 = branchEvalIn_fired ? _GEN_5663 : reservedRegMap2_3; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6313 = branchEvalIn_fired ? _GEN_5664 : reservedRegMap2_4; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6314 = branchEvalIn_fired ? _GEN_5665 : reservedRegMap2_5; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6315 = branchEvalIn_fired ? _GEN_5666 : reservedRegMap2_6; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6316 = branchEvalIn_fired ? _GEN_5667 : reservedRegMap2_7; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6317 = branchEvalIn_fired ? _GEN_5668 : reservedRegMap2_8; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6318 = branchEvalIn_fired ? _GEN_5669 : reservedRegMap2_9; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6319 = branchEvalIn_fired ? _GEN_5670 : reservedRegMap2_10; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6320 = branchEvalIn_fired ? _GEN_5671 : reservedRegMap2_11; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6321 = branchEvalIn_fired ? _GEN_5672 : reservedRegMap2_12; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6322 = branchEvalIn_fired ? _GEN_5673 : reservedRegMap2_13; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6323 = branchEvalIn_fired ? _GEN_5674 : reservedRegMap2_14; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6324 = branchEvalIn_fired ? _GEN_5675 : reservedRegMap2_15; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6325 = branchEvalIn_fired ? _GEN_5676 : reservedRegMap2_16; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6326 = branchEvalIn_fired ? _GEN_5677 : reservedRegMap2_17; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6327 = branchEvalIn_fired ? _GEN_5678 : reservedRegMap2_18; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6328 = branchEvalIn_fired ? _GEN_5679 : reservedRegMap2_19; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6329 = branchEvalIn_fired ? _GEN_5680 : reservedRegMap2_20; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6330 = branchEvalIn_fired ? _GEN_5681 : reservedRegMap2_21; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6331 = branchEvalIn_fired ? _GEN_5682 : reservedRegMap2_22; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6332 = branchEvalIn_fired ? _GEN_5683 : reservedRegMap2_23; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6333 = branchEvalIn_fired ? _GEN_5684 : reservedRegMap2_24; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6334 = branchEvalIn_fired ? _GEN_5685 : reservedRegMap2_25; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6335 = branchEvalIn_fired ? _GEN_5686 : reservedRegMap2_26; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6336 = branchEvalIn_fired ? _GEN_5687 : reservedRegMap2_27; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6337 = branchEvalIn_fired ? _GEN_5688 : reservedRegMap2_28; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6338 = branchEvalIn_fired ? _GEN_5689 : reservedRegMap2_29; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6339 = branchEvalIn_fired ? _GEN_5690 : reservedRegMap2_30; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6340 = branchEvalIn_fired ? _GEN_5691 : reservedRegMap2_31; // @[decode.scala 318:28 363:28]
  wire [5:0] _GEN_6341 = branchEvalIn_fired ? _GEN_5692 : reservedRegMap3_0; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6342 = branchEvalIn_fired ? _GEN_5693 : reservedRegMap3_1; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6343 = branchEvalIn_fired ? _GEN_5694 : reservedRegMap3_2; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6344 = branchEvalIn_fired ? _GEN_5695 : reservedRegMap3_3; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6345 = branchEvalIn_fired ? _GEN_5696 : reservedRegMap3_4; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6346 = branchEvalIn_fired ? _GEN_5697 : reservedRegMap3_5; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6347 = branchEvalIn_fired ? _GEN_5698 : reservedRegMap3_6; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6348 = branchEvalIn_fired ? _GEN_5699 : reservedRegMap3_7; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6349 = branchEvalIn_fired ? _GEN_5700 : reservedRegMap3_8; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6350 = branchEvalIn_fired ? _GEN_5701 : reservedRegMap3_9; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6351 = branchEvalIn_fired ? _GEN_5702 : reservedRegMap3_10; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6352 = branchEvalIn_fired ? _GEN_5703 : reservedRegMap3_11; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6353 = branchEvalIn_fired ? _GEN_5704 : reservedRegMap3_12; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6354 = branchEvalIn_fired ? _GEN_5705 : reservedRegMap3_13; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6355 = branchEvalIn_fired ? _GEN_5706 : reservedRegMap3_14; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6356 = branchEvalIn_fired ? _GEN_5707 : reservedRegMap3_15; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6357 = branchEvalIn_fired ? _GEN_5708 : reservedRegMap3_16; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6358 = branchEvalIn_fired ? _GEN_5709 : reservedRegMap3_17; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6359 = branchEvalIn_fired ? _GEN_5710 : reservedRegMap3_18; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6360 = branchEvalIn_fired ? _GEN_5711 : reservedRegMap3_19; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6361 = branchEvalIn_fired ? _GEN_5712 : reservedRegMap3_20; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6362 = branchEvalIn_fired ? _GEN_5713 : reservedRegMap3_21; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6363 = branchEvalIn_fired ? _GEN_5714 : reservedRegMap3_22; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6364 = branchEvalIn_fired ? _GEN_5715 : reservedRegMap3_23; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6365 = branchEvalIn_fired ? _GEN_5716 : reservedRegMap3_24; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6366 = branchEvalIn_fired ? _GEN_5717 : reservedRegMap3_25; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6367 = branchEvalIn_fired ? _GEN_5718 : reservedRegMap3_26; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6368 = branchEvalIn_fired ? _GEN_5719 : reservedRegMap3_27; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6369 = branchEvalIn_fired ? _GEN_5720 : reservedRegMap3_28; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6370 = branchEvalIn_fired ? _GEN_5721 : reservedRegMap3_29; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6371 = branchEvalIn_fired ? _GEN_5722 : reservedRegMap3_30; // @[decode.scala 319:28 363:28]
  wire [5:0] _GEN_6372 = branchEvalIn_fired ? _GEN_5723 : reservedRegMap3_31; // @[decode.scala 319:28 363:28]
  wire  _GEN_6373 = branchEvalIn_fired ? _GEN_5724 : reservedFreeList1_0; // @[decode.scala 363:28 322:30]
  wire  _GEN_6374 = branchEvalIn_fired ? _GEN_5725 : reservedFreeList1_1; // @[decode.scala 363:28 322:30]
  wire  _GEN_6375 = branchEvalIn_fired ? _GEN_5726 : reservedFreeList1_2; // @[decode.scala 363:28 322:30]
  wire  _GEN_6376 = branchEvalIn_fired ? _GEN_5727 : reservedFreeList1_3; // @[decode.scala 363:28 322:30]
  wire  _GEN_6377 = branchEvalIn_fired ? _GEN_5728 : reservedFreeList1_4; // @[decode.scala 363:28 322:30]
  wire  _GEN_6378 = branchEvalIn_fired ? _GEN_5729 : reservedFreeList1_5; // @[decode.scala 363:28 322:30]
  wire  _GEN_6379 = branchEvalIn_fired ? _GEN_5730 : reservedFreeList1_6; // @[decode.scala 363:28 322:30]
  wire  _GEN_6380 = branchEvalIn_fired ? _GEN_5731 : reservedFreeList1_7; // @[decode.scala 363:28 322:30]
  wire  _GEN_6381 = branchEvalIn_fired ? _GEN_5732 : reservedFreeList1_8; // @[decode.scala 363:28 322:30]
  wire  _GEN_6382 = branchEvalIn_fired ? _GEN_5733 : reservedFreeList1_9; // @[decode.scala 363:28 322:30]
  wire  _GEN_6383 = branchEvalIn_fired ? _GEN_5734 : reservedFreeList1_10; // @[decode.scala 363:28 322:30]
  wire  _GEN_6384 = branchEvalIn_fired ? _GEN_5735 : reservedFreeList1_11; // @[decode.scala 363:28 322:30]
  wire  _GEN_6385 = branchEvalIn_fired ? _GEN_5736 : reservedFreeList1_12; // @[decode.scala 363:28 322:30]
  wire  _GEN_6386 = branchEvalIn_fired ? _GEN_5737 : reservedFreeList1_13; // @[decode.scala 363:28 322:30]
  wire  _GEN_6387 = branchEvalIn_fired ? _GEN_5738 : reservedFreeList1_14; // @[decode.scala 363:28 322:30]
  wire  _GEN_6388 = branchEvalIn_fired ? _GEN_5739 : reservedFreeList1_15; // @[decode.scala 363:28 322:30]
  wire  _GEN_6389 = branchEvalIn_fired ? _GEN_5740 : reservedFreeList1_16; // @[decode.scala 363:28 322:30]
  wire  _GEN_6390 = branchEvalIn_fired ? _GEN_5741 : reservedFreeList1_17; // @[decode.scala 363:28 322:30]
  wire  _GEN_6391 = branchEvalIn_fired ? _GEN_5742 : reservedFreeList1_18; // @[decode.scala 363:28 322:30]
  wire  _GEN_6392 = branchEvalIn_fired ? _GEN_5743 : reservedFreeList1_19; // @[decode.scala 363:28 322:30]
  wire  _GEN_6393 = branchEvalIn_fired ? _GEN_5744 : reservedFreeList1_20; // @[decode.scala 363:28 322:30]
  wire  _GEN_6394 = branchEvalIn_fired ? _GEN_5745 : reservedFreeList1_21; // @[decode.scala 363:28 322:30]
  wire  _GEN_6395 = branchEvalIn_fired ? _GEN_5746 : reservedFreeList1_22; // @[decode.scala 363:28 322:30]
  wire  _GEN_6396 = branchEvalIn_fired ? _GEN_5747 : reservedFreeList1_23; // @[decode.scala 363:28 322:30]
  wire  _GEN_6397 = branchEvalIn_fired ? _GEN_5748 : reservedFreeList1_24; // @[decode.scala 363:28 322:30]
  wire  _GEN_6398 = branchEvalIn_fired ? _GEN_5749 : reservedFreeList1_25; // @[decode.scala 363:28 322:30]
  wire  _GEN_6399 = branchEvalIn_fired ? _GEN_5750 : reservedFreeList1_26; // @[decode.scala 363:28 322:30]
  wire  _GEN_6400 = branchEvalIn_fired ? _GEN_5751 : reservedFreeList1_27; // @[decode.scala 363:28 322:30]
  wire  _GEN_6401 = branchEvalIn_fired ? _GEN_5752 : reservedFreeList1_28; // @[decode.scala 363:28 322:30]
  wire  _GEN_6402 = branchEvalIn_fired ? _GEN_5753 : reservedFreeList1_29; // @[decode.scala 363:28 322:30]
  wire  _GEN_6403 = branchEvalIn_fired ? _GEN_5754 : reservedFreeList1_30; // @[decode.scala 363:28 322:30]
  wire  _GEN_6404 = branchEvalIn_fired ? _GEN_5755 : reservedFreeList1_31; // @[decode.scala 363:28 322:30]
  wire  _GEN_6405 = branchEvalIn_fired ? _GEN_5756 : reservedFreeList1_32; // @[decode.scala 363:28 322:30]
  wire  _GEN_6406 = branchEvalIn_fired ? _GEN_5757 : reservedFreeList1_33; // @[decode.scala 363:28 322:30]
  wire  _GEN_6407 = branchEvalIn_fired ? _GEN_5758 : reservedFreeList1_34; // @[decode.scala 363:28 322:30]
  wire  _GEN_6408 = branchEvalIn_fired ? _GEN_5759 : reservedFreeList1_35; // @[decode.scala 363:28 322:30]
  wire  _GEN_6409 = branchEvalIn_fired ? _GEN_5760 : reservedFreeList1_36; // @[decode.scala 363:28 322:30]
  wire  _GEN_6410 = branchEvalIn_fired ? _GEN_5761 : reservedFreeList1_37; // @[decode.scala 363:28 322:30]
  wire  _GEN_6411 = branchEvalIn_fired ? _GEN_5762 : reservedFreeList1_38; // @[decode.scala 363:28 322:30]
  wire  _GEN_6412 = branchEvalIn_fired ? _GEN_5763 : reservedFreeList1_39; // @[decode.scala 363:28 322:30]
  wire  _GEN_6413 = branchEvalIn_fired ? _GEN_5764 : reservedFreeList1_40; // @[decode.scala 363:28 322:30]
  wire  _GEN_6414 = branchEvalIn_fired ? _GEN_5765 : reservedFreeList1_41; // @[decode.scala 363:28 322:30]
  wire  _GEN_6415 = branchEvalIn_fired ? _GEN_5766 : reservedFreeList1_42; // @[decode.scala 363:28 322:30]
  wire  _GEN_6416 = branchEvalIn_fired ? _GEN_5767 : reservedFreeList1_43; // @[decode.scala 363:28 322:30]
  wire  _GEN_6417 = branchEvalIn_fired ? _GEN_5768 : reservedFreeList1_44; // @[decode.scala 363:28 322:30]
  wire  _GEN_6418 = branchEvalIn_fired ? _GEN_5769 : reservedFreeList1_45; // @[decode.scala 363:28 322:30]
  wire  _GEN_6419 = branchEvalIn_fired ? _GEN_5770 : reservedFreeList1_46; // @[decode.scala 363:28 322:30]
  wire  _GEN_6420 = branchEvalIn_fired ? _GEN_5771 : reservedFreeList1_47; // @[decode.scala 363:28 322:30]
  wire  _GEN_6421 = branchEvalIn_fired ? _GEN_5772 : reservedFreeList1_48; // @[decode.scala 363:28 322:30]
  wire  _GEN_6422 = branchEvalIn_fired ? _GEN_5773 : reservedFreeList1_49; // @[decode.scala 363:28 322:30]
  wire  _GEN_6423 = branchEvalIn_fired ? _GEN_5774 : reservedFreeList1_50; // @[decode.scala 363:28 322:30]
  wire  _GEN_6424 = branchEvalIn_fired ? _GEN_5775 : reservedFreeList1_51; // @[decode.scala 363:28 322:30]
  wire  _GEN_6425 = branchEvalIn_fired ? _GEN_5776 : reservedFreeList1_52; // @[decode.scala 363:28 322:30]
  wire  _GEN_6426 = branchEvalIn_fired ? _GEN_5777 : reservedFreeList1_53; // @[decode.scala 363:28 322:30]
  wire  _GEN_6427 = branchEvalIn_fired ? _GEN_5778 : reservedFreeList1_54; // @[decode.scala 363:28 322:30]
  wire  _GEN_6428 = branchEvalIn_fired ? _GEN_5779 : reservedFreeList1_55; // @[decode.scala 363:28 322:30]
  wire  _GEN_6429 = branchEvalIn_fired ? _GEN_5780 : reservedFreeList1_56; // @[decode.scala 363:28 322:30]
  wire  _GEN_6430 = branchEvalIn_fired ? _GEN_5781 : reservedFreeList1_57; // @[decode.scala 363:28 322:30]
  wire  _GEN_6431 = branchEvalIn_fired ? _GEN_5782 : reservedFreeList1_58; // @[decode.scala 363:28 322:30]
  wire  _GEN_6432 = branchEvalIn_fired ? _GEN_5783 : reservedFreeList1_59; // @[decode.scala 363:28 322:30]
  wire  _GEN_6433 = branchEvalIn_fired ? _GEN_5784 : reservedFreeList1_60; // @[decode.scala 363:28 322:30]
  wire  _GEN_6434 = branchEvalIn_fired ? _GEN_5785 : reservedFreeList1_61; // @[decode.scala 363:28 322:30]
  wire  _GEN_6435 = branchEvalIn_fired ? _GEN_5786 : reservedFreeList1_62; // @[decode.scala 363:28 322:30]
  wire  _GEN_6437 = branchEvalIn_fired ? _GEN_5788 : reservedFreeList2_0; // @[decode.scala 363:28 323:30]
  wire  _GEN_6438 = branchEvalIn_fired ? _GEN_5789 : reservedFreeList2_1; // @[decode.scala 363:28 323:30]
  wire  _GEN_6439 = branchEvalIn_fired ? _GEN_5790 : reservedFreeList2_2; // @[decode.scala 363:28 323:30]
  wire  _GEN_6440 = branchEvalIn_fired ? _GEN_5791 : reservedFreeList2_3; // @[decode.scala 363:28 323:30]
  wire  _GEN_6441 = branchEvalIn_fired ? _GEN_5792 : reservedFreeList2_4; // @[decode.scala 363:28 323:30]
  wire  _GEN_6442 = branchEvalIn_fired ? _GEN_5793 : reservedFreeList2_5; // @[decode.scala 363:28 323:30]
  wire  _GEN_6443 = branchEvalIn_fired ? _GEN_5794 : reservedFreeList2_6; // @[decode.scala 363:28 323:30]
  wire  _GEN_6444 = branchEvalIn_fired ? _GEN_5795 : reservedFreeList2_7; // @[decode.scala 363:28 323:30]
  wire  _GEN_6445 = branchEvalIn_fired ? _GEN_5796 : reservedFreeList2_8; // @[decode.scala 363:28 323:30]
  wire  _GEN_6446 = branchEvalIn_fired ? _GEN_5797 : reservedFreeList2_9; // @[decode.scala 363:28 323:30]
  wire  _GEN_6447 = branchEvalIn_fired ? _GEN_5798 : reservedFreeList2_10; // @[decode.scala 363:28 323:30]
  wire  _GEN_6448 = branchEvalIn_fired ? _GEN_5799 : reservedFreeList2_11; // @[decode.scala 363:28 323:30]
  wire  _GEN_6449 = branchEvalIn_fired ? _GEN_5800 : reservedFreeList2_12; // @[decode.scala 363:28 323:30]
  wire  _GEN_6450 = branchEvalIn_fired ? _GEN_5801 : reservedFreeList2_13; // @[decode.scala 363:28 323:30]
  wire  _GEN_6451 = branchEvalIn_fired ? _GEN_5802 : reservedFreeList2_14; // @[decode.scala 363:28 323:30]
  wire  _GEN_6452 = branchEvalIn_fired ? _GEN_5803 : reservedFreeList2_15; // @[decode.scala 363:28 323:30]
  wire  _GEN_6453 = branchEvalIn_fired ? _GEN_5804 : reservedFreeList2_16; // @[decode.scala 363:28 323:30]
  wire  _GEN_6454 = branchEvalIn_fired ? _GEN_5805 : reservedFreeList2_17; // @[decode.scala 363:28 323:30]
  wire  _GEN_6455 = branchEvalIn_fired ? _GEN_5806 : reservedFreeList2_18; // @[decode.scala 363:28 323:30]
  wire  _GEN_6456 = branchEvalIn_fired ? _GEN_5807 : reservedFreeList2_19; // @[decode.scala 363:28 323:30]
  wire  _GEN_6457 = branchEvalIn_fired ? _GEN_5808 : reservedFreeList2_20; // @[decode.scala 363:28 323:30]
  wire  _GEN_6458 = branchEvalIn_fired ? _GEN_5809 : reservedFreeList2_21; // @[decode.scala 363:28 323:30]
  wire  _GEN_6459 = branchEvalIn_fired ? _GEN_5810 : reservedFreeList2_22; // @[decode.scala 363:28 323:30]
  wire  _GEN_6460 = branchEvalIn_fired ? _GEN_5811 : reservedFreeList2_23; // @[decode.scala 363:28 323:30]
  wire  _GEN_6461 = branchEvalIn_fired ? _GEN_5812 : reservedFreeList2_24; // @[decode.scala 363:28 323:30]
  wire  _GEN_6462 = branchEvalIn_fired ? _GEN_5813 : reservedFreeList2_25; // @[decode.scala 363:28 323:30]
  wire  _GEN_6463 = branchEvalIn_fired ? _GEN_5814 : reservedFreeList2_26; // @[decode.scala 363:28 323:30]
  wire  _GEN_6464 = branchEvalIn_fired ? _GEN_5815 : reservedFreeList2_27; // @[decode.scala 363:28 323:30]
  wire  _GEN_6465 = branchEvalIn_fired ? _GEN_5816 : reservedFreeList2_28; // @[decode.scala 363:28 323:30]
  wire  _GEN_6466 = branchEvalIn_fired ? _GEN_5817 : reservedFreeList2_29; // @[decode.scala 363:28 323:30]
  wire  _GEN_6467 = branchEvalIn_fired ? _GEN_5818 : reservedFreeList2_30; // @[decode.scala 363:28 323:30]
  wire  _GEN_6468 = branchEvalIn_fired ? _GEN_5819 : reservedFreeList2_31; // @[decode.scala 363:28 323:30]
  wire  _GEN_6469 = branchEvalIn_fired ? _GEN_5820 : reservedFreeList2_32; // @[decode.scala 363:28 323:30]
  wire  _GEN_6470 = branchEvalIn_fired ? _GEN_5821 : reservedFreeList2_33; // @[decode.scala 363:28 323:30]
  wire  _GEN_6471 = branchEvalIn_fired ? _GEN_5822 : reservedFreeList2_34; // @[decode.scala 363:28 323:30]
  wire  _GEN_6472 = branchEvalIn_fired ? _GEN_5823 : reservedFreeList2_35; // @[decode.scala 363:28 323:30]
  wire  _GEN_6473 = branchEvalIn_fired ? _GEN_5824 : reservedFreeList2_36; // @[decode.scala 363:28 323:30]
  wire  _GEN_6474 = branchEvalIn_fired ? _GEN_5825 : reservedFreeList2_37; // @[decode.scala 363:28 323:30]
  wire  _GEN_6475 = branchEvalIn_fired ? _GEN_5826 : reservedFreeList2_38; // @[decode.scala 363:28 323:30]
  wire  _GEN_6476 = branchEvalIn_fired ? _GEN_5827 : reservedFreeList2_39; // @[decode.scala 363:28 323:30]
  wire  _GEN_6477 = branchEvalIn_fired ? _GEN_5828 : reservedFreeList2_40; // @[decode.scala 363:28 323:30]
  wire  _GEN_6478 = branchEvalIn_fired ? _GEN_5829 : reservedFreeList2_41; // @[decode.scala 363:28 323:30]
  wire  _GEN_6479 = branchEvalIn_fired ? _GEN_5830 : reservedFreeList2_42; // @[decode.scala 363:28 323:30]
  wire  _GEN_6480 = branchEvalIn_fired ? _GEN_5831 : reservedFreeList2_43; // @[decode.scala 363:28 323:30]
  wire  _GEN_6481 = branchEvalIn_fired ? _GEN_5832 : reservedFreeList2_44; // @[decode.scala 363:28 323:30]
  wire  _GEN_6482 = branchEvalIn_fired ? _GEN_5833 : reservedFreeList2_45; // @[decode.scala 363:28 323:30]
  wire  _GEN_6483 = branchEvalIn_fired ? _GEN_5834 : reservedFreeList2_46; // @[decode.scala 363:28 323:30]
  wire  _GEN_6484 = branchEvalIn_fired ? _GEN_5835 : reservedFreeList2_47; // @[decode.scala 363:28 323:30]
  wire  _GEN_6485 = branchEvalIn_fired ? _GEN_5836 : reservedFreeList2_48; // @[decode.scala 363:28 323:30]
  wire  _GEN_6486 = branchEvalIn_fired ? _GEN_5837 : reservedFreeList2_49; // @[decode.scala 363:28 323:30]
  wire  _GEN_6487 = branchEvalIn_fired ? _GEN_5838 : reservedFreeList2_50; // @[decode.scala 363:28 323:30]
  wire  _GEN_6488 = branchEvalIn_fired ? _GEN_5839 : reservedFreeList2_51; // @[decode.scala 363:28 323:30]
  wire  _GEN_6489 = branchEvalIn_fired ? _GEN_5840 : reservedFreeList2_52; // @[decode.scala 363:28 323:30]
  wire  _GEN_6490 = branchEvalIn_fired ? _GEN_5841 : reservedFreeList2_53; // @[decode.scala 363:28 323:30]
  wire  _GEN_6491 = branchEvalIn_fired ? _GEN_5842 : reservedFreeList2_54; // @[decode.scala 363:28 323:30]
  wire  _GEN_6492 = branchEvalIn_fired ? _GEN_5843 : reservedFreeList2_55; // @[decode.scala 363:28 323:30]
  wire  _GEN_6493 = branchEvalIn_fired ? _GEN_5844 : reservedFreeList2_56; // @[decode.scala 363:28 323:30]
  wire  _GEN_6494 = branchEvalIn_fired ? _GEN_5845 : reservedFreeList2_57; // @[decode.scala 363:28 323:30]
  wire  _GEN_6495 = branchEvalIn_fired ? _GEN_5846 : reservedFreeList2_58; // @[decode.scala 363:28 323:30]
  wire  _GEN_6496 = branchEvalIn_fired ? _GEN_5847 : reservedFreeList2_59; // @[decode.scala 363:28 323:30]
  wire  _GEN_6497 = branchEvalIn_fired ? _GEN_5848 : reservedFreeList2_60; // @[decode.scala 363:28 323:30]
  wire  _GEN_6498 = branchEvalIn_fired ? _GEN_5849 : reservedFreeList2_61; // @[decode.scala 363:28 323:30]
  wire  _GEN_6499 = branchEvalIn_fired ? _GEN_5850 : reservedFreeList2_62; // @[decode.scala 363:28 323:30]
  wire  _GEN_6501 = branchEvalIn_fired ? _GEN_5852 : reservedFreeList3_0; // @[decode.scala 363:28 324:30]
  wire  _GEN_6502 = branchEvalIn_fired ? _GEN_5853 : reservedFreeList3_1; // @[decode.scala 363:28 324:30]
  wire  _GEN_6503 = branchEvalIn_fired ? _GEN_5854 : reservedFreeList3_2; // @[decode.scala 363:28 324:30]
  wire  _GEN_6504 = branchEvalIn_fired ? _GEN_5855 : reservedFreeList3_3; // @[decode.scala 363:28 324:30]
  wire  _GEN_6505 = branchEvalIn_fired ? _GEN_5856 : reservedFreeList3_4; // @[decode.scala 363:28 324:30]
  wire  _GEN_6506 = branchEvalIn_fired ? _GEN_5857 : reservedFreeList3_5; // @[decode.scala 363:28 324:30]
  wire  _GEN_6507 = branchEvalIn_fired ? _GEN_5858 : reservedFreeList3_6; // @[decode.scala 363:28 324:30]
  wire  _GEN_6508 = branchEvalIn_fired ? _GEN_5859 : reservedFreeList3_7; // @[decode.scala 363:28 324:30]
  wire  _GEN_6509 = branchEvalIn_fired ? _GEN_5860 : reservedFreeList3_8; // @[decode.scala 363:28 324:30]
  wire  _GEN_6510 = branchEvalIn_fired ? _GEN_5861 : reservedFreeList3_9; // @[decode.scala 363:28 324:30]
  wire  _GEN_6511 = branchEvalIn_fired ? _GEN_5862 : reservedFreeList3_10; // @[decode.scala 363:28 324:30]
  wire  _GEN_6512 = branchEvalIn_fired ? _GEN_5863 : reservedFreeList3_11; // @[decode.scala 363:28 324:30]
  wire  _GEN_6513 = branchEvalIn_fired ? _GEN_5864 : reservedFreeList3_12; // @[decode.scala 363:28 324:30]
  wire  _GEN_6514 = branchEvalIn_fired ? _GEN_5865 : reservedFreeList3_13; // @[decode.scala 363:28 324:30]
  wire  _GEN_6515 = branchEvalIn_fired ? _GEN_5866 : reservedFreeList3_14; // @[decode.scala 363:28 324:30]
  wire  _GEN_6516 = branchEvalIn_fired ? _GEN_5867 : reservedFreeList3_15; // @[decode.scala 363:28 324:30]
  wire  _GEN_6517 = branchEvalIn_fired ? _GEN_5868 : reservedFreeList3_16; // @[decode.scala 363:28 324:30]
  wire  _GEN_6518 = branchEvalIn_fired ? _GEN_5869 : reservedFreeList3_17; // @[decode.scala 363:28 324:30]
  wire  _GEN_6519 = branchEvalIn_fired ? _GEN_5870 : reservedFreeList3_18; // @[decode.scala 363:28 324:30]
  wire  _GEN_6520 = branchEvalIn_fired ? _GEN_5871 : reservedFreeList3_19; // @[decode.scala 363:28 324:30]
  wire  _GEN_6521 = branchEvalIn_fired ? _GEN_5872 : reservedFreeList3_20; // @[decode.scala 363:28 324:30]
  wire  _GEN_6522 = branchEvalIn_fired ? _GEN_5873 : reservedFreeList3_21; // @[decode.scala 363:28 324:30]
  wire  _GEN_6523 = branchEvalIn_fired ? _GEN_5874 : reservedFreeList3_22; // @[decode.scala 363:28 324:30]
  wire  _GEN_6524 = branchEvalIn_fired ? _GEN_5875 : reservedFreeList3_23; // @[decode.scala 363:28 324:30]
  wire  _GEN_6525 = branchEvalIn_fired ? _GEN_5876 : reservedFreeList3_24; // @[decode.scala 363:28 324:30]
  wire  _GEN_6526 = branchEvalIn_fired ? _GEN_5877 : reservedFreeList3_25; // @[decode.scala 363:28 324:30]
  wire  _GEN_6527 = branchEvalIn_fired ? _GEN_5878 : reservedFreeList3_26; // @[decode.scala 363:28 324:30]
  wire  _GEN_6528 = branchEvalIn_fired ? _GEN_5879 : reservedFreeList3_27; // @[decode.scala 363:28 324:30]
  wire  _GEN_6529 = branchEvalIn_fired ? _GEN_5880 : reservedFreeList3_28; // @[decode.scala 363:28 324:30]
  wire  _GEN_6530 = branchEvalIn_fired ? _GEN_5881 : reservedFreeList3_29; // @[decode.scala 363:28 324:30]
  wire  _GEN_6531 = branchEvalIn_fired ? _GEN_5882 : reservedFreeList3_30; // @[decode.scala 363:28 324:30]
  wire  _GEN_6532 = branchEvalIn_fired ? _GEN_5883 : reservedFreeList3_31; // @[decode.scala 363:28 324:30]
  wire  _GEN_6533 = branchEvalIn_fired ? _GEN_5884 : reservedFreeList3_32; // @[decode.scala 363:28 324:30]
  wire  _GEN_6534 = branchEvalIn_fired ? _GEN_5885 : reservedFreeList3_33; // @[decode.scala 363:28 324:30]
  wire  _GEN_6535 = branchEvalIn_fired ? _GEN_5886 : reservedFreeList3_34; // @[decode.scala 363:28 324:30]
  wire  _GEN_6536 = branchEvalIn_fired ? _GEN_5887 : reservedFreeList3_35; // @[decode.scala 363:28 324:30]
  wire  _GEN_6537 = branchEvalIn_fired ? _GEN_5888 : reservedFreeList3_36; // @[decode.scala 363:28 324:30]
  wire  _GEN_6538 = branchEvalIn_fired ? _GEN_5889 : reservedFreeList3_37; // @[decode.scala 363:28 324:30]
  wire  _GEN_6539 = branchEvalIn_fired ? _GEN_5890 : reservedFreeList3_38; // @[decode.scala 363:28 324:30]
  wire  _GEN_6540 = branchEvalIn_fired ? _GEN_5891 : reservedFreeList3_39; // @[decode.scala 363:28 324:30]
  wire  _GEN_6541 = branchEvalIn_fired ? _GEN_5892 : reservedFreeList3_40; // @[decode.scala 363:28 324:30]
  wire  _GEN_6542 = branchEvalIn_fired ? _GEN_5893 : reservedFreeList3_41; // @[decode.scala 363:28 324:30]
  wire  _GEN_6543 = branchEvalIn_fired ? _GEN_5894 : reservedFreeList3_42; // @[decode.scala 363:28 324:30]
  wire  _GEN_6544 = branchEvalIn_fired ? _GEN_5895 : reservedFreeList3_43; // @[decode.scala 363:28 324:30]
  wire  _GEN_6545 = branchEvalIn_fired ? _GEN_5896 : reservedFreeList3_44; // @[decode.scala 363:28 324:30]
  wire  _GEN_6546 = branchEvalIn_fired ? _GEN_5897 : reservedFreeList3_45; // @[decode.scala 363:28 324:30]
  wire  _GEN_6547 = branchEvalIn_fired ? _GEN_5898 : reservedFreeList3_46; // @[decode.scala 363:28 324:30]
  wire  _GEN_6548 = branchEvalIn_fired ? _GEN_5899 : reservedFreeList3_47; // @[decode.scala 363:28 324:30]
  wire  _GEN_6549 = branchEvalIn_fired ? _GEN_5900 : reservedFreeList3_48; // @[decode.scala 363:28 324:30]
  wire  _GEN_6550 = branchEvalIn_fired ? _GEN_5901 : reservedFreeList3_49; // @[decode.scala 363:28 324:30]
  wire  _GEN_6551 = branchEvalIn_fired ? _GEN_5902 : reservedFreeList3_50; // @[decode.scala 363:28 324:30]
  wire  _GEN_6552 = branchEvalIn_fired ? _GEN_5903 : reservedFreeList3_51; // @[decode.scala 363:28 324:30]
  wire  _GEN_6553 = branchEvalIn_fired ? _GEN_5904 : reservedFreeList3_52; // @[decode.scala 363:28 324:30]
  wire  _GEN_6554 = branchEvalIn_fired ? _GEN_5905 : reservedFreeList3_53; // @[decode.scala 363:28 324:30]
  wire  _GEN_6555 = branchEvalIn_fired ? _GEN_5906 : reservedFreeList3_54; // @[decode.scala 363:28 324:30]
  wire  _GEN_6556 = branchEvalIn_fired ? _GEN_5907 : reservedFreeList3_55; // @[decode.scala 363:28 324:30]
  wire  _GEN_6557 = branchEvalIn_fired ? _GEN_5908 : reservedFreeList3_56; // @[decode.scala 363:28 324:30]
  wire  _GEN_6558 = branchEvalIn_fired ? _GEN_5909 : reservedFreeList3_57; // @[decode.scala 363:28 324:30]
  wire  _GEN_6559 = branchEvalIn_fired ? _GEN_5910 : reservedFreeList3_58; // @[decode.scala 363:28 324:30]
  wire  _GEN_6560 = branchEvalIn_fired ? _GEN_5911 : reservedFreeList3_59; // @[decode.scala 363:28 324:30]
  wire  _GEN_6561 = branchEvalIn_fired ? _GEN_5912 : reservedFreeList3_60; // @[decode.scala 363:28 324:30]
  wire  _GEN_6562 = branchEvalIn_fired ? _GEN_5913 : reservedFreeList3_61; // @[decode.scala 363:28 324:30]
  wire  _GEN_6563 = branchEvalIn_fired ? _GEN_5914 : reservedFreeList3_62; // @[decode.scala 363:28 324:30]
  wire  _GEN_6565 = branchEvalIn_fired ? _GEN_5916 : reservedValidList1_0; // @[decode.scala 363:28 327:31]
  wire  _GEN_6566 = branchEvalIn_fired ? _GEN_5917 : reservedValidList1_1; // @[decode.scala 363:28 327:31]
  wire  _GEN_6567 = branchEvalIn_fired ? _GEN_5918 : reservedValidList1_2; // @[decode.scala 363:28 327:31]
  wire  _GEN_6568 = branchEvalIn_fired ? _GEN_5919 : reservedValidList1_3; // @[decode.scala 363:28 327:31]
  wire  _GEN_6569 = branchEvalIn_fired ? _GEN_5920 : reservedValidList1_4; // @[decode.scala 363:28 327:31]
  wire  _GEN_6570 = branchEvalIn_fired ? _GEN_5921 : reservedValidList1_5; // @[decode.scala 363:28 327:31]
  wire  _GEN_6571 = branchEvalIn_fired ? _GEN_5922 : reservedValidList1_6; // @[decode.scala 363:28 327:31]
  wire  _GEN_6572 = branchEvalIn_fired ? _GEN_5923 : reservedValidList1_7; // @[decode.scala 363:28 327:31]
  wire  _GEN_6573 = branchEvalIn_fired ? _GEN_5924 : reservedValidList1_8; // @[decode.scala 363:28 327:31]
  wire  _GEN_6574 = branchEvalIn_fired ? _GEN_5925 : reservedValidList1_9; // @[decode.scala 363:28 327:31]
  wire  _GEN_6575 = branchEvalIn_fired ? _GEN_5926 : reservedValidList1_10; // @[decode.scala 363:28 327:31]
  wire  _GEN_6576 = branchEvalIn_fired ? _GEN_5927 : reservedValidList1_11; // @[decode.scala 363:28 327:31]
  wire  _GEN_6577 = branchEvalIn_fired ? _GEN_5928 : reservedValidList1_12; // @[decode.scala 363:28 327:31]
  wire  _GEN_6578 = branchEvalIn_fired ? _GEN_5929 : reservedValidList1_13; // @[decode.scala 363:28 327:31]
  wire  _GEN_6579 = branchEvalIn_fired ? _GEN_5930 : reservedValidList1_14; // @[decode.scala 363:28 327:31]
  wire  _GEN_6580 = branchEvalIn_fired ? _GEN_5931 : reservedValidList1_15; // @[decode.scala 363:28 327:31]
  wire  _GEN_6581 = branchEvalIn_fired ? _GEN_5932 : reservedValidList1_16; // @[decode.scala 363:28 327:31]
  wire  _GEN_6582 = branchEvalIn_fired ? _GEN_5933 : reservedValidList1_17; // @[decode.scala 363:28 327:31]
  wire  _GEN_6583 = branchEvalIn_fired ? _GEN_5934 : reservedValidList1_18; // @[decode.scala 363:28 327:31]
  wire  _GEN_6584 = branchEvalIn_fired ? _GEN_5935 : reservedValidList1_19; // @[decode.scala 363:28 327:31]
  wire  _GEN_6585 = branchEvalIn_fired ? _GEN_5936 : reservedValidList1_20; // @[decode.scala 363:28 327:31]
  wire  _GEN_6586 = branchEvalIn_fired ? _GEN_5937 : reservedValidList1_21; // @[decode.scala 363:28 327:31]
  wire  _GEN_6587 = branchEvalIn_fired ? _GEN_5938 : reservedValidList1_22; // @[decode.scala 363:28 327:31]
  wire  _GEN_6588 = branchEvalIn_fired ? _GEN_5939 : reservedValidList1_23; // @[decode.scala 363:28 327:31]
  wire  _GEN_6589 = branchEvalIn_fired ? _GEN_5940 : reservedValidList1_24; // @[decode.scala 363:28 327:31]
  wire  _GEN_6590 = branchEvalIn_fired ? _GEN_5941 : reservedValidList1_25; // @[decode.scala 363:28 327:31]
  wire  _GEN_6591 = branchEvalIn_fired ? _GEN_5942 : reservedValidList1_26; // @[decode.scala 363:28 327:31]
  wire  _GEN_6592 = branchEvalIn_fired ? _GEN_5943 : reservedValidList1_27; // @[decode.scala 363:28 327:31]
  wire  _GEN_6593 = branchEvalIn_fired ? _GEN_5944 : reservedValidList1_28; // @[decode.scala 363:28 327:31]
  wire  _GEN_6594 = branchEvalIn_fired ? _GEN_5945 : reservedValidList1_29; // @[decode.scala 363:28 327:31]
  wire  _GEN_6595 = branchEvalIn_fired ? _GEN_5946 : reservedValidList1_30; // @[decode.scala 363:28 327:31]
  wire  _GEN_6596 = branchEvalIn_fired ? _GEN_5947 : reservedValidList1_31; // @[decode.scala 363:28 327:31]
  wire  _GEN_6597 = branchEvalIn_fired ? _GEN_5948 : reservedValidList1_32; // @[decode.scala 363:28 327:31]
  wire  _GEN_6598 = branchEvalIn_fired ? _GEN_5949 : reservedValidList1_33; // @[decode.scala 363:28 327:31]
  wire  _GEN_6599 = branchEvalIn_fired ? _GEN_5950 : reservedValidList1_34; // @[decode.scala 363:28 327:31]
  wire  _GEN_6600 = branchEvalIn_fired ? _GEN_5951 : reservedValidList1_35; // @[decode.scala 363:28 327:31]
  wire  _GEN_6601 = branchEvalIn_fired ? _GEN_5952 : reservedValidList1_36; // @[decode.scala 363:28 327:31]
  wire  _GEN_6602 = branchEvalIn_fired ? _GEN_5953 : reservedValidList1_37; // @[decode.scala 363:28 327:31]
  wire  _GEN_6603 = branchEvalIn_fired ? _GEN_5954 : reservedValidList1_38; // @[decode.scala 363:28 327:31]
  wire  _GEN_6604 = branchEvalIn_fired ? _GEN_5955 : reservedValidList1_39; // @[decode.scala 363:28 327:31]
  wire  _GEN_6605 = branchEvalIn_fired ? _GEN_5956 : reservedValidList1_40; // @[decode.scala 363:28 327:31]
  wire  _GEN_6606 = branchEvalIn_fired ? _GEN_5957 : reservedValidList1_41; // @[decode.scala 363:28 327:31]
  wire  _GEN_6607 = branchEvalIn_fired ? _GEN_5958 : reservedValidList1_42; // @[decode.scala 363:28 327:31]
  wire  _GEN_6608 = branchEvalIn_fired ? _GEN_5959 : reservedValidList1_43; // @[decode.scala 363:28 327:31]
  wire  _GEN_6609 = branchEvalIn_fired ? _GEN_5960 : reservedValidList1_44; // @[decode.scala 363:28 327:31]
  wire  _GEN_6610 = branchEvalIn_fired ? _GEN_5961 : reservedValidList1_45; // @[decode.scala 363:28 327:31]
  wire  _GEN_6611 = branchEvalIn_fired ? _GEN_5962 : reservedValidList1_46; // @[decode.scala 363:28 327:31]
  wire  _GEN_6612 = branchEvalIn_fired ? _GEN_5963 : reservedValidList1_47; // @[decode.scala 363:28 327:31]
  wire  _GEN_6613 = branchEvalIn_fired ? _GEN_5964 : reservedValidList1_48; // @[decode.scala 363:28 327:31]
  wire  _GEN_6614 = branchEvalIn_fired ? _GEN_5965 : reservedValidList1_49; // @[decode.scala 363:28 327:31]
  wire  _GEN_6615 = branchEvalIn_fired ? _GEN_5966 : reservedValidList1_50; // @[decode.scala 363:28 327:31]
  wire  _GEN_6616 = branchEvalIn_fired ? _GEN_5967 : reservedValidList1_51; // @[decode.scala 363:28 327:31]
  wire  _GEN_6617 = branchEvalIn_fired ? _GEN_5968 : reservedValidList1_52; // @[decode.scala 363:28 327:31]
  wire  _GEN_6618 = branchEvalIn_fired ? _GEN_5969 : reservedValidList1_53; // @[decode.scala 363:28 327:31]
  wire  _GEN_6619 = branchEvalIn_fired ? _GEN_5970 : reservedValidList1_54; // @[decode.scala 363:28 327:31]
  wire  _GEN_6620 = branchEvalIn_fired ? _GEN_5971 : reservedValidList1_55; // @[decode.scala 363:28 327:31]
  wire  _GEN_6621 = branchEvalIn_fired ? _GEN_5972 : reservedValidList1_56; // @[decode.scala 363:28 327:31]
  wire  _GEN_6622 = branchEvalIn_fired ? _GEN_5973 : reservedValidList1_57; // @[decode.scala 363:28 327:31]
  wire  _GEN_6623 = branchEvalIn_fired ? _GEN_5974 : reservedValidList1_58; // @[decode.scala 363:28 327:31]
  wire  _GEN_6624 = branchEvalIn_fired ? _GEN_5975 : reservedValidList1_59; // @[decode.scala 363:28 327:31]
  wire  _GEN_6625 = branchEvalIn_fired ? _GEN_5976 : reservedValidList1_60; // @[decode.scala 363:28 327:31]
  wire  _GEN_6626 = branchEvalIn_fired ? _GEN_5977 : reservedValidList1_61; // @[decode.scala 363:28 327:31]
  wire  _GEN_6627 = branchEvalIn_fired ? _GEN_5978 : reservedValidList1_62; // @[decode.scala 363:28 327:31]
  wire  _GEN_6628 = branchEvalIn_fired ? _GEN_5979 : reservedValidList1_63; // @[decode.scala 363:28 327:31]
  wire  _GEN_6629 = branchEvalIn_fired ? _GEN_5980 : reservedValidList2_0; // @[decode.scala 363:28 328:31]
  wire  _GEN_6630 = branchEvalIn_fired ? _GEN_5981 : reservedValidList2_1; // @[decode.scala 363:28 328:31]
  wire  _GEN_6631 = branchEvalIn_fired ? _GEN_5982 : reservedValidList2_2; // @[decode.scala 363:28 328:31]
  wire  _GEN_6632 = branchEvalIn_fired ? _GEN_5983 : reservedValidList2_3; // @[decode.scala 363:28 328:31]
  wire  _GEN_6633 = branchEvalIn_fired ? _GEN_5984 : reservedValidList2_4; // @[decode.scala 363:28 328:31]
  wire  _GEN_6634 = branchEvalIn_fired ? _GEN_5985 : reservedValidList2_5; // @[decode.scala 363:28 328:31]
  wire  _GEN_6635 = branchEvalIn_fired ? _GEN_5986 : reservedValidList2_6; // @[decode.scala 363:28 328:31]
  wire  _GEN_6636 = branchEvalIn_fired ? _GEN_5987 : reservedValidList2_7; // @[decode.scala 363:28 328:31]
  wire  _GEN_6637 = branchEvalIn_fired ? _GEN_5988 : reservedValidList2_8; // @[decode.scala 363:28 328:31]
  wire  _GEN_6638 = branchEvalIn_fired ? _GEN_5989 : reservedValidList2_9; // @[decode.scala 363:28 328:31]
  wire  _GEN_6639 = branchEvalIn_fired ? _GEN_5990 : reservedValidList2_10; // @[decode.scala 363:28 328:31]
  wire  _GEN_6640 = branchEvalIn_fired ? _GEN_5991 : reservedValidList2_11; // @[decode.scala 363:28 328:31]
  wire  _GEN_6641 = branchEvalIn_fired ? _GEN_5992 : reservedValidList2_12; // @[decode.scala 363:28 328:31]
  wire  _GEN_6642 = branchEvalIn_fired ? _GEN_5993 : reservedValidList2_13; // @[decode.scala 363:28 328:31]
  wire  _GEN_6643 = branchEvalIn_fired ? _GEN_5994 : reservedValidList2_14; // @[decode.scala 363:28 328:31]
  wire  _GEN_6644 = branchEvalIn_fired ? _GEN_5995 : reservedValidList2_15; // @[decode.scala 363:28 328:31]
  wire  _GEN_6645 = branchEvalIn_fired ? _GEN_5996 : reservedValidList2_16; // @[decode.scala 363:28 328:31]
  wire  _GEN_6646 = branchEvalIn_fired ? _GEN_5997 : reservedValidList2_17; // @[decode.scala 363:28 328:31]
  wire  _GEN_6647 = branchEvalIn_fired ? _GEN_5998 : reservedValidList2_18; // @[decode.scala 363:28 328:31]
  wire  _GEN_6648 = branchEvalIn_fired ? _GEN_5999 : reservedValidList2_19; // @[decode.scala 363:28 328:31]
  wire  _GEN_6649 = branchEvalIn_fired ? _GEN_6000 : reservedValidList2_20; // @[decode.scala 363:28 328:31]
  wire  _GEN_6650 = branchEvalIn_fired ? _GEN_6001 : reservedValidList2_21; // @[decode.scala 363:28 328:31]
  wire  _GEN_6651 = branchEvalIn_fired ? _GEN_6002 : reservedValidList2_22; // @[decode.scala 363:28 328:31]
  wire  _GEN_6652 = branchEvalIn_fired ? _GEN_6003 : reservedValidList2_23; // @[decode.scala 363:28 328:31]
  wire  _GEN_6653 = branchEvalIn_fired ? _GEN_6004 : reservedValidList2_24; // @[decode.scala 363:28 328:31]
  wire  _GEN_6654 = branchEvalIn_fired ? _GEN_6005 : reservedValidList2_25; // @[decode.scala 363:28 328:31]
  wire  _GEN_6655 = branchEvalIn_fired ? _GEN_6006 : reservedValidList2_26; // @[decode.scala 363:28 328:31]
  wire  _GEN_6656 = branchEvalIn_fired ? _GEN_6007 : reservedValidList2_27; // @[decode.scala 363:28 328:31]
  wire  _GEN_6657 = branchEvalIn_fired ? _GEN_6008 : reservedValidList2_28; // @[decode.scala 363:28 328:31]
  wire  _GEN_6658 = branchEvalIn_fired ? _GEN_6009 : reservedValidList2_29; // @[decode.scala 363:28 328:31]
  wire  _GEN_6659 = branchEvalIn_fired ? _GEN_6010 : reservedValidList2_30; // @[decode.scala 363:28 328:31]
  wire  _GEN_6660 = branchEvalIn_fired ? _GEN_6011 : reservedValidList2_31; // @[decode.scala 363:28 328:31]
  wire  _GEN_6661 = branchEvalIn_fired ? _GEN_6012 : reservedValidList2_32; // @[decode.scala 363:28 328:31]
  wire  _GEN_6662 = branchEvalIn_fired ? _GEN_6013 : reservedValidList2_33; // @[decode.scala 363:28 328:31]
  wire  _GEN_6663 = branchEvalIn_fired ? _GEN_6014 : reservedValidList2_34; // @[decode.scala 363:28 328:31]
  wire  _GEN_6664 = branchEvalIn_fired ? _GEN_6015 : reservedValidList2_35; // @[decode.scala 363:28 328:31]
  wire  _GEN_6665 = branchEvalIn_fired ? _GEN_6016 : reservedValidList2_36; // @[decode.scala 363:28 328:31]
  wire  _GEN_6666 = branchEvalIn_fired ? _GEN_6017 : reservedValidList2_37; // @[decode.scala 363:28 328:31]
  wire  _GEN_6667 = branchEvalIn_fired ? _GEN_6018 : reservedValidList2_38; // @[decode.scala 363:28 328:31]
  wire  _GEN_6668 = branchEvalIn_fired ? _GEN_6019 : reservedValidList2_39; // @[decode.scala 363:28 328:31]
  wire  _GEN_6669 = branchEvalIn_fired ? _GEN_6020 : reservedValidList2_40; // @[decode.scala 363:28 328:31]
  wire  _GEN_6670 = branchEvalIn_fired ? _GEN_6021 : reservedValidList2_41; // @[decode.scala 363:28 328:31]
  wire  _GEN_6671 = branchEvalIn_fired ? _GEN_6022 : reservedValidList2_42; // @[decode.scala 363:28 328:31]
  wire  _GEN_6672 = branchEvalIn_fired ? _GEN_6023 : reservedValidList2_43; // @[decode.scala 363:28 328:31]
  wire  _GEN_6673 = branchEvalIn_fired ? _GEN_6024 : reservedValidList2_44; // @[decode.scala 363:28 328:31]
  wire  _GEN_6674 = branchEvalIn_fired ? _GEN_6025 : reservedValidList2_45; // @[decode.scala 363:28 328:31]
  wire  _GEN_6675 = branchEvalIn_fired ? _GEN_6026 : reservedValidList2_46; // @[decode.scala 363:28 328:31]
  wire  _GEN_6676 = branchEvalIn_fired ? _GEN_6027 : reservedValidList2_47; // @[decode.scala 363:28 328:31]
  wire  _GEN_6677 = branchEvalIn_fired ? _GEN_6028 : reservedValidList2_48; // @[decode.scala 363:28 328:31]
  wire  _GEN_6678 = branchEvalIn_fired ? _GEN_6029 : reservedValidList2_49; // @[decode.scala 363:28 328:31]
  wire  _GEN_6679 = branchEvalIn_fired ? _GEN_6030 : reservedValidList2_50; // @[decode.scala 363:28 328:31]
  wire  _GEN_6680 = branchEvalIn_fired ? _GEN_6031 : reservedValidList2_51; // @[decode.scala 363:28 328:31]
  wire  _GEN_6681 = branchEvalIn_fired ? _GEN_6032 : reservedValidList2_52; // @[decode.scala 363:28 328:31]
  wire  _GEN_6682 = branchEvalIn_fired ? _GEN_6033 : reservedValidList2_53; // @[decode.scala 363:28 328:31]
  wire  _GEN_6683 = branchEvalIn_fired ? _GEN_6034 : reservedValidList2_54; // @[decode.scala 363:28 328:31]
  wire  _GEN_6684 = branchEvalIn_fired ? _GEN_6035 : reservedValidList2_55; // @[decode.scala 363:28 328:31]
  wire  _GEN_6685 = branchEvalIn_fired ? _GEN_6036 : reservedValidList2_56; // @[decode.scala 363:28 328:31]
  wire  _GEN_6686 = branchEvalIn_fired ? _GEN_6037 : reservedValidList2_57; // @[decode.scala 363:28 328:31]
  wire  _GEN_6687 = branchEvalIn_fired ? _GEN_6038 : reservedValidList2_58; // @[decode.scala 363:28 328:31]
  wire  _GEN_6688 = branchEvalIn_fired ? _GEN_6039 : reservedValidList2_59; // @[decode.scala 363:28 328:31]
  wire  _GEN_6689 = branchEvalIn_fired ? _GEN_6040 : reservedValidList2_60; // @[decode.scala 363:28 328:31]
  wire  _GEN_6690 = branchEvalIn_fired ? _GEN_6041 : reservedValidList2_61; // @[decode.scala 363:28 328:31]
  wire  _GEN_6691 = branchEvalIn_fired ? _GEN_6042 : reservedValidList2_62; // @[decode.scala 363:28 328:31]
  wire  _GEN_6692 = branchEvalIn_fired ? _GEN_6043 : reservedValidList2_63; // @[decode.scala 363:28 328:31]
  wire  _GEN_6693 = branchEvalIn_fired ? _GEN_6044 : reservedValidList3_0; // @[decode.scala 363:28 329:31]
  wire  _GEN_6694 = branchEvalIn_fired ? _GEN_6045 : reservedValidList3_1; // @[decode.scala 363:28 329:31]
  wire  _GEN_6695 = branchEvalIn_fired ? _GEN_6046 : reservedValidList3_2; // @[decode.scala 363:28 329:31]
  wire  _GEN_6696 = branchEvalIn_fired ? _GEN_6047 : reservedValidList3_3; // @[decode.scala 363:28 329:31]
  wire  _GEN_6697 = branchEvalIn_fired ? _GEN_6048 : reservedValidList3_4; // @[decode.scala 363:28 329:31]
  wire  _GEN_6698 = branchEvalIn_fired ? _GEN_6049 : reservedValidList3_5; // @[decode.scala 363:28 329:31]
  wire  _GEN_6699 = branchEvalIn_fired ? _GEN_6050 : reservedValidList3_6; // @[decode.scala 363:28 329:31]
  wire  _GEN_6700 = branchEvalIn_fired ? _GEN_6051 : reservedValidList3_7; // @[decode.scala 363:28 329:31]
  wire  _GEN_6701 = branchEvalIn_fired ? _GEN_6052 : reservedValidList3_8; // @[decode.scala 363:28 329:31]
  wire  _GEN_6702 = branchEvalIn_fired ? _GEN_6053 : reservedValidList3_9; // @[decode.scala 363:28 329:31]
  wire  _GEN_6703 = branchEvalIn_fired ? _GEN_6054 : reservedValidList3_10; // @[decode.scala 363:28 329:31]
  wire  _GEN_6704 = branchEvalIn_fired ? _GEN_6055 : reservedValidList3_11; // @[decode.scala 363:28 329:31]
  wire  _GEN_6705 = branchEvalIn_fired ? _GEN_6056 : reservedValidList3_12; // @[decode.scala 363:28 329:31]
  wire  _GEN_6706 = branchEvalIn_fired ? _GEN_6057 : reservedValidList3_13; // @[decode.scala 363:28 329:31]
  wire  _GEN_6707 = branchEvalIn_fired ? _GEN_6058 : reservedValidList3_14; // @[decode.scala 363:28 329:31]
  wire  _GEN_6708 = branchEvalIn_fired ? _GEN_6059 : reservedValidList3_15; // @[decode.scala 363:28 329:31]
  wire  _GEN_6709 = branchEvalIn_fired ? _GEN_6060 : reservedValidList3_16; // @[decode.scala 363:28 329:31]
  wire  _GEN_6710 = branchEvalIn_fired ? _GEN_6061 : reservedValidList3_17; // @[decode.scala 363:28 329:31]
  wire  _GEN_6711 = branchEvalIn_fired ? _GEN_6062 : reservedValidList3_18; // @[decode.scala 363:28 329:31]
  wire  _GEN_6712 = branchEvalIn_fired ? _GEN_6063 : reservedValidList3_19; // @[decode.scala 363:28 329:31]
  wire  _GEN_6713 = branchEvalIn_fired ? _GEN_6064 : reservedValidList3_20; // @[decode.scala 363:28 329:31]
  wire  _GEN_6714 = branchEvalIn_fired ? _GEN_6065 : reservedValidList3_21; // @[decode.scala 363:28 329:31]
  wire  _GEN_6715 = branchEvalIn_fired ? _GEN_6066 : reservedValidList3_22; // @[decode.scala 363:28 329:31]
  wire  _GEN_6716 = branchEvalIn_fired ? _GEN_6067 : reservedValidList3_23; // @[decode.scala 363:28 329:31]
  wire  _GEN_6717 = branchEvalIn_fired ? _GEN_6068 : reservedValidList3_24; // @[decode.scala 363:28 329:31]
  wire  _GEN_6718 = branchEvalIn_fired ? _GEN_6069 : reservedValidList3_25; // @[decode.scala 363:28 329:31]
  wire  _GEN_6719 = branchEvalIn_fired ? _GEN_6070 : reservedValidList3_26; // @[decode.scala 363:28 329:31]
  wire  _GEN_6720 = branchEvalIn_fired ? _GEN_6071 : reservedValidList3_27; // @[decode.scala 363:28 329:31]
  wire  _GEN_6721 = branchEvalIn_fired ? _GEN_6072 : reservedValidList3_28; // @[decode.scala 363:28 329:31]
  wire  _GEN_6722 = branchEvalIn_fired ? _GEN_6073 : reservedValidList3_29; // @[decode.scala 363:28 329:31]
  wire  _GEN_6723 = branchEvalIn_fired ? _GEN_6074 : reservedValidList3_30; // @[decode.scala 363:28 329:31]
  wire  _GEN_6724 = branchEvalIn_fired ? _GEN_6075 : reservedValidList3_31; // @[decode.scala 363:28 329:31]
  wire  _GEN_6725 = branchEvalIn_fired ? _GEN_6076 : reservedValidList3_32; // @[decode.scala 363:28 329:31]
  wire  _GEN_6726 = branchEvalIn_fired ? _GEN_6077 : reservedValidList3_33; // @[decode.scala 363:28 329:31]
  wire  _GEN_6727 = branchEvalIn_fired ? _GEN_6078 : reservedValidList3_34; // @[decode.scala 363:28 329:31]
  wire  _GEN_6728 = branchEvalIn_fired ? _GEN_6079 : reservedValidList3_35; // @[decode.scala 363:28 329:31]
  wire  _GEN_6729 = branchEvalIn_fired ? _GEN_6080 : reservedValidList3_36; // @[decode.scala 363:28 329:31]
  wire  _GEN_6730 = branchEvalIn_fired ? _GEN_6081 : reservedValidList3_37; // @[decode.scala 363:28 329:31]
  wire  _GEN_6731 = branchEvalIn_fired ? _GEN_6082 : reservedValidList3_38; // @[decode.scala 363:28 329:31]
  wire  _GEN_6732 = branchEvalIn_fired ? _GEN_6083 : reservedValidList3_39; // @[decode.scala 363:28 329:31]
  wire  _GEN_6733 = branchEvalIn_fired ? _GEN_6084 : reservedValidList3_40; // @[decode.scala 363:28 329:31]
  wire  _GEN_6734 = branchEvalIn_fired ? _GEN_6085 : reservedValidList3_41; // @[decode.scala 363:28 329:31]
  wire  _GEN_6735 = branchEvalIn_fired ? _GEN_6086 : reservedValidList3_42; // @[decode.scala 363:28 329:31]
  wire  _GEN_6736 = branchEvalIn_fired ? _GEN_6087 : reservedValidList3_43; // @[decode.scala 363:28 329:31]
  wire  _GEN_6737 = branchEvalIn_fired ? _GEN_6088 : reservedValidList3_44; // @[decode.scala 363:28 329:31]
  wire  _GEN_6738 = branchEvalIn_fired ? _GEN_6089 : reservedValidList3_45; // @[decode.scala 363:28 329:31]
  wire  _GEN_6739 = branchEvalIn_fired ? _GEN_6090 : reservedValidList3_46; // @[decode.scala 363:28 329:31]
  wire  _GEN_6740 = branchEvalIn_fired ? _GEN_6091 : reservedValidList3_47; // @[decode.scala 363:28 329:31]
  wire  _GEN_6741 = branchEvalIn_fired ? _GEN_6092 : reservedValidList3_48; // @[decode.scala 363:28 329:31]
  wire  _GEN_6742 = branchEvalIn_fired ? _GEN_6093 : reservedValidList3_49; // @[decode.scala 363:28 329:31]
  wire  _GEN_6743 = branchEvalIn_fired ? _GEN_6094 : reservedValidList3_50; // @[decode.scala 363:28 329:31]
  wire  _GEN_6744 = branchEvalIn_fired ? _GEN_6095 : reservedValidList3_51; // @[decode.scala 363:28 329:31]
  wire  _GEN_6745 = branchEvalIn_fired ? _GEN_6096 : reservedValidList3_52; // @[decode.scala 363:28 329:31]
  wire  _GEN_6746 = branchEvalIn_fired ? _GEN_6097 : reservedValidList3_53; // @[decode.scala 363:28 329:31]
  wire  _GEN_6747 = branchEvalIn_fired ? _GEN_6098 : reservedValidList3_54; // @[decode.scala 363:28 329:31]
  wire  _GEN_6748 = branchEvalIn_fired ? _GEN_6099 : reservedValidList3_55; // @[decode.scala 363:28 329:31]
  wire  _GEN_6749 = branchEvalIn_fired ? _GEN_6100 : reservedValidList3_56; // @[decode.scala 363:28 329:31]
  wire  _GEN_6750 = branchEvalIn_fired ? _GEN_6101 : reservedValidList3_57; // @[decode.scala 363:28 329:31]
  wire  _GEN_6751 = branchEvalIn_fired ? _GEN_6102 : reservedValidList3_58; // @[decode.scala 363:28 329:31]
  wire  _GEN_6752 = branchEvalIn_fired ? _GEN_6103 : reservedValidList3_59; // @[decode.scala 363:28 329:31]
  wire  _GEN_6753 = branchEvalIn_fired ? _GEN_6104 : reservedValidList3_60; // @[decode.scala 363:28 329:31]
  wire  _GEN_6754 = branchEvalIn_fired ? _GEN_6105 : reservedValidList3_61; // @[decode.scala 363:28 329:31]
  wire  _GEN_6755 = branchEvalIn_fired ? _GEN_6106 : reservedValidList3_62; // @[decode.scala 363:28 329:31]
  wire  _GEN_6756 = branchEvalIn_fired ? _GEN_6107 : reservedValidList3_63; // @[decode.scala 363:28 329:31]
  wire [4:0] _bitPosition_T_1 = ~_toExec_branchMask_T; // @[decode.scala 417:34]
  wire [2:0] _bitPosition_T_7 = _bitPosition_T_1[3] ? 3'h3 : 3'h4; // @[Mux.scala 47:70]
  wire [2:0] _bitPosition_T_8 = _bitPosition_T_1[2] ? 3'h2 : _bitPosition_T_7; // @[Mux.scala 47:70]
  wire [2:0] _bitPosition_T_9 = _bitPosition_T_1[1] ? 3'h1 : _bitPosition_T_8; // @[Mux.scala 47:70]
  wire [2:0] _bitPosition_T_10 = _bitPosition_T_1[0] ? 3'h0 : _bitPosition_T_9; // @[Mux.scala 47:70]
  wire  _T_191 = _T_442 | _T_444 | _T_441; // @[decode.scala 420:50]
  wire [1:0] bitPosition = _bitPosition_T_10[1:0];
  wire  _GEN_16095 = 2'h0 == bitPosition; // @[decode.scala 423:{44,44}]
  wire  _GEN_6757 = 2'h0 == bitPosition | _GEN_6109; // @[decode.scala 423:{44,44}]
  wire  _GEN_16096 = 2'h1 == bitPosition; // @[decode.scala 423:{44,44}]
  wire  _GEN_6758 = 2'h1 == bitPosition | _GEN_6110; // @[decode.scala 423:{44,44}]
  wire  _GEN_16097 = 2'h2 == bitPosition; // @[decode.scala 423:{44,44}]
  wire  _GEN_6759 = 2'h2 == bitPosition | _GEN_6111; // @[decode.scala 423:{44,44}]
  wire  _GEN_16098 = 2'h3 == bitPosition; // @[decode.scala 423:{44,44}]
  wire  _GEN_6760 = 2'h3 == bitPosition | _GEN_6112; // @[decode.scala 423:{44,44}]
  wire [2:0] _GEN_16099 = {{1'd0}, bitPosition}; // @[decode.scala 423:{44,44}]
  wire  _GEN_6761 = 3'h4 == _GEN_16099 | _GEN_6113; // @[decode.scala 423:{44,44}]
  wire [4:0] _GEN_6762 = _GEN_16098 ? 5'h8 : branchPCMask; // @[decode.scala 424:27 225:29 428:32]
  wire [4:0] _GEN_6763 = _GEN_16097 ? 5'h4 : _GEN_6762; // @[decode.scala 424:27 427:32]
  wire [4:0] _GEN_6764 = _GEN_16096 ? 5'h2 : _GEN_6763; // @[decode.scala 424:27 426:32]
  wire  _GEN_6798 = 6'h0 == freeRegAddr ? 1'h0 : PRFFreeList_0; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6799 = 6'h1 == freeRegAddr ? 1'h0 : PRFFreeList_1; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6800 = 6'h2 == freeRegAddr ? 1'h0 : PRFFreeList_2; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6801 = 6'h3 == freeRegAddr ? 1'h0 : PRFFreeList_3; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6802 = 6'h4 == freeRegAddr ? 1'h0 : PRFFreeList_4; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6803 = 6'h5 == freeRegAddr ? 1'h0 : PRFFreeList_5; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6804 = 6'h6 == freeRegAddr ? 1'h0 : PRFFreeList_6; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6805 = 6'h7 == freeRegAddr ? 1'h0 : PRFFreeList_7; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6806 = 6'h8 == freeRegAddr ? 1'h0 : PRFFreeList_8; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6807 = 6'h9 == freeRegAddr ? 1'h0 : PRFFreeList_9; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6808 = 6'ha == freeRegAddr ? 1'h0 : PRFFreeList_10; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6809 = 6'hb == freeRegAddr ? 1'h0 : PRFFreeList_11; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6810 = 6'hc == freeRegAddr ? 1'h0 : PRFFreeList_12; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6811 = 6'hd == freeRegAddr ? 1'h0 : PRFFreeList_13; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6812 = 6'he == freeRegAddr ? 1'h0 : PRFFreeList_14; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6813 = 6'hf == freeRegAddr ? 1'h0 : PRFFreeList_15; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6814 = 6'h10 == freeRegAddr ? 1'h0 : PRFFreeList_16; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6815 = 6'h11 == freeRegAddr ? 1'h0 : PRFFreeList_17; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6816 = 6'h12 == freeRegAddr ? 1'h0 : PRFFreeList_18; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6817 = 6'h13 == freeRegAddr ? 1'h0 : PRFFreeList_19; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6818 = 6'h14 == freeRegAddr ? 1'h0 : PRFFreeList_20; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6819 = 6'h15 == freeRegAddr ? 1'h0 : PRFFreeList_21; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6820 = 6'h16 == freeRegAddr ? 1'h0 : PRFFreeList_22; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6821 = 6'h17 == freeRegAddr ? 1'h0 : PRFFreeList_23; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6822 = 6'h18 == freeRegAddr ? 1'h0 : PRFFreeList_24; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6823 = 6'h19 == freeRegAddr ? 1'h0 : PRFFreeList_25; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6824 = 6'h1a == freeRegAddr ? 1'h0 : PRFFreeList_26; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6825 = 6'h1b == freeRegAddr ? 1'h0 : PRFFreeList_27; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6826 = 6'h1c == freeRegAddr ? 1'h0 : PRFFreeList_28; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6827 = 6'h1d == freeRegAddr ? 1'h0 : PRFFreeList_29; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6828 = 6'h1e == freeRegAddr ? 1'h0 : PRFFreeList_30; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6829 = 6'h1f == freeRegAddr ? 1'h0 : PRFFreeList_31; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6830 = 6'h20 == freeRegAddr ? 1'h0 : PRFFreeList_32; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6831 = 6'h21 == freeRegAddr ? 1'h0 : PRFFreeList_33; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6832 = 6'h22 == freeRegAddr ? 1'h0 : PRFFreeList_34; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6833 = 6'h23 == freeRegAddr ? 1'h0 : PRFFreeList_35; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6834 = 6'h24 == freeRegAddr ? 1'h0 : PRFFreeList_36; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6835 = 6'h25 == freeRegAddr ? 1'h0 : PRFFreeList_37; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6836 = 6'h26 == freeRegAddr ? 1'h0 : PRFFreeList_38; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6837 = 6'h27 == freeRegAddr ? 1'h0 : PRFFreeList_39; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6838 = 6'h28 == freeRegAddr ? 1'h0 : PRFFreeList_40; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6839 = 6'h29 == freeRegAddr ? 1'h0 : PRFFreeList_41; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6840 = 6'h2a == freeRegAddr ? 1'h0 : PRFFreeList_42; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6841 = 6'h2b == freeRegAddr ? 1'h0 : PRFFreeList_43; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6842 = 6'h2c == freeRegAddr ? 1'h0 : PRFFreeList_44; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6843 = 6'h2d == freeRegAddr ? 1'h0 : PRFFreeList_45; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6844 = 6'h2e == freeRegAddr ? 1'h0 : PRFFreeList_46; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6845 = 6'h2f == freeRegAddr ? 1'h0 : PRFFreeList_47; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6846 = 6'h30 == freeRegAddr ? 1'h0 : PRFFreeList_48; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6847 = 6'h31 == freeRegAddr ? 1'h0 : PRFFreeList_49; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6848 = 6'h32 == freeRegAddr ? 1'h0 : PRFFreeList_50; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6849 = 6'h33 == freeRegAddr ? 1'h0 : PRFFreeList_51; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6850 = 6'h34 == freeRegAddr ? 1'h0 : PRFFreeList_52; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6851 = 6'h35 == freeRegAddr ? 1'h0 : PRFFreeList_53; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6852 = 6'h36 == freeRegAddr ? 1'h0 : PRFFreeList_54; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6853 = 6'h37 == freeRegAddr ? 1'h0 : PRFFreeList_55; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6854 = 6'h38 == freeRegAddr ? 1'h0 : PRFFreeList_56; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6855 = 6'h39 == freeRegAddr ? 1'h0 : PRFFreeList_57; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6856 = 6'h3a == freeRegAddr ? 1'h0 : PRFFreeList_58; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6857 = 6'h3b == freeRegAddr ? 1'h0 : PRFFreeList_59; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6858 = 6'h3c == freeRegAddr ? 1'h0 : PRFFreeList_60; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6859 = 6'h3d == freeRegAddr ? 1'h0 : PRFFreeList_61; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6860 = 6'h3e == freeRegAddr ? 1'h0 : PRFFreeList_62; // @[decode.scala 434:30 438:{45,45}]
  wire  _GEN_6862 = 6'h0 == freeRegAddr ? 1'h0 : PRFValidList_0; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6863 = 6'h1 == freeRegAddr ? 1'h0 : PRFValidList_1; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6864 = 6'h2 == freeRegAddr ? 1'h0 : PRFValidList_2; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6865 = 6'h3 == freeRegAddr ? 1'h0 : PRFValidList_3; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6866 = 6'h4 == freeRegAddr ? 1'h0 : PRFValidList_4; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6867 = 6'h5 == freeRegAddr ? 1'h0 : PRFValidList_5; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6868 = 6'h6 == freeRegAddr ? 1'h0 : PRFValidList_6; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6869 = 6'h7 == freeRegAddr ? 1'h0 : PRFValidList_7; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6870 = 6'h8 == freeRegAddr ? 1'h0 : PRFValidList_8; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6871 = 6'h9 == freeRegAddr ? 1'h0 : PRFValidList_9; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6872 = 6'ha == freeRegAddr ? 1'h0 : PRFValidList_10; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6873 = 6'hb == freeRegAddr ? 1'h0 : PRFValidList_11; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6874 = 6'hc == freeRegAddr ? 1'h0 : PRFValidList_12; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6875 = 6'hd == freeRegAddr ? 1'h0 : PRFValidList_13; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6876 = 6'he == freeRegAddr ? 1'h0 : PRFValidList_14; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6877 = 6'hf == freeRegAddr ? 1'h0 : PRFValidList_15; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6878 = 6'h10 == freeRegAddr ? 1'h0 : PRFValidList_16; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6879 = 6'h11 == freeRegAddr ? 1'h0 : PRFValidList_17; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6880 = 6'h12 == freeRegAddr ? 1'h0 : PRFValidList_18; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6881 = 6'h13 == freeRegAddr ? 1'h0 : PRFValidList_19; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6882 = 6'h14 == freeRegAddr ? 1'h0 : PRFValidList_20; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6883 = 6'h15 == freeRegAddr ? 1'h0 : PRFValidList_21; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6884 = 6'h16 == freeRegAddr ? 1'h0 : PRFValidList_22; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6885 = 6'h17 == freeRegAddr ? 1'h0 : PRFValidList_23; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6886 = 6'h18 == freeRegAddr ? 1'h0 : PRFValidList_24; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6887 = 6'h19 == freeRegAddr ? 1'h0 : PRFValidList_25; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6888 = 6'h1a == freeRegAddr ? 1'h0 : PRFValidList_26; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6889 = 6'h1b == freeRegAddr ? 1'h0 : PRFValidList_27; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6890 = 6'h1c == freeRegAddr ? 1'h0 : PRFValidList_28; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6891 = 6'h1d == freeRegAddr ? 1'h0 : PRFValidList_29; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6892 = 6'h1e == freeRegAddr ? 1'h0 : PRFValidList_30; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6893 = 6'h1f == freeRegAddr ? 1'h0 : PRFValidList_31; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6894 = 6'h20 == freeRegAddr ? 1'h0 : PRFValidList_32; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6895 = 6'h21 == freeRegAddr ? 1'h0 : PRFValidList_33; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6896 = 6'h22 == freeRegAddr ? 1'h0 : PRFValidList_34; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6897 = 6'h23 == freeRegAddr ? 1'h0 : PRFValidList_35; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6898 = 6'h24 == freeRegAddr ? 1'h0 : PRFValidList_36; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6899 = 6'h25 == freeRegAddr ? 1'h0 : PRFValidList_37; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6900 = 6'h26 == freeRegAddr ? 1'h0 : PRFValidList_38; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6901 = 6'h27 == freeRegAddr ? 1'h0 : PRFValidList_39; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6902 = 6'h28 == freeRegAddr ? 1'h0 : PRFValidList_40; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6903 = 6'h29 == freeRegAddr ? 1'h0 : PRFValidList_41; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6904 = 6'h2a == freeRegAddr ? 1'h0 : PRFValidList_42; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6905 = 6'h2b == freeRegAddr ? 1'h0 : PRFValidList_43; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6906 = 6'h2c == freeRegAddr ? 1'h0 : PRFValidList_44; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6907 = 6'h2d == freeRegAddr ? 1'h0 : PRFValidList_45; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6908 = 6'h2e == freeRegAddr ? 1'h0 : PRFValidList_46; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6909 = 6'h2f == freeRegAddr ? 1'h0 : PRFValidList_47; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6910 = 6'h30 == freeRegAddr ? 1'h0 : PRFValidList_48; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6911 = 6'h31 == freeRegAddr ? 1'h0 : PRFValidList_49; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6912 = 6'h32 == freeRegAddr ? 1'h0 : PRFValidList_50; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6913 = 6'h33 == freeRegAddr ? 1'h0 : PRFValidList_51; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6914 = 6'h34 == freeRegAddr ? 1'h0 : PRFValidList_52; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6915 = 6'h35 == freeRegAddr ? 1'h0 : PRFValidList_53; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6916 = 6'h36 == freeRegAddr ? 1'h0 : PRFValidList_54; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6917 = 6'h37 == freeRegAddr ? 1'h0 : PRFValidList_55; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6918 = 6'h38 == freeRegAddr ? 1'h0 : PRFValidList_56; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6919 = 6'h39 == freeRegAddr ? 1'h0 : PRFValidList_57; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6920 = 6'h3a == freeRegAddr ? 1'h0 : PRFValidList_58; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6921 = 6'h3b == freeRegAddr ? 1'h0 : PRFValidList_59; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6922 = 6'h3c == freeRegAddr ? 1'h0 : PRFValidList_60; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6923 = 6'h3d == freeRegAddr ? 1'h0 : PRFValidList_61; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6924 = 6'h3e == freeRegAddr ? 1'h0 : PRFValidList_62; // @[decode.scala 435:30 439:{45,45}]
  wire  _GEN_6925 = 6'h3f == freeRegAddr ? 1'h0 : PRFValidList_63; // @[decode.scala 435:30 439:{45,45}]
  wire [5:0] _GEN_6926 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_850 : frontEndRegMap_0; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6927 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_851 : frontEndRegMap_1; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6928 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_852 : frontEndRegMap_2; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6929 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_853 : frontEndRegMap_3; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6930 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_854 : frontEndRegMap_4; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6931 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_855 : frontEndRegMap_5; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6932 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_856 : frontEndRegMap_6; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6933 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_857 : frontEndRegMap_7; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6934 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_858 : frontEndRegMap_8; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6935 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_859 : frontEndRegMap_9; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6936 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_860 : frontEndRegMap_10; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6937 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_861 : frontEndRegMap_11; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6938 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_862 : frontEndRegMap_12; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6939 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_863 : frontEndRegMap_13; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6940 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_864 : frontEndRegMap_14; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6941 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_865 : frontEndRegMap_15; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6942 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_866 : frontEndRegMap_16; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6943 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_867 : frontEndRegMap_17; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6944 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_868 : frontEndRegMap_18; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6945 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_869 : frontEndRegMap_19; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6946 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_870 : frontEndRegMap_20; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6947 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_871 : frontEndRegMap_21; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6948 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_872 : frontEndRegMap_22; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6949 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_873 : frontEndRegMap_23; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6950 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_874 : frontEndRegMap_24; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6951 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_875 : frontEndRegMap_25; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6952 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_876 : frontEndRegMap_26; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6953 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_877 : frontEndRegMap_27; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6954 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_878 : frontEndRegMap_28; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6955 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_879 : frontEndRegMap_29; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6956 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_880 : frontEndRegMap_30; // @[decode.scala 433:30 436:44]
  wire [5:0] _GEN_6957 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_881 : frontEndRegMap_31; // @[decode.scala 433:30 436:44]
  wire  _GEN_6958 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6798 : PRFFreeList_0; // @[decode.scala 434:30 436:44]
  wire  _GEN_6959 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6799 : PRFFreeList_1; // @[decode.scala 434:30 436:44]
  wire  _GEN_6960 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6800 : PRFFreeList_2; // @[decode.scala 434:30 436:44]
  wire  _GEN_6961 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6801 : PRFFreeList_3; // @[decode.scala 434:30 436:44]
  wire  _GEN_6962 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6802 : PRFFreeList_4; // @[decode.scala 434:30 436:44]
  wire  _GEN_6963 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6803 : PRFFreeList_5; // @[decode.scala 434:30 436:44]
  wire  _GEN_6964 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6804 : PRFFreeList_6; // @[decode.scala 434:30 436:44]
  wire  _GEN_6965 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6805 : PRFFreeList_7; // @[decode.scala 434:30 436:44]
  wire  _GEN_6966 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6806 : PRFFreeList_8; // @[decode.scala 434:30 436:44]
  wire  _GEN_6967 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6807 : PRFFreeList_9; // @[decode.scala 434:30 436:44]
  wire  _GEN_6968 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6808 : PRFFreeList_10; // @[decode.scala 434:30 436:44]
  wire  _GEN_6969 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6809 : PRFFreeList_11; // @[decode.scala 434:30 436:44]
  wire  _GEN_6970 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6810 : PRFFreeList_12; // @[decode.scala 434:30 436:44]
  wire  _GEN_6971 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6811 : PRFFreeList_13; // @[decode.scala 434:30 436:44]
  wire  _GEN_6972 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6812 : PRFFreeList_14; // @[decode.scala 434:30 436:44]
  wire  _GEN_6973 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6813 : PRFFreeList_15; // @[decode.scala 434:30 436:44]
  wire  _GEN_6974 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6814 : PRFFreeList_16; // @[decode.scala 434:30 436:44]
  wire  _GEN_6975 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6815 : PRFFreeList_17; // @[decode.scala 434:30 436:44]
  wire  _GEN_6976 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6816 : PRFFreeList_18; // @[decode.scala 434:30 436:44]
  wire  _GEN_6977 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6817 : PRFFreeList_19; // @[decode.scala 434:30 436:44]
  wire  _GEN_6978 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6818 : PRFFreeList_20; // @[decode.scala 434:30 436:44]
  wire  _GEN_6979 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6819 : PRFFreeList_21; // @[decode.scala 434:30 436:44]
  wire  _GEN_6980 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6820 : PRFFreeList_22; // @[decode.scala 434:30 436:44]
  wire  _GEN_6981 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6821 : PRFFreeList_23; // @[decode.scala 434:30 436:44]
  wire  _GEN_6982 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6822 : PRFFreeList_24; // @[decode.scala 434:30 436:44]
  wire  _GEN_6983 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6823 : PRFFreeList_25; // @[decode.scala 434:30 436:44]
  wire  _GEN_6984 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6824 : PRFFreeList_26; // @[decode.scala 434:30 436:44]
  wire  _GEN_6985 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6825 : PRFFreeList_27; // @[decode.scala 434:30 436:44]
  wire  _GEN_6986 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6826 : PRFFreeList_28; // @[decode.scala 434:30 436:44]
  wire  _GEN_6987 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6827 : PRFFreeList_29; // @[decode.scala 434:30 436:44]
  wire  _GEN_6988 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6828 : PRFFreeList_30; // @[decode.scala 434:30 436:44]
  wire  _GEN_6989 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6829 : PRFFreeList_31; // @[decode.scala 434:30 436:44]
  wire  _GEN_6990 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6830 : PRFFreeList_32; // @[decode.scala 434:30 436:44]
  wire  _GEN_6991 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6831 : PRFFreeList_33; // @[decode.scala 434:30 436:44]
  wire  _GEN_6992 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6832 : PRFFreeList_34; // @[decode.scala 434:30 436:44]
  wire  _GEN_6993 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6833 : PRFFreeList_35; // @[decode.scala 434:30 436:44]
  wire  _GEN_6994 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6834 : PRFFreeList_36; // @[decode.scala 434:30 436:44]
  wire  _GEN_6995 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6835 : PRFFreeList_37; // @[decode.scala 434:30 436:44]
  wire  _GEN_6996 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6836 : PRFFreeList_38; // @[decode.scala 434:30 436:44]
  wire  _GEN_6997 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6837 : PRFFreeList_39; // @[decode.scala 434:30 436:44]
  wire  _GEN_6998 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6838 : PRFFreeList_40; // @[decode.scala 434:30 436:44]
  wire  _GEN_6999 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6839 : PRFFreeList_41; // @[decode.scala 434:30 436:44]
  wire  _GEN_7000 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6840 : PRFFreeList_42; // @[decode.scala 434:30 436:44]
  wire  _GEN_7001 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6841 : PRFFreeList_43; // @[decode.scala 434:30 436:44]
  wire  _GEN_7002 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6842 : PRFFreeList_44; // @[decode.scala 434:30 436:44]
  wire  _GEN_7003 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6843 : PRFFreeList_45; // @[decode.scala 434:30 436:44]
  wire  _GEN_7004 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6844 : PRFFreeList_46; // @[decode.scala 434:30 436:44]
  wire  _GEN_7005 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6845 : PRFFreeList_47; // @[decode.scala 434:30 436:44]
  wire  _GEN_7006 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6846 : PRFFreeList_48; // @[decode.scala 434:30 436:44]
  wire  _GEN_7007 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6847 : PRFFreeList_49; // @[decode.scala 434:30 436:44]
  wire  _GEN_7008 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6848 : PRFFreeList_50; // @[decode.scala 434:30 436:44]
  wire  _GEN_7009 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6849 : PRFFreeList_51; // @[decode.scala 434:30 436:44]
  wire  _GEN_7010 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6850 : PRFFreeList_52; // @[decode.scala 434:30 436:44]
  wire  _GEN_7011 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6851 : PRFFreeList_53; // @[decode.scala 434:30 436:44]
  wire  _GEN_7012 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6852 : PRFFreeList_54; // @[decode.scala 434:30 436:44]
  wire  _GEN_7013 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6853 : PRFFreeList_55; // @[decode.scala 434:30 436:44]
  wire  _GEN_7014 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6854 : PRFFreeList_56; // @[decode.scala 434:30 436:44]
  wire  _GEN_7015 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6855 : PRFFreeList_57; // @[decode.scala 434:30 436:44]
  wire  _GEN_7016 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6856 : PRFFreeList_58; // @[decode.scala 434:30 436:44]
  wire  _GEN_7017 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6857 : PRFFreeList_59; // @[decode.scala 434:30 436:44]
  wire  _GEN_7018 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6858 : PRFFreeList_60; // @[decode.scala 434:30 436:44]
  wire  _GEN_7019 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6859 : PRFFreeList_61; // @[decode.scala 434:30 436:44]
  wire  _GEN_7020 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6860 : PRFFreeList_62; // @[decode.scala 434:30 436:44]
  wire  _GEN_7022 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6862 : PRFValidList_0; // @[decode.scala 435:30 436:44]
  wire  _GEN_7023 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6863 : PRFValidList_1; // @[decode.scala 435:30 436:44]
  wire  _GEN_7024 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6864 : PRFValidList_2; // @[decode.scala 435:30 436:44]
  wire  _GEN_7025 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6865 : PRFValidList_3; // @[decode.scala 435:30 436:44]
  wire  _GEN_7026 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6866 : PRFValidList_4; // @[decode.scala 435:30 436:44]
  wire  _GEN_7027 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6867 : PRFValidList_5; // @[decode.scala 435:30 436:44]
  wire  _GEN_7028 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6868 : PRFValidList_6; // @[decode.scala 435:30 436:44]
  wire  _GEN_7029 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6869 : PRFValidList_7; // @[decode.scala 435:30 436:44]
  wire  _GEN_7030 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6870 : PRFValidList_8; // @[decode.scala 435:30 436:44]
  wire  _GEN_7031 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6871 : PRFValidList_9; // @[decode.scala 435:30 436:44]
  wire  _GEN_7032 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6872 : PRFValidList_10; // @[decode.scala 435:30 436:44]
  wire  _GEN_7033 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6873 : PRFValidList_11; // @[decode.scala 435:30 436:44]
  wire  _GEN_7034 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6874 : PRFValidList_12; // @[decode.scala 435:30 436:44]
  wire  _GEN_7035 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6875 : PRFValidList_13; // @[decode.scala 435:30 436:44]
  wire  _GEN_7036 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6876 : PRFValidList_14; // @[decode.scala 435:30 436:44]
  wire  _GEN_7037 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6877 : PRFValidList_15; // @[decode.scala 435:30 436:44]
  wire  _GEN_7038 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6878 : PRFValidList_16; // @[decode.scala 435:30 436:44]
  wire  _GEN_7039 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6879 : PRFValidList_17; // @[decode.scala 435:30 436:44]
  wire  _GEN_7040 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6880 : PRFValidList_18; // @[decode.scala 435:30 436:44]
  wire  _GEN_7041 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6881 : PRFValidList_19; // @[decode.scala 435:30 436:44]
  wire  _GEN_7042 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6882 : PRFValidList_20; // @[decode.scala 435:30 436:44]
  wire  _GEN_7043 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6883 : PRFValidList_21; // @[decode.scala 435:30 436:44]
  wire  _GEN_7044 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6884 : PRFValidList_22; // @[decode.scala 435:30 436:44]
  wire  _GEN_7045 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6885 : PRFValidList_23; // @[decode.scala 435:30 436:44]
  wire  _GEN_7046 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6886 : PRFValidList_24; // @[decode.scala 435:30 436:44]
  wire  _GEN_7047 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6887 : PRFValidList_25; // @[decode.scala 435:30 436:44]
  wire  _GEN_7048 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6888 : PRFValidList_26; // @[decode.scala 435:30 436:44]
  wire  _GEN_7049 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6889 : PRFValidList_27; // @[decode.scala 435:30 436:44]
  wire  _GEN_7050 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6890 : PRFValidList_28; // @[decode.scala 435:30 436:44]
  wire  _GEN_7051 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6891 : PRFValidList_29; // @[decode.scala 435:30 436:44]
  wire  _GEN_7052 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6892 : PRFValidList_30; // @[decode.scala 435:30 436:44]
  wire  _GEN_7053 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6893 : PRFValidList_31; // @[decode.scala 435:30 436:44]
  wire  _GEN_7054 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6894 : PRFValidList_32; // @[decode.scala 435:30 436:44]
  wire  _GEN_7055 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6895 : PRFValidList_33; // @[decode.scala 435:30 436:44]
  wire  _GEN_7056 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6896 : PRFValidList_34; // @[decode.scala 435:30 436:44]
  wire  _GEN_7057 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6897 : PRFValidList_35; // @[decode.scala 435:30 436:44]
  wire  _GEN_7058 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6898 : PRFValidList_36; // @[decode.scala 435:30 436:44]
  wire  _GEN_7059 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6899 : PRFValidList_37; // @[decode.scala 435:30 436:44]
  wire  _GEN_7060 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6900 : PRFValidList_38; // @[decode.scala 435:30 436:44]
  wire  _GEN_7061 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6901 : PRFValidList_39; // @[decode.scala 435:30 436:44]
  wire  _GEN_7062 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6902 : PRFValidList_40; // @[decode.scala 435:30 436:44]
  wire  _GEN_7063 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6903 : PRFValidList_41; // @[decode.scala 435:30 436:44]
  wire  _GEN_7064 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6904 : PRFValidList_42; // @[decode.scala 435:30 436:44]
  wire  _GEN_7065 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6905 : PRFValidList_43; // @[decode.scala 435:30 436:44]
  wire  _GEN_7066 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6906 : PRFValidList_44; // @[decode.scala 435:30 436:44]
  wire  _GEN_7067 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6907 : PRFValidList_45; // @[decode.scala 435:30 436:44]
  wire  _GEN_7068 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6908 : PRFValidList_46; // @[decode.scala 435:30 436:44]
  wire  _GEN_7069 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6909 : PRFValidList_47; // @[decode.scala 435:30 436:44]
  wire  _GEN_7070 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6910 : PRFValidList_48; // @[decode.scala 435:30 436:44]
  wire  _GEN_7071 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6911 : PRFValidList_49; // @[decode.scala 435:30 436:44]
  wire  _GEN_7072 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6912 : PRFValidList_50; // @[decode.scala 435:30 436:44]
  wire  _GEN_7073 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6913 : PRFValidList_51; // @[decode.scala 435:30 436:44]
  wire  _GEN_7074 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6914 : PRFValidList_52; // @[decode.scala 435:30 436:44]
  wire  _GEN_7075 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6915 : PRFValidList_53; // @[decode.scala 435:30 436:44]
  wire  _GEN_7076 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6916 : PRFValidList_54; // @[decode.scala 435:30 436:44]
  wire  _GEN_7077 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6917 : PRFValidList_55; // @[decode.scala 435:30 436:44]
  wire  _GEN_7078 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6918 : PRFValidList_56; // @[decode.scala 435:30 436:44]
  wire  _GEN_7079 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6919 : PRFValidList_57; // @[decode.scala 435:30 436:44]
  wire  _GEN_7080 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6920 : PRFValidList_58; // @[decode.scala 435:30 436:44]
  wire  _GEN_7081 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6921 : PRFValidList_59; // @[decode.scala 435:30 436:44]
  wire  _GEN_7082 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6922 : PRFValidList_60; // @[decode.scala 435:30 436:44]
  wire  _GEN_7083 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6923 : PRFValidList_61; // @[decode.scala 435:30 436:44]
  wire  _GEN_7084 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6924 : PRFValidList_62; // @[decode.scala 435:30 436:44]
  wire  _GEN_7085 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_6925 : PRFValidList_63; // @[decode.scala 435:30 436:44]
  wire [5:0] _GEN_8046 = 3'h3 == branchTracker ? _GEN_6926 : reservedRegMap4_0; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8047 = 3'h3 == branchTracker ? _GEN_6927 : reservedRegMap4_1; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8048 = 3'h3 == branchTracker ? _GEN_6928 : reservedRegMap4_2; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8049 = 3'h3 == branchTracker ? _GEN_6929 : reservedRegMap4_3; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8050 = 3'h3 == branchTracker ? _GEN_6930 : reservedRegMap4_4; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8051 = 3'h3 == branchTracker ? _GEN_6931 : reservedRegMap4_5; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8052 = 3'h3 == branchTracker ? _GEN_6932 : reservedRegMap4_6; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8053 = 3'h3 == branchTracker ? _GEN_6933 : reservedRegMap4_7; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8054 = 3'h3 == branchTracker ? _GEN_6934 : reservedRegMap4_8; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8055 = 3'h3 == branchTracker ? _GEN_6935 : reservedRegMap4_9; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8056 = 3'h3 == branchTracker ? _GEN_6936 : reservedRegMap4_10; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8057 = 3'h3 == branchTracker ? _GEN_6937 : reservedRegMap4_11; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8058 = 3'h3 == branchTracker ? _GEN_6938 : reservedRegMap4_12; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8059 = 3'h3 == branchTracker ? _GEN_6939 : reservedRegMap4_13; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8060 = 3'h3 == branchTracker ? _GEN_6940 : reservedRegMap4_14; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8061 = 3'h3 == branchTracker ? _GEN_6941 : reservedRegMap4_15; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8062 = 3'h3 == branchTracker ? _GEN_6942 : reservedRegMap4_16; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8063 = 3'h3 == branchTracker ? _GEN_6943 : reservedRegMap4_17; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8064 = 3'h3 == branchTracker ? _GEN_6944 : reservedRegMap4_18; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8065 = 3'h3 == branchTracker ? _GEN_6945 : reservedRegMap4_19; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8066 = 3'h3 == branchTracker ? _GEN_6946 : reservedRegMap4_20; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8067 = 3'h3 == branchTracker ? _GEN_6947 : reservedRegMap4_21; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8068 = 3'h3 == branchTracker ? _GEN_6948 : reservedRegMap4_22; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8069 = 3'h3 == branchTracker ? _GEN_6949 : reservedRegMap4_23; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8070 = 3'h3 == branchTracker ? _GEN_6950 : reservedRegMap4_24; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8071 = 3'h3 == branchTracker ? _GEN_6951 : reservedRegMap4_25; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8072 = 3'h3 == branchTracker ? _GEN_6952 : reservedRegMap4_26; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8073 = 3'h3 == branchTracker ? _GEN_6953 : reservedRegMap4_27; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8074 = 3'h3 == branchTracker ? _GEN_6954 : reservedRegMap4_28; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8075 = 3'h3 == branchTracker ? _GEN_6955 : reservedRegMap4_29; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8076 = 3'h3 == branchTracker ? _GEN_6956 : reservedRegMap4_30; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8077 = 3'h3 == branchTracker ? _GEN_6957 : reservedRegMap4_31; // @[decode.scala 320:28 431:29]
  wire  _GEN_8078 = 3'h3 == branchTracker ? _GEN_6958 : reservedFreeList4_0; // @[decode.scala 431:29 325:30]
  wire  _GEN_8079 = 3'h3 == branchTracker ? _GEN_6959 : reservedFreeList4_1; // @[decode.scala 431:29 325:30]
  wire  _GEN_8080 = 3'h3 == branchTracker ? _GEN_6960 : reservedFreeList4_2; // @[decode.scala 431:29 325:30]
  wire  _GEN_8081 = 3'h3 == branchTracker ? _GEN_6961 : reservedFreeList4_3; // @[decode.scala 431:29 325:30]
  wire  _GEN_8082 = 3'h3 == branchTracker ? _GEN_6962 : reservedFreeList4_4; // @[decode.scala 431:29 325:30]
  wire  _GEN_8083 = 3'h3 == branchTracker ? _GEN_6963 : reservedFreeList4_5; // @[decode.scala 431:29 325:30]
  wire  _GEN_8084 = 3'h3 == branchTracker ? _GEN_6964 : reservedFreeList4_6; // @[decode.scala 431:29 325:30]
  wire  _GEN_8085 = 3'h3 == branchTracker ? _GEN_6965 : reservedFreeList4_7; // @[decode.scala 431:29 325:30]
  wire  _GEN_8086 = 3'h3 == branchTracker ? _GEN_6966 : reservedFreeList4_8; // @[decode.scala 431:29 325:30]
  wire  _GEN_8087 = 3'h3 == branchTracker ? _GEN_6967 : reservedFreeList4_9; // @[decode.scala 431:29 325:30]
  wire  _GEN_8088 = 3'h3 == branchTracker ? _GEN_6968 : reservedFreeList4_10; // @[decode.scala 431:29 325:30]
  wire  _GEN_8089 = 3'h3 == branchTracker ? _GEN_6969 : reservedFreeList4_11; // @[decode.scala 431:29 325:30]
  wire  _GEN_8090 = 3'h3 == branchTracker ? _GEN_6970 : reservedFreeList4_12; // @[decode.scala 431:29 325:30]
  wire  _GEN_8091 = 3'h3 == branchTracker ? _GEN_6971 : reservedFreeList4_13; // @[decode.scala 431:29 325:30]
  wire  _GEN_8092 = 3'h3 == branchTracker ? _GEN_6972 : reservedFreeList4_14; // @[decode.scala 431:29 325:30]
  wire  _GEN_8093 = 3'h3 == branchTracker ? _GEN_6973 : reservedFreeList4_15; // @[decode.scala 431:29 325:30]
  wire  _GEN_8094 = 3'h3 == branchTracker ? _GEN_6974 : reservedFreeList4_16; // @[decode.scala 431:29 325:30]
  wire  _GEN_8095 = 3'h3 == branchTracker ? _GEN_6975 : reservedFreeList4_17; // @[decode.scala 431:29 325:30]
  wire  _GEN_8096 = 3'h3 == branchTracker ? _GEN_6976 : reservedFreeList4_18; // @[decode.scala 431:29 325:30]
  wire  _GEN_8097 = 3'h3 == branchTracker ? _GEN_6977 : reservedFreeList4_19; // @[decode.scala 431:29 325:30]
  wire  _GEN_8098 = 3'h3 == branchTracker ? _GEN_6978 : reservedFreeList4_20; // @[decode.scala 431:29 325:30]
  wire  _GEN_8099 = 3'h3 == branchTracker ? _GEN_6979 : reservedFreeList4_21; // @[decode.scala 431:29 325:30]
  wire  _GEN_8100 = 3'h3 == branchTracker ? _GEN_6980 : reservedFreeList4_22; // @[decode.scala 431:29 325:30]
  wire  _GEN_8101 = 3'h3 == branchTracker ? _GEN_6981 : reservedFreeList4_23; // @[decode.scala 431:29 325:30]
  wire  _GEN_8102 = 3'h3 == branchTracker ? _GEN_6982 : reservedFreeList4_24; // @[decode.scala 431:29 325:30]
  wire  _GEN_8103 = 3'h3 == branchTracker ? _GEN_6983 : reservedFreeList4_25; // @[decode.scala 431:29 325:30]
  wire  _GEN_8104 = 3'h3 == branchTracker ? _GEN_6984 : reservedFreeList4_26; // @[decode.scala 431:29 325:30]
  wire  _GEN_8105 = 3'h3 == branchTracker ? _GEN_6985 : reservedFreeList4_27; // @[decode.scala 431:29 325:30]
  wire  _GEN_8106 = 3'h3 == branchTracker ? _GEN_6986 : reservedFreeList4_28; // @[decode.scala 431:29 325:30]
  wire  _GEN_8107 = 3'h3 == branchTracker ? _GEN_6987 : reservedFreeList4_29; // @[decode.scala 431:29 325:30]
  wire  _GEN_8108 = 3'h3 == branchTracker ? _GEN_6988 : reservedFreeList4_30; // @[decode.scala 431:29 325:30]
  wire  _GEN_8109 = 3'h3 == branchTracker ? _GEN_6989 : reservedFreeList4_31; // @[decode.scala 431:29 325:30]
  wire  _GEN_8110 = 3'h3 == branchTracker ? _GEN_6990 : reservedFreeList4_32; // @[decode.scala 431:29 325:30]
  wire  _GEN_8111 = 3'h3 == branchTracker ? _GEN_6991 : reservedFreeList4_33; // @[decode.scala 431:29 325:30]
  wire  _GEN_8112 = 3'h3 == branchTracker ? _GEN_6992 : reservedFreeList4_34; // @[decode.scala 431:29 325:30]
  wire  _GEN_8113 = 3'h3 == branchTracker ? _GEN_6993 : reservedFreeList4_35; // @[decode.scala 431:29 325:30]
  wire  _GEN_8114 = 3'h3 == branchTracker ? _GEN_6994 : reservedFreeList4_36; // @[decode.scala 431:29 325:30]
  wire  _GEN_8115 = 3'h3 == branchTracker ? _GEN_6995 : reservedFreeList4_37; // @[decode.scala 431:29 325:30]
  wire  _GEN_8116 = 3'h3 == branchTracker ? _GEN_6996 : reservedFreeList4_38; // @[decode.scala 431:29 325:30]
  wire  _GEN_8117 = 3'h3 == branchTracker ? _GEN_6997 : reservedFreeList4_39; // @[decode.scala 431:29 325:30]
  wire  _GEN_8118 = 3'h3 == branchTracker ? _GEN_6998 : reservedFreeList4_40; // @[decode.scala 431:29 325:30]
  wire  _GEN_8119 = 3'h3 == branchTracker ? _GEN_6999 : reservedFreeList4_41; // @[decode.scala 431:29 325:30]
  wire  _GEN_8120 = 3'h3 == branchTracker ? _GEN_7000 : reservedFreeList4_42; // @[decode.scala 431:29 325:30]
  wire  _GEN_8121 = 3'h3 == branchTracker ? _GEN_7001 : reservedFreeList4_43; // @[decode.scala 431:29 325:30]
  wire  _GEN_8122 = 3'h3 == branchTracker ? _GEN_7002 : reservedFreeList4_44; // @[decode.scala 431:29 325:30]
  wire  _GEN_8123 = 3'h3 == branchTracker ? _GEN_7003 : reservedFreeList4_45; // @[decode.scala 431:29 325:30]
  wire  _GEN_8124 = 3'h3 == branchTracker ? _GEN_7004 : reservedFreeList4_46; // @[decode.scala 431:29 325:30]
  wire  _GEN_8125 = 3'h3 == branchTracker ? _GEN_7005 : reservedFreeList4_47; // @[decode.scala 431:29 325:30]
  wire  _GEN_8126 = 3'h3 == branchTracker ? _GEN_7006 : reservedFreeList4_48; // @[decode.scala 431:29 325:30]
  wire  _GEN_8127 = 3'h3 == branchTracker ? _GEN_7007 : reservedFreeList4_49; // @[decode.scala 431:29 325:30]
  wire  _GEN_8128 = 3'h3 == branchTracker ? _GEN_7008 : reservedFreeList4_50; // @[decode.scala 431:29 325:30]
  wire  _GEN_8129 = 3'h3 == branchTracker ? _GEN_7009 : reservedFreeList4_51; // @[decode.scala 431:29 325:30]
  wire  _GEN_8130 = 3'h3 == branchTracker ? _GEN_7010 : reservedFreeList4_52; // @[decode.scala 431:29 325:30]
  wire  _GEN_8131 = 3'h3 == branchTracker ? _GEN_7011 : reservedFreeList4_53; // @[decode.scala 431:29 325:30]
  wire  _GEN_8132 = 3'h3 == branchTracker ? _GEN_7012 : reservedFreeList4_54; // @[decode.scala 431:29 325:30]
  wire  _GEN_8133 = 3'h3 == branchTracker ? _GEN_7013 : reservedFreeList4_55; // @[decode.scala 431:29 325:30]
  wire  _GEN_8134 = 3'h3 == branchTracker ? _GEN_7014 : reservedFreeList4_56; // @[decode.scala 431:29 325:30]
  wire  _GEN_8135 = 3'h3 == branchTracker ? _GEN_7015 : reservedFreeList4_57; // @[decode.scala 431:29 325:30]
  wire  _GEN_8136 = 3'h3 == branchTracker ? _GEN_7016 : reservedFreeList4_58; // @[decode.scala 431:29 325:30]
  wire  _GEN_8137 = 3'h3 == branchTracker ? _GEN_7017 : reservedFreeList4_59; // @[decode.scala 431:29 325:30]
  wire  _GEN_8138 = 3'h3 == branchTracker ? _GEN_7018 : reservedFreeList4_60; // @[decode.scala 431:29 325:30]
  wire  _GEN_8139 = 3'h3 == branchTracker ? _GEN_7019 : reservedFreeList4_61; // @[decode.scala 431:29 325:30]
  wire  _GEN_8140 = 3'h3 == branchTracker ? _GEN_7020 : reservedFreeList4_62; // @[decode.scala 431:29 325:30]
  wire  _GEN_8142 = 3'h3 == branchTracker ? _GEN_7022 : reservedValidList4_0; // @[decode.scala 431:29 330:31]
  wire  _GEN_8143 = 3'h3 == branchTracker ? _GEN_7023 : reservedValidList4_1; // @[decode.scala 431:29 330:31]
  wire  _GEN_8144 = 3'h3 == branchTracker ? _GEN_7024 : reservedValidList4_2; // @[decode.scala 431:29 330:31]
  wire  _GEN_8145 = 3'h3 == branchTracker ? _GEN_7025 : reservedValidList4_3; // @[decode.scala 431:29 330:31]
  wire  _GEN_8146 = 3'h3 == branchTracker ? _GEN_7026 : reservedValidList4_4; // @[decode.scala 431:29 330:31]
  wire  _GEN_8147 = 3'h3 == branchTracker ? _GEN_7027 : reservedValidList4_5; // @[decode.scala 431:29 330:31]
  wire  _GEN_8148 = 3'h3 == branchTracker ? _GEN_7028 : reservedValidList4_6; // @[decode.scala 431:29 330:31]
  wire  _GEN_8149 = 3'h3 == branchTracker ? _GEN_7029 : reservedValidList4_7; // @[decode.scala 431:29 330:31]
  wire  _GEN_8150 = 3'h3 == branchTracker ? _GEN_7030 : reservedValidList4_8; // @[decode.scala 431:29 330:31]
  wire  _GEN_8151 = 3'h3 == branchTracker ? _GEN_7031 : reservedValidList4_9; // @[decode.scala 431:29 330:31]
  wire  _GEN_8152 = 3'h3 == branchTracker ? _GEN_7032 : reservedValidList4_10; // @[decode.scala 431:29 330:31]
  wire  _GEN_8153 = 3'h3 == branchTracker ? _GEN_7033 : reservedValidList4_11; // @[decode.scala 431:29 330:31]
  wire  _GEN_8154 = 3'h3 == branchTracker ? _GEN_7034 : reservedValidList4_12; // @[decode.scala 431:29 330:31]
  wire  _GEN_8155 = 3'h3 == branchTracker ? _GEN_7035 : reservedValidList4_13; // @[decode.scala 431:29 330:31]
  wire  _GEN_8156 = 3'h3 == branchTracker ? _GEN_7036 : reservedValidList4_14; // @[decode.scala 431:29 330:31]
  wire  _GEN_8157 = 3'h3 == branchTracker ? _GEN_7037 : reservedValidList4_15; // @[decode.scala 431:29 330:31]
  wire  _GEN_8158 = 3'h3 == branchTracker ? _GEN_7038 : reservedValidList4_16; // @[decode.scala 431:29 330:31]
  wire  _GEN_8159 = 3'h3 == branchTracker ? _GEN_7039 : reservedValidList4_17; // @[decode.scala 431:29 330:31]
  wire  _GEN_8160 = 3'h3 == branchTracker ? _GEN_7040 : reservedValidList4_18; // @[decode.scala 431:29 330:31]
  wire  _GEN_8161 = 3'h3 == branchTracker ? _GEN_7041 : reservedValidList4_19; // @[decode.scala 431:29 330:31]
  wire  _GEN_8162 = 3'h3 == branchTracker ? _GEN_7042 : reservedValidList4_20; // @[decode.scala 431:29 330:31]
  wire  _GEN_8163 = 3'h3 == branchTracker ? _GEN_7043 : reservedValidList4_21; // @[decode.scala 431:29 330:31]
  wire  _GEN_8164 = 3'h3 == branchTracker ? _GEN_7044 : reservedValidList4_22; // @[decode.scala 431:29 330:31]
  wire  _GEN_8165 = 3'h3 == branchTracker ? _GEN_7045 : reservedValidList4_23; // @[decode.scala 431:29 330:31]
  wire  _GEN_8166 = 3'h3 == branchTracker ? _GEN_7046 : reservedValidList4_24; // @[decode.scala 431:29 330:31]
  wire  _GEN_8167 = 3'h3 == branchTracker ? _GEN_7047 : reservedValidList4_25; // @[decode.scala 431:29 330:31]
  wire  _GEN_8168 = 3'h3 == branchTracker ? _GEN_7048 : reservedValidList4_26; // @[decode.scala 431:29 330:31]
  wire  _GEN_8169 = 3'h3 == branchTracker ? _GEN_7049 : reservedValidList4_27; // @[decode.scala 431:29 330:31]
  wire  _GEN_8170 = 3'h3 == branchTracker ? _GEN_7050 : reservedValidList4_28; // @[decode.scala 431:29 330:31]
  wire  _GEN_8171 = 3'h3 == branchTracker ? _GEN_7051 : reservedValidList4_29; // @[decode.scala 431:29 330:31]
  wire  _GEN_8172 = 3'h3 == branchTracker ? _GEN_7052 : reservedValidList4_30; // @[decode.scala 431:29 330:31]
  wire  _GEN_8173 = 3'h3 == branchTracker ? _GEN_7053 : reservedValidList4_31; // @[decode.scala 431:29 330:31]
  wire  _GEN_8174 = 3'h3 == branchTracker ? _GEN_7054 : reservedValidList4_32; // @[decode.scala 431:29 330:31]
  wire  _GEN_8175 = 3'h3 == branchTracker ? _GEN_7055 : reservedValidList4_33; // @[decode.scala 431:29 330:31]
  wire  _GEN_8176 = 3'h3 == branchTracker ? _GEN_7056 : reservedValidList4_34; // @[decode.scala 431:29 330:31]
  wire  _GEN_8177 = 3'h3 == branchTracker ? _GEN_7057 : reservedValidList4_35; // @[decode.scala 431:29 330:31]
  wire  _GEN_8178 = 3'h3 == branchTracker ? _GEN_7058 : reservedValidList4_36; // @[decode.scala 431:29 330:31]
  wire  _GEN_8179 = 3'h3 == branchTracker ? _GEN_7059 : reservedValidList4_37; // @[decode.scala 431:29 330:31]
  wire  _GEN_8180 = 3'h3 == branchTracker ? _GEN_7060 : reservedValidList4_38; // @[decode.scala 431:29 330:31]
  wire  _GEN_8181 = 3'h3 == branchTracker ? _GEN_7061 : reservedValidList4_39; // @[decode.scala 431:29 330:31]
  wire  _GEN_8182 = 3'h3 == branchTracker ? _GEN_7062 : reservedValidList4_40; // @[decode.scala 431:29 330:31]
  wire  _GEN_8183 = 3'h3 == branchTracker ? _GEN_7063 : reservedValidList4_41; // @[decode.scala 431:29 330:31]
  wire  _GEN_8184 = 3'h3 == branchTracker ? _GEN_7064 : reservedValidList4_42; // @[decode.scala 431:29 330:31]
  wire  _GEN_8185 = 3'h3 == branchTracker ? _GEN_7065 : reservedValidList4_43; // @[decode.scala 431:29 330:31]
  wire  _GEN_8186 = 3'h3 == branchTracker ? _GEN_7066 : reservedValidList4_44; // @[decode.scala 431:29 330:31]
  wire  _GEN_8187 = 3'h3 == branchTracker ? _GEN_7067 : reservedValidList4_45; // @[decode.scala 431:29 330:31]
  wire  _GEN_8188 = 3'h3 == branchTracker ? _GEN_7068 : reservedValidList4_46; // @[decode.scala 431:29 330:31]
  wire  _GEN_8189 = 3'h3 == branchTracker ? _GEN_7069 : reservedValidList4_47; // @[decode.scala 431:29 330:31]
  wire  _GEN_8190 = 3'h3 == branchTracker ? _GEN_7070 : reservedValidList4_48; // @[decode.scala 431:29 330:31]
  wire  _GEN_8191 = 3'h3 == branchTracker ? _GEN_7071 : reservedValidList4_49; // @[decode.scala 431:29 330:31]
  wire  _GEN_8192 = 3'h3 == branchTracker ? _GEN_7072 : reservedValidList4_50; // @[decode.scala 431:29 330:31]
  wire  _GEN_8193 = 3'h3 == branchTracker ? _GEN_7073 : reservedValidList4_51; // @[decode.scala 431:29 330:31]
  wire  _GEN_8194 = 3'h3 == branchTracker ? _GEN_7074 : reservedValidList4_52; // @[decode.scala 431:29 330:31]
  wire  _GEN_8195 = 3'h3 == branchTracker ? _GEN_7075 : reservedValidList4_53; // @[decode.scala 431:29 330:31]
  wire  _GEN_8196 = 3'h3 == branchTracker ? _GEN_7076 : reservedValidList4_54; // @[decode.scala 431:29 330:31]
  wire  _GEN_8197 = 3'h3 == branchTracker ? _GEN_7077 : reservedValidList4_55; // @[decode.scala 431:29 330:31]
  wire  _GEN_8198 = 3'h3 == branchTracker ? _GEN_7078 : reservedValidList4_56; // @[decode.scala 431:29 330:31]
  wire  _GEN_8199 = 3'h3 == branchTracker ? _GEN_7079 : reservedValidList4_57; // @[decode.scala 431:29 330:31]
  wire  _GEN_8200 = 3'h3 == branchTracker ? _GEN_7080 : reservedValidList4_58; // @[decode.scala 431:29 330:31]
  wire  _GEN_8201 = 3'h3 == branchTracker ? _GEN_7081 : reservedValidList4_59; // @[decode.scala 431:29 330:31]
  wire  _GEN_8202 = 3'h3 == branchTracker ? _GEN_7082 : reservedValidList4_60; // @[decode.scala 431:29 330:31]
  wire  _GEN_8203 = 3'h3 == branchTracker ? _GEN_7083 : reservedValidList4_61; // @[decode.scala 431:29 330:31]
  wire  _GEN_8204 = 3'h3 == branchTracker ? _GEN_7084 : reservedValidList4_62; // @[decode.scala 431:29 330:31]
  wire  _GEN_8205 = 3'h3 == branchTracker ? _GEN_7085 : reservedValidList4_63; // @[decode.scala 431:29 330:31]
  wire [5:0] _GEN_8206 = 3'h2 == branchTracker ? _GEN_6926 : _GEN_6341; // @[decode.scala 431:29]
  wire [5:0] _GEN_8207 = 3'h2 == branchTracker ? _GEN_6927 : _GEN_6342; // @[decode.scala 431:29]
  wire [5:0] _GEN_8208 = 3'h2 == branchTracker ? _GEN_6928 : _GEN_6343; // @[decode.scala 431:29]
  wire [5:0] _GEN_8209 = 3'h2 == branchTracker ? _GEN_6929 : _GEN_6344; // @[decode.scala 431:29]
  wire [5:0] _GEN_8210 = 3'h2 == branchTracker ? _GEN_6930 : _GEN_6345; // @[decode.scala 431:29]
  wire [5:0] _GEN_8211 = 3'h2 == branchTracker ? _GEN_6931 : _GEN_6346; // @[decode.scala 431:29]
  wire [5:0] _GEN_8212 = 3'h2 == branchTracker ? _GEN_6932 : _GEN_6347; // @[decode.scala 431:29]
  wire [5:0] _GEN_8213 = 3'h2 == branchTracker ? _GEN_6933 : _GEN_6348; // @[decode.scala 431:29]
  wire [5:0] _GEN_8214 = 3'h2 == branchTracker ? _GEN_6934 : _GEN_6349; // @[decode.scala 431:29]
  wire [5:0] _GEN_8215 = 3'h2 == branchTracker ? _GEN_6935 : _GEN_6350; // @[decode.scala 431:29]
  wire [5:0] _GEN_8216 = 3'h2 == branchTracker ? _GEN_6936 : _GEN_6351; // @[decode.scala 431:29]
  wire [5:0] _GEN_8217 = 3'h2 == branchTracker ? _GEN_6937 : _GEN_6352; // @[decode.scala 431:29]
  wire [5:0] _GEN_8218 = 3'h2 == branchTracker ? _GEN_6938 : _GEN_6353; // @[decode.scala 431:29]
  wire [5:0] _GEN_8219 = 3'h2 == branchTracker ? _GEN_6939 : _GEN_6354; // @[decode.scala 431:29]
  wire [5:0] _GEN_8220 = 3'h2 == branchTracker ? _GEN_6940 : _GEN_6355; // @[decode.scala 431:29]
  wire [5:0] _GEN_8221 = 3'h2 == branchTracker ? _GEN_6941 : _GEN_6356; // @[decode.scala 431:29]
  wire [5:0] _GEN_8222 = 3'h2 == branchTracker ? _GEN_6942 : _GEN_6357; // @[decode.scala 431:29]
  wire [5:0] _GEN_8223 = 3'h2 == branchTracker ? _GEN_6943 : _GEN_6358; // @[decode.scala 431:29]
  wire [5:0] _GEN_8224 = 3'h2 == branchTracker ? _GEN_6944 : _GEN_6359; // @[decode.scala 431:29]
  wire [5:0] _GEN_8225 = 3'h2 == branchTracker ? _GEN_6945 : _GEN_6360; // @[decode.scala 431:29]
  wire [5:0] _GEN_8226 = 3'h2 == branchTracker ? _GEN_6946 : _GEN_6361; // @[decode.scala 431:29]
  wire [5:0] _GEN_8227 = 3'h2 == branchTracker ? _GEN_6947 : _GEN_6362; // @[decode.scala 431:29]
  wire [5:0] _GEN_8228 = 3'h2 == branchTracker ? _GEN_6948 : _GEN_6363; // @[decode.scala 431:29]
  wire [5:0] _GEN_8229 = 3'h2 == branchTracker ? _GEN_6949 : _GEN_6364; // @[decode.scala 431:29]
  wire [5:0] _GEN_8230 = 3'h2 == branchTracker ? _GEN_6950 : _GEN_6365; // @[decode.scala 431:29]
  wire [5:0] _GEN_8231 = 3'h2 == branchTracker ? _GEN_6951 : _GEN_6366; // @[decode.scala 431:29]
  wire [5:0] _GEN_8232 = 3'h2 == branchTracker ? _GEN_6952 : _GEN_6367; // @[decode.scala 431:29]
  wire [5:0] _GEN_8233 = 3'h2 == branchTracker ? _GEN_6953 : _GEN_6368; // @[decode.scala 431:29]
  wire [5:0] _GEN_8234 = 3'h2 == branchTracker ? _GEN_6954 : _GEN_6369; // @[decode.scala 431:29]
  wire [5:0] _GEN_8235 = 3'h2 == branchTracker ? _GEN_6955 : _GEN_6370; // @[decode.scala 431:29]
  wire [5:0] _GEN_8236 = 3'h2 == branchTracker ? _GEN_6956 : _GEN_6371; // @[decode.scala 431:29]
  wire [5:0] _GEN_8237 = 3'h2 == branchTracker ? _GEN_6957 : _GEN_6372; // @[decode.scala 431:29]
  wire  _GEN_8238 = 3'h2 == branchTracker ? _GEN_6958 : _GEN_6501; // @[decode.scala 431:29]
  wire  _GEN_8239 = 3'h2 == branchTracker ? _GEN_6959 : _GEN_6502; // @[decode.scala 431:29]
  wire  _GEN_8240 = 3'h2 == branchTracker ? _GEN_6960 : _GEN_6503; // @[decode.scala 431:29]
  wire  _GEN_8241 = 3'h2 == branchTracker ? _GEN_6961 : _GEN_6504; // @[decode.scala 431:29]
  wire  _GEN_8242 = 3'h2 == branchTracker ? _GEN_6962 : _GEN_6505; // @[decode.scala 431:29]
  wire  _GEN_8243 = 3'h2 == branchTracker ? _GEN_6963 : _GEN_6506; // @[decode.scala 431:29]
  wire  _GEN_8244 = 3'h2 == branchTracker ? _GEN_6964 : _GEN_6507; // @[decode.scala 431:29]
  wire  _GEN_8245 = 3'h2 == branchTracker ? _GEN_6965 : _GEN_6508; // @[decode.scala 431:29]
  wire  _GEN_8246 = 3'h2 == branchTracker ? _GEN_6966 : _GEN_6509; // @[decode.scala 431:29]
  wire  _GEN_8247 = 3'h2 == branchTracker ? _GEN_6967 : _GEN_6510; // @[decode.scala 431:29]
  wire  _GEN_8248 = 3'h2 == branchTracker ? _GEN_6968 : _GEN_6511; // @[decode.scala 431:29]
  wire  _GEN_8249 = 3'h2 == branchTracker ? _GEN_6969 : _GEN_6512; // @[decode.scala 431:29]
  wire  _GEN_8250 = 3'h2 == branchTracker ? _GEN_6970 : _GEN_6513; // @[decode.scala 431:29]
  wire  _GEN_8251 = 3'h2 == branchTracker ? _GEN_6971 : _GEN_6514; // @[decode.scala 431:29]
  wire  _GEN_8252 = 3'h2 == branchTracker ? _GEN_6972 : _GEN_6515; // @[decode.scala 431:29]
  wire  _GEN_8253 = 3'h2 == branchTracker ? _GEN_6973 : _GEN_6516; // @[decode.scala 431:29]
  wire  _GEN_8254 = 3'h2 == branchTracker ? _GEN_6974 : _GEN_6517; // @[decode.scala 431:29]
  wire  _GEN_8255 = 3'h2 == branchTracker ? _GEN_6975 : _GEN_6518; // @[decode.scala 431:29]
  wire  _GEN_8256 = 3'h2 == branchTracker ? _GEN_6976 : _GEN_6519; // @[decode.scala 431:29]
  wire  _GEN_8257 = 3'h2 == branchTracker ? _GEN_6977 : _GEN_6520; // @[decode.scala 431:29]
  wire  _GEN_8258 = 3'h2 == branchTracker ? _GEN_6978 : _GEN_6521; // @[decode.scala 431:29]
  wire  _GEN_8259 = 3'h2 == branchTracker ? _GEN_6979 : _GEN_6522; // @[decode.scala 431:29]
  wire  _GEN_8260 = 3'h2 == branchTracker ? _GEN_6980 : _GEN_6523; // @[decode.scala 431:29]
  wire  _GEN_8261 = 3'h2 == branchTracker ? _GEN_6981 : _GEN_6524; // @[decode.scala 431:29]
  wire  _GEN_8262 = 3'h2 == branchTracker ? _GEN_6982 : _GEN_6525; // @[decode.scala 431:29]
  wire  _GEN_8263 = 3'h2 == branchTracker ? _GEN_6983 : _GEN_6526; // @[decode.scala 431:29]
  wire  _GEN_8264 = 3'h2 == branchTracker ? _GEN_6984 : _GEN_6527; // @[decode.scala 431:29]
  wire  _GEN_8265 = 3'h2 == branchTracker ? _GEN_6985 : _GEN_6528; // @[decode.scala 431:29]
  wire  _GEN_8266 = 3'h2 == branchTracker ? _GEN_6986 : _GEN_6529; // @[decode.scala 431:29]
  wire  _GEN_8267 = 3'h2 == branchTracker ? _GEN_6987 : _GEN_6530; // @[decode.scala 431:29]
  wire  _GEN_8268 = 3'h2 == branchTracker ? _GEN_6988 : _GEN_6531; // @[decode.scala 431:29]
  wire  _GEN_8269 = 3'h2 == branchTracker ? _GEN_6989 : _GEN_6532; // @[decode.scala 431:29]
  wire  _GEN_8270 = 3'h2 == branchTracker ? _GEN_6990 : _GEN_6533; // @[decode.scala 431:29]
  wire  _GEN_8271 = 3'h2 == branchTracker ? _GEN_6991 : _GEN_6534; // @[decode.scala 431:29]
  wire  _GEN_8272 = 3'h2 == branchTracker ? _GEN_6992 : _GEN_6535; // @[decode.scala 431:29]
  wire  _GEN_8273 = 3'h2 == branchTracker ? _GEN_6993 : _GEN_6536; // @[decode.scala 431:29]
  wire  _GEN_8274 = 3'h2 == branchTracker ? _GEN_6994 : _GEN_6537; // @[decode.scala 431:29]
  wire  _GEN_8275 = 3'h2 == branchTracker ? _GEN_6995 : _GEN_6538; // @[decode.scala 431:29]
  wire  _GEN_8276 = 3'h2 == branchTracker ? _GEN_6996 : _GEN_6539; // @[decode.scala 431:29]
  wire  _GEN_8277 = 3'h2 == branchTracker ? _GEN_6997 : _GEN_6540; // @[decode.scala 431:29]
  wire  _GEN_8278 = 3'h2 == branchTracker ? _GEN_6998 : _GEN_6541; // @[decode.scala 431:29]
  wire  _GEN_8279 = 3'h2 == branchTracker ? _GEN_6999 : _GEN_6542; // @[decode.scala 431:29]
  wire  _GEN_8280 = 3'h2 == branchTracker ? _GEN_7000 : _GEN_6543; // @[decode.scala 431:29]
  wire  _GEN_8281 = 3'h2 == branchTracker ? _GEN_7001 : _GEN_6544; // @[decode.scala 431:29]
  wire  _GEN_8282 = 3'h2 == branchTracker ? _GEN_7002 : _GEN_6545; // @[decode.scala 431:29]
  wire  _GEN_8283 = 3'h2 == branchTracker ? _GEN_7003 : _GEN_6546; // @[decode.scala 431:29]
  wire  _GEN_8284 = 3'h2 == branchTracker ? _GEN_7004 : _GEN_6547; // @[decode.scala 431:29]
  wire  _GEN_8285 = 3'h2 == branchTracker ? _GEN_7005 : _GEN_6548; // @[decode.scala 431:29]
  wire  _GEN_8286 = 3'h2 == branchTracker ? _GEN_7006 : _GEN_6549; // @[decode.scala 431:29]
  wire  _GEN_8287 = 3'h2 == branchTracker ? _GEN_7007 : _GEN_6550; // @[decode.scala 431:29]
  wire  _GEN_8288 = 3'h2 == branchTracker ? _GEN_7008 : _GEN_6551; // @[decode.scala 431:29]
  wire  _GEN_8289 = 3'h2 == branchTracker ? _GEN_7009 : _GEN_6552; // @[decode.scala 431:29]
  wire  _GEN_8290 = 3'h2 == branchTracker ? _GEN_7010 : _GEN_6553; // @[decode.scala 431:29]
  wire  _GEN_8291 = 3'h2 == branchTracker ? _GEN_7011 : _GEN_6554; // @[decode.scala 431:29]
  wire  _GEN_8292 = 3'h2 == branchTracker ? _GEN_7012 : _GEN_6555; // @[decode.scala 431:29]
  wire  _GEN_8293 = 3'h2 == branchTracker ? _GEN_7013 : _GEN_6556; // @[decode.scala 431:29]
  wire  _GEN_8294 = 3'h2 == branchTracker ? _GEN_7014 : _GEN_6557; // @[decode.scala 431:29]
  wire  _GEN_8295 = 3'h2 == branchTracker ? _GEN_7015 : _GEN_6558; // @[decode.scala 431:29]
  wire  _GEN_8296 = 3'h2 == branchTracker ? _GEN_7016 : _GEN_6559; // @[decode.scala 431:29]
  wire  _GEN_8297 = 3'h2 == branchTracker ? _GEN_7017 : _GEN_6560; // @[decode.scala 431:29]
  wire  _GEN_8298 = 3'h2 == branchTracker ? _GEN_7018 : _GEN_6561; // @[decode.scala 431:29]
  wire  _GEN_8299 = 3'h2 == branchTracker ? _GEN_7019 : _GEN_6562; // @[decode.scala 431:29]
  wire  _GEN_8300 = 3'h2 == branchTracker ? _GEN_7020 : _GEN_6563; // @[decode.scala 431:29]
  wire  _GEN_8302 = 3'h2 == branchTracker ? _GEN_7022 : _GEN_6693; // @[decode.scala 431:29]
  wire  _GEN_8303 = 3'h2 == branchTracker ? _GEN_7023 : _GEN_6694; // @[decode.scala 431:29]
  wire  _GEN_8304 = 3'h2 == branchTracker ? _GEN_7024 : _GEN_6695; // @[decode.scala 431:29]
  wire  _GEN_8305 = 3'h2 == branchTracker ? _GEN_7025 : _GEN_6696; // @[decode.scala 431:29]
  wire  _GEN_8306 = 3'h2 == branchTracker ? _GEN_7026 : _GEN_6697; // @[decode.scala 431:29]
  wire  _GEN_8307 = 3'h2 == branchTracker ? _GEN_7027 : _GEN_6698; // @[decode.scala 431:29]
  wire  _GEN_8308 = 3'h2 == branchTracker ? _GEN_7028 : _GEN_6699; // @[decode.scala 431:29]
  wire  _GEN_8309 = 3'h2 == branchTracker ? _GEN_7029 : _GEN_6700; // @[decode.scala 431:29]
  wire  _GEN_8310 = 3'h2 == branchTracker ? _GEN_7030 : _GEN_6701; // @[decode.scala 431:29]
  wire  _GEN_8311 = 3'h2 == branchTracker ? _GEN_7031 : _GEN_6702; // @[decode.scala 431:29]
  wire  _GEN_8312 = 3'h2 == branchTracker ? _GEN_7032 : _GEN_6703; // @[decode.scala 431:29]
  wire  _GEN_8313 = 3'h2 == branchTracker ? _GEN_7033 : _GEN_6704; // @[decode.scala 431:29]
  wire  _GEN_8314 = 3'h2 == branchTracker ? _GEN_7034 : _GEN_6705; // @[decode.scala 431:29]
  wire  _GEN_8315 = 3'h2 == branchTracker ? _GEN_7035 : _GEN_6706; // @[decode.scala 431:29]
  wire  _GEN_8316 = 3'h2 == branchTracker ? _GEN_7036 : _GEN_6707; // @[decode.scala 431:29]
  wire  _GEN_8317 = 3'h2 == branchTracker ? _GEN_7037 : _GEN_6708; // @[decode.scala 431:29]
  wire  _GEN_8318 = 3'h2 == branchTracker ? _GEN_7038 : _GEN_6709; // @[decode.scala 431:29]
  wire  _GEN_8319 = 3'h2 == branchTracker ? _GEN_7039 : _GEN_6710; // @[decode.scala 431:29]
  wire  _GEN_8320 = 3'h2 == branchTracker ? _GEN_7040 : _GEN_6711; // @[decode.scala 431:29]
  wire  _GEN_8321 = 3'h2 == branchTracker ? _GEN_7041 : _GEN_6712; // @[decode.scala 431:29]
  wire  _GEN_8322 = 3'h2 == branchTracker ? _GEN_7042 : _GEN_6713; // @[decode.scala 431:29]
  wire  _GEN_8323 = 3'h2 == branchTracker ? _GEN_7043 : _GEN_6714; // @[decode.scala 431:29]
  wire  _GEN_8324 = 3'h2 == branchTracker ? _GEN_7044 : _GEN_6715; // @[decode.scala 431:29]
  wire  _GEN_8325 = 3'h2 == branchTracker ? _GEN_7045 : _GEN_6716; // @[decode.scala 431:29]
  wire  _GEN_8326 = 3'h2 == branchTracker ? _GEN_7046 : _GEN_6717; // @[decode.scala 431:29]
  wire  _GEN_8327 = 3'h2 == branchTracker ? _GEN_7047 : _GEN_6718; // @[decode.scala 431:29]
  wire  _GEN_8328 = 3'h2 == branchTracker ? _GEN_7048 : _GEN_6719; // @[decode.scala 431:29]
  wire  _GEN_8329 = 3'h2 == branchTracker ? _GEN_7049 : _GEN_6720; // @[decode.scala 431:29]
  wire  _GEN_8330 = 3'h2 == branchTracker ? _GEN_7050 : _GEN_6721; // @[decode.scala 431:29]
  wire  _GEN_8331 = 3'h2 == branchTracker ? _GEN_7051 : _GEN_6722; // @[decode.scala 431:29]
  wire  _GEN_8332 = 3'h2 == branchTracker ? _GEN_7052 : _GEN_6723; // @[decode.scala 431:29]
  wire  _GEN_8333 = 3'h2 == branchTracker ? _GEN_7053 : _GEN_6724; // @[decode.scala 431:29]
  wire  _GEN_8334 = 3'h2 == branchTracker ? _GEN_7054 : _GEN_6725; // @[decode.scala 431:29]
  wire  _GEN_8335 = 3'h2 == branchTracker ? _GEN_7055 : _GEN_6726; // @[decode.scala 431:29]
  wire  _GEN_8336 = 3'h2 == branchTracker ? _GEN_7056 : _GEN_6727; // @[decode.scala 431:29]
  wire  _GEN_8337 = 3'h2 == branchTracker ? _GEN_7057 : _GEN_6728; // @[decode.scala 431:29]
  wire  _GEN_8338 = 3'h2 == branchTracker ? _GEN_7058 : _GEN_6729; // @[decode.scala 431:29]
  wire  _GEN_8339 = 3'h2 == branchTracker ? _GEN_7059 : _GEN_6730; // @[decode.scala 431:29]
  wire  _GEN_8340 = 3'h2 == branchTracker ? _GEN_7060 : _GEN_6731; // @[decode.scala 431:29]
  wire  _GEN_8341 = 3'h2 == branchTracker ? _GEN_7061 : _GEN_6732; // @[decode.scala 431:29]
  wire  _GEN_8342 = 3'h2 == branchTracker ? _GEN_7062 : _GEN_6733; // @[decode.scala 431:29]
  wire  _GEN_8343 = 3'h2 == branchTracker ? _GEN_7063 : _GEN_6734; // @[decode.scala 431:29]
  wire  _GEN_8344 = 3'h2 == branchTracker ? _GEN_7064 : _GEN_6735; // @[decode.scala 431:29]
  wire  _GEN_8345 = 3'h2 == branchTracker ? _GEN_7065 : _GEN_6736; // @[decode.scala 431:29]
  wire  _GEN_8346 = 3'h2 == branchTracker ? _GEN_7066 : _GEN_6737; // @[decode.scala 431:29]
  wire  _GEN_8347 = 3'h2 == branchTracker ? _GEN_7067 : _GEN_6738; // @[decode.scala 431:29]
  wire  _GEN_8348 = 3'h2 == branchTracker ? _GEN_7068 : _GEN_6739; // @[decode.scala 431:29]
  wire  _GEN_8349 = 3'h2 == branchTracker ? _GEN_7069 : _GEN_6740; // @[decode.scala 431:29]
  wire  _GEN_8350 = 3'h2 == branchTracker ? _GEN_7070 : _GEN_6741; // @[decode.scala 431:29]
  wire  _GEN_8351 = 3'h2 == branchTracker ? _GEN_7071 : _GEN_6742; // @[decode.scala 431:29]
  wire  _GEN_8352 = 3'h2 == branchTracker ? _GEN_7072 : _GEN_6743; // @[decode.scala 431:29]
  wire  _GEN_8353 = 3'h2 == branchTracker ? _GEN_7073 : _GEN_6744; // @[decode.scala 431:29]
  wire  _GEN_8354 = 3'h2 == branchTracker ? _GEN_7074 : _GEN_6745; // @[decode.scala 431:29]
  wire  _GEN_8355 = 3'h2 == branchTracker ? _GEN_7075 : _GEN_6746; // @[decode.scala 431:29]
  wire  _GEN_8356 = 3'h2 == branchTracker ? _GEN_7076 : _GEN_6747; // @[decode.scala 431:29]
  wire  _GEN_8357 = 3'h2 == branchTracker ? _GEN_7077 : _GEN_6748; // @[decode.scala 431:29]
  wire  _GEN_8358 = 3'h2 == branchTracker ? _GEN_7078 : _GEN_6749; // @[decode.scala 431:29]
  wire  _GEN_8359 = 3'h2 == branchTracker ? _GEN_7079 : _GEN_6750; // @[decode.scala 431:29]
  wire  _GEN_8360 = 3'h2 == branchTracker ? _GEN_7080 : _GEN_6751; // @[decode.scala 431:29]
  wire  _GEN_8361 = 3'h2 == branchTracker ? _GEN_7081 : _GEN_6752; // @[decode.scala 431:29]
  wire  _GEN_8362 = 3'h2 == branchTracker ? _GEN_7082 : _GEN_6753; // @[decode.scala 431:29]
  wire  _GEN_8363 = 3'h2 == branchTracker ? _GEN_7083 : _GEN_6754; // @[decode.scala 431:29]
  wire  _GEN_8364 = 3'h2 == branchTracker ? _GEN_7084 : _GEN_6755; // @[decode.scala 431:29]
  wire  _GEN_8365 = 3'h2 == branchTracker ? _GEN_7085 : _GEN_6756; // @[decode.scala 431:29]
  wire [5:0] _GEN_8366 = 3'h2 == branchTracker ? reservedRegMap4_0 : _GEN_8046; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8367 = 3'h2 == branchTracker ? reservedRegMap4_1 : _GEN_8047; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8368 = 3'h2 == branchTracker ? reservedRegMap4_2 : _GEN_8048; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8369 = 3'h2 == branchTracker ? reservedRegMap4_3 : _GEN_8049; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8370 = 3'h2 == branchTracker ? reservedRegMap4_4 : _GEN_8050; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8371 = 3'h2 == branchTracker ? reservedRegMap4_5 : _GEN_8051; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8372 = 3'h2 == branchTracker ? reservedRegMap4_6 : _GEN_8052; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8373 = 3'h2 == branchTracker ? reservedRegMap4_7 : _GEN_8053; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8374 = 3'h2 == branchTracker ? reservedRegMap4_8 : _GEN_8054; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8375 = 3'h2 == branchTracker ? reservedRegMap4_9 : _GEN_8055; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8376 = 3'h2 == branchTracker ? reservedRegMap4_10 : _GEN_8056; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8377 = 3'h2 == branchTracker ? reservedRegMap4_11 : _GEN_8057; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8378 = 3'h2 == branchTracker ? reservedRegMap4_12 : _GEN_8058; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8379 = 3'h2 == branchTracker ? reservedRegMap4_13 : _GEN_8059; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8380 = 3'h2 == branchTracker ? reservedRegMap4_14 : _GEN_8060; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8381 = 3'h2 == branchTracker ? reservedRegMap4_15 : _GEN_8061; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8382 = 3'h2 == branchTracker ? reservedRegMap4_16 : _GEN_8062; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8383 = 3'h2 == branchTracker ? reservedRegMap4_17 : _GEN_8063; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8384 = 3'h2 == branchTracker ? reservedRegMap4_18 : _GEN_8064; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8385 = 3'h2 == branchTracker ? reservedRegMap4_19 : _GEN_8065; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8386 = 3'h2 == branchTracker ? reservedRegMap4_20 : _GEN_8066; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8387 = 3'h2 == branchTracker ? reservedRegMap4_21 : _GEN_8067; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8388 = 3'h2 == branchTracker ? reservedRegMap4_22 : _GEN_8068; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8389 = 3'h2 == branchTracker ? reservedRegMap4_23 : _GEN_8069; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8390 = 3'h2 == branchTracker ? reservedRegMap4_24 : _GEN_8070; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8391 = 3'h2 == branchTracker ? reservedRegMap4_25 : _GEN_8071; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8392 = 3'h2 == branchTracker ? reservedRegMap4_26 : _GEN_8072; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8393 = 3'h2 == branchTracker ? reservedRegMap4_27 : _GEN_8073; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8394 = 3'h2 == branchTracker ? reservedRegMap4_28 : _GEN_8074; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8395 = 3'h2 == branchTracker ? reservedRegMap4_29 : _GEN_8075; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8396 = 3'h2 == branchTracker ? reservedRegMap4_30 : _GEN_8076; // @[decode.scala 320:28 431:29]
  wire [5:0] _GEN_8397 = 3'h2 == branchTracker ? reservedRegMap4_31 : _GEN_8077; // @[decode.scala 320:28 431:29]
  wire  _GEN_8398 = 3'h2 == branchTracker ? reservedFreeList4_0 : _GEN_8078; // @[decode.scala 431:29 325:30]
  wire  _GEN_8399 = 3'h2 == branchTracker ? reservedFreeList4_1 : _GEN_8079; // @[decode.scala 431:29 325:30]
  wire  _GEN_8400 = 3'h2 == branchTracker ? reservedFreeList4_2 : _GEN_8080; // @[decode.scala 431:29 325:30]
  wire  _GEN_8401 = 3'h2 == branchTracker ? reservedFreeList4_3 : _GEN_8081; // @[decode.scala 431:29 325:30]
  wire  _GEN_8402 = 3'h2 == branchTracker ? reservedFreeList4_4 : _GEN_8082; // @[decode.scala 431:29 325:30]
  wire  _GEN_8403 = 3'h2 == branchTracker ? reservedFreeList4_5 : _GEN_8083; // @[decode.scala 431:29 325:30]
  wire  _GEN_8404 = 3'h2 == branchTracker ? reservedFreeList4_6 : _GEN_8084; // @[decode.scala 431:29 325:30]
  wire  _GEN_8405 = 3'h2 == branchTracker ? reservedFreeList4_7 : _GEN_8085; // @[decode.scala 431:29 325:30]
  wire  _GEN_8406 = 3'h2 == branchTracker ? reservedFreeList4_8 : _GEN_8086; // @[decode.scala 431:29 325:30]
  wire  _GEN_8407 = 3'h2 == branchTracker ? reservedFreeList4_9 : _GEN_8087; // @[decode.scala 431:29 325:30]
  wire  _GEN_8408 = 3'h2 == branchTracker ? reservedFreeList4_10 : _GEN_8088; // @[decode.scala 431:29 325:30]
  wire  _GEN_8409 = 3'h2 == branchTracker ? reservedFreeList4_11 : _GEN_8089; // @[decode.scala 431:29 325:30]
  wire  _GEN_8410 = 3'h2 == branchTracker ? reservedFreeList4_12 : _GEN_8090; // @[decode.scala 431:29 325:30]
  wire  _GEN_8411 = 3'h2 == branchTracker ? reservedFreeList4_13 : _GEN_8091; // @[decode.scala 431:29 325:30]
  wire  _GEN_8412 = 3'h2 == branchTracker ? reservedFreeList4_14 : _GEN_8092; // @[decode.scala 431:29 325:30]
  wire  _GEN_8413 = 3'h2 == branchTracker ? reservedFreeList4_15 : _GEN_8093; // @[decode.scala 431:29 325:30]
  wire  _GEN_8414 = 3'h2 == branchTracker ? reservedFreeList4_16 : _GEN_8094; // @[decode.scala 431:29 325:30]
  wire  _GEN_8415 = 3'h2 == branchTracker ? reservedFreeList4_17 : _GEN_8095; // @[decode.scala 431:29 325:30]
  wire  _GEN_8416 = 3'h2 == branchTracker ? reservedFreeList4_18 : _GEN_8096; // @[decode.scala 431:29 325:30]
  wire  _GEN_8417 = 3'h2 == branchTracker ? reservedFreeList4_19 : _GEN_8097; // @[decode.scala 431:29 325:30]
  wire  _GEN_8418 = 3'h2 == branchTracker ? reservedFreeList4_20 : _GEN_8098; // @[decode.scala 431:29 325:30]
  wire  _GEN_8419 = 3'h2 == branchTracker ? reservedFreeList4_21 : _GEN_8099; // @[decode.scala 431:29 325:30]
  wire  _GEN_8420 = 3'h2 == branchTracker ? reservedFreeList4_22 : _GEN_8100; // @[decode.scala 431:29 325:30]
  wire  _GEN_8421 = 3'h2 == branchTracker ? reservedFreeList4_23 : _GEN_8101; // @[decode.scala 431:29 325:30]
  wire  _GEN_8422 = 3'h2 == branchTracker ? reservedFreeList4_24 : _GEN_8102; // @[decode.scala 431:29 325:30]
  wire  _GEN_8423 = 3'h2 == branchTracker ? reservedFreeList4_25 : _GEN_8103; // @[decode.scala 431:29 325:30]
  wire  _GEN_8424 = 3'h2 == branchTracker ? reservedFreeList4_26 : _GEN_8104; // @[decode.scala 431:29 325:30]
  wire  _GEN_8425 = 3'h2 == branchTracker ? reservedFreeList4_27 : _GEN_8105; // @[decode.scala 431:29 325:30]
  wire  _GEN_8426 = 3'h2 == branchTracker ? reservedFreeList4_28 : _GEN_8106; // @[decode.scala 431:29 325:30]
  wire  _GEN_8427 = 3'h2 == branchTracker ? reservedFreeList4_29 : _GEN_8107; // @[decode.scala 431:29 325:30]
  wire  _GEN_8428 = 3'h2 == branchTracker ? reservedFreeList4_30 : _GEN_8108; // @[decode.scala 431:29 325:30]
  wire  _GEN_8429 = 3'h2 == branchTracker ? reservedFreeList4_31 : _GEN_8109; // @[decode.scala 431:29 325:30]
  wire  _GEN_8430 = 3'h2 == branchTracker ? reservedFreeList4_32 : _GEN_8110; // @[decode.scala 431:29 325:30]
  wire  _GEN_8431 = 3'h2 == branchTracker ? reservedFreeList4_33 : _GEN_8111; // @[decode.scala 431:29 325:30]
  wire  _GEN_8432 = 3'h2 == branchTracker ? reservedFreeList4_34 : _GEN_8112; // @[decode.scala 431:29 325:30]
  wire  _GEN_8433 = 3'h2 == branchTracker ? reservedFreeList4_35 : _GEN_8113; // @[decode.scala 431:29 325:30]
  wire  _GEN_8434 = 3'h2 == branchTracker ? reservedFreeList4_36 : _GEN_8114; // @[decode.scala 431:29 325:30]
  wire  _GEN_8435 = 3'h2 == branchTracker ? reservedFreeList4_37 : _GEN_8115; // @[decode.scala 431:29 325:30]
  wire  _GEN_8436 = 3'h2 == branchTracker ? reservedFreeList4_38 : _GEN_8116; // @[decode.scala 431:29 325:30]
  wire  _GEN_8437 = 3'h2 == branchTracker ? reservedFreeList4_39 : _GEN_8117; // @[decode.scala 431:29 325:30]
  wire  _GEN_8438 = 3'h2 == branchTracker ? reservedFreeList4_40 : _GEN_8118; // @[decode.scala 431:29 325:30]
  wire  _GEN_8439 = 3'h2 == branchTracker ? reservedFreeList4_41 : _GEN_8119; // @[decode.scala 431:29 325:30]
  wire  _GEN_8440 = 3'h2 == branchTracker ? reservedFreeList4_42 : _GEN_8120; // @[decode.scala 431:29 325:30]
  wire  _GEN_8441 = 3'h2 == branchTracker ? reservedFreeList4_43 : _GEN_8121; // @[decode.scala 431:29 325:30]
  wire  _GEN_8442 = 3'h2 == branchTracker ? reservedFreeList4_44 : _GEN_8122; // @[decode.scala 431:29 325:30]
  wire  _GEN_8443 = 3'h2 == branchTracker ? reservedFreeList4_45 : _GEN_8123; // @[decode.scala 431:29 325:30]
  wire  _GEN_8444 = 3'h2 == branchTracker ? reservedFreeList4_46 : _GEN_8124; // @[decode.scala 431:29 325:30]
  wire  _GEN_8445 = 3'h2 == branchTracker ? reservedFreeList4_47 : _GEN_8125; // @[decode.scala 431:29 325:30]
  wire  _GEN_8446 = 3'h2 == branchTracker ? reservedFreeList4_48 : _GEN_8126; // @[decode.scala 431:29 325:30]
  wire  _GEN_8447 = 3'h2 == branchTracker ? reservedFreeList4_49 : _GEN_8127; // @[decode.scala 431:29 325:30]
  wire  _GEN_8448 = 3'h2 == branchTracker ? reservedFreeList4_50 : _GEN_8128; // @[decode.scala 431:29 325:30]
  wire  _GEN_8449 = 3'h2 == branchTracker ? reservedFreeList4_51 : _GEN_8129; // @[decode.scala 431:29 325:30]
  wire  _GEN_8450 = 3'h2 == branchTracker ? reservedFreeList4_52 : _GEN_8130; // @[decode.scala 431:29 325:30]
  wire  _GEN_8451 = 3'h2 == branchTracker ? reservedFreeList4_53 : _GEN_8131; // @[decode.scala 431:29 325:30]
  wire  _GEN_8452 = 3'h2 == branchTracker ? reservedFreeList4_54 : _GEN_8132; // @[decode.scala 431:29 325:30]
  wire  _GEN_8453 = 3'h2 == branchTracker ? reservedFreeList4_55 : _GEN_8133; // @[decode.scala 431:29 325:30]
  wire  _GEN_8454 = 3'h2 == branchTracker ? reservedFreeList4_56 : _GEN_8134; // @[decode.scala 431:29 325:30]
  wire  _GEN_8455 = 3'h2 == branchTracker ? reservedFreeList4_57 : _GEN_8135; // @[decode.scala 431:29 325:30]
  wire  _GEN_8456 = 3'h2 == branchTracker ? reservedFreeList4_58 : _GEN_8136; // @[decode.scala 431:29 325:30]
  wire  _GEN_8457 = 3'h2 == branchTracker ? reservedFreeList4_59 : _GEN_8137; // @[decode.scala 431:29 325:30]
  wire  _GEN_8458 = 3'h2 == branchTracker ? reservedFreeList4_60 : _GEN_8138; // @[decode.scala 431:29 325:30]
  wire  _GEN_8459 = 3'h2 == branchTracker ? reservedFreeList4_61 : _GEN_8139; // @[decode.scala 431:29 325:30]
  wire  _GEN_8460 = 3'h2 == branchTracker ? reservedFreeList4_62 : _GEN_8140; // @[decode.scala 431:29 325:30]
  wire  _GEN_8462 = 3'h2 == branchTracker ? reservedValidList4_0 : _GEN_8142; // @[decode.scala 431:29 330:31]
  wire  _GEN_8463 = 3'h2 == branchTracker ? reservedValidList4_1 : _GEN_8143; // @[decode.scala 431:29 330:31]
  wire  _GEN_8464 = 3'h2 == branchTracker ? reservedValidList4_2 : _GEN_8144; // @[decode.scala 431:29 330:31]
  wire  _GEN_8465 = 3'h2 == branchTracker ? reservedValidList4_3 : _GEN_8145; // @[decode.scala 431:29 330:31]
  wire  _GEN_8466 = 3'h2 == branchTracker ? reservedValidList4_4 : _GEN_8146; // @[decode.scala 431:29 330:31]
  wire  _GEN_8467 = 3'h2 == branchTracker ? reservedValidList4_5 : _GEN_8147; // @[decode.scala 431:29 330:31]
  wire  _GEN_8468 = 3'h2 == branchTracker ? reservedValidList4_6 : _GEN_8148; // @[decode.scala 431:29 330:31]
  wire  _GEN_8469 = 3'h2 == branchTracker ? reservedValidList4_7 : _GEN_8149; // @[decode.scala 431:29 330:31]
  wire  _GEN_8470 = 3'h2 == branchTracker ? reservedValidList4_8 : _GEN_8150; // @[decode.scala 431:29 330:31]
  wire  _GEN_8471 = 3'h2 == branchTracker ? reservedValidList4_9 : _GEN_8151; // @[decode.scala 431:29 330:31]
  wire  _GEN_8472 = 3'h2 == branchTracker ? reservedValidList4_10 : _GEN_8152; // @[decode.scala 431:29 330:31]
  wire  _GEN_8473 = 3'h2 == branchTracker ? reservedValidList4_11 : _GEN_8153; // @[decode.scala 431:29 330:31]
  wire  _GEN_8474 = 3'h2 == branchTracker ? reservedValidList4_12 : _GEN_8154; // @[decode.scala 431:29 330:31]
  wire  _GEN_8475 = 3'h2 == branchTracker ? reservedValidList4_13 : _GEN_8155; // @[decode.scala 431:29 330:31]
  wire  _GEN_8476 = 3'h2 == branchTracker ? reservedValidList4_14 : _GEN_8156; // @[decode.scala 431:29 330:31]
  wire  _GEN_8477 = 3'h2 == branchTracker ? reservedValidList4_15 : _GEN_8157; // @[decode.scala 431:29 330:31]
  wire  _GEN_8478 = 3'h2 == branchTracker ? reservedValidList4_16 : _GEN_8158; // @[decode.scala 431:29 330:31]
  wire  _GEN_8479 = 3'h2 == branchTracker ? reservedValidList4_17 : _GEN_8159; // @[decode.scala 431:29 330:31]
  wire  _GEN_8480 = 3'h2 == branchTracker ? reservedValidList4_18 : _GEN_8160; // @[decode.scala 431:29 330:31]
  wire  _GEN_8481 = 3'h2 == branchTracker ? reservedValidList4_19 : _GEN_8161; // @[decode.scala 431:29 330:31]
  wire  _GEN_8482 = 3'h2 == branchTracker ? reservedValidList4_20 : _GEN_8162; // @[decode.scala 431:29 330:31]
  wire  _GEN_8483 = 3'h2 == branchTracker ? reservedValidList4_21 : _GEN_8163; // @[decode.scala 431:29 330:31]
  wire  _GEN_8484 = 3'h2 == branchTracker ? reservedValidList4_22 : _GEN_8164; // @[decode.scala 431:29 330:31]
  wire  _GEN_8485 = 3'h2 == branchTracker ? reservedValidList4_23 : _GEN_8165; // @[decode.scala 431:29 330:31]
  wire  _GEN_8486 = 3'h2 == branchTracker ? reservedValidList4_24 : _GEN_8166; // @[decode.scala 431:29 330:31]
  wire  _GEN_8487 = 3'h2 == branchTracker ? reservedValidList4_25 : _GEN_8167; // @[decode.scala 431:29 330:31]
  wire  _GEN_8488 = 3'h2 == branchTracker ? reservedValidList4_26 : _GEN_8168; // @[decode.scala 431:29 330:31]
  wire  _GEN_8489 = 3'h2 == branchTracker ? reservedValidList4_27 : _GEN_8169; // @[decode.scala 431:29 330:31]
  wire  _GEN_8490 = 3'h2 == branchTracker ? reservedValidList4_28 : _GEN_8170; // @[decode.scala 431:29 330:31]
  wire  _GEN_8491 = 3'h2 == branchTracker ? reservedValidList4_29 : _GEN_8171; // @[decode.scala 431:29 330:31]
  wire  _GEN_8492 = 3'h2 == branchTracker ? reservedValidList4_30 : _GEN_8172; // @[decode.scala 431:29 330:31]
  wire  _GEN_8493 = 3'h2 == branchTracker ? reservedValidList4_31 : _GEN_8173; // @[decode.scala 431:29 330:31]
  wire  _GEN_8494 = 3'h2 == branchTracker ? reservedValidList4_32 : _GEN_8174; // @[decode.scala 431:29 330:31]
  wire  _GEN_8495 = 3'h2 == branchTracker ? reservedValidList4_33 : _GEN_8175; // @[decode.scala 431:29 330:31]
  wire  _GEN_8496 = 3'h2 == branchTracker ? reservedValidList4_34 : _GEN_8176; // @[decode.scala 431:29 330:31]
  wire  _GEN_8497 = 3'h2 == branchTracker ? reservedValidList4_35 : _GEN_8177; // @[decode.scala 431:29 330:31]
  wire  _GEN_8498 = 3'h2 == branchTracker ? reservedValidList4_36 : _GEN_8178; // @[decode.scala 431:29 330:31]
  wire  _GEN_8499 = 3'h2 == branchTracker ? reservedValidList4_37 : _GEN_8179; // @[decode.scala 431:29 330:31]
  wire  _GEN_8500 = 3'h2 == branchTracker ? reservedValidList4_38 : _GEN_8180; // @[decode.scala 431:29 330:31]
  wire  _GEN_8501 = 3'h2 == branchTracker ? reservedValidList4_39 : _GEN_8181; // @[decode.scala 431:29 330:31]
  wire  _GEN_8502 = 3'h2 == branchTracker ? reservedValidList4_40 : _GEN_8182; // @[decode.scala 431:29 330:31]
  wire  _GEN_8503 = 3'h2 == branchTracker ? reservedValidList4_41 : _GEN_8183; // @[decode.scala 431:29 330:31]
  wire  _GEN_8504 = 3'h2 == branchTracker ? reservedValidList4_42 : _GEN_8184; // @[decode.scala 431:29 330:31]
  wire  _GEN_8505 = 3'h2 == branchTracker ? reservedValidList4_43 : _GEN_8185; // @[decode.scala 431:29 330:31]
  wire  _GEN_8506 = 3'h2 == branchTracker ? reservedValidList4_44 : _GEN_8186; // @[decode.scala 431:29 330:31]
  wire  _GEN_8507 = 3'h2 == branchTracker ? reservedValidList4_45 : _GEN_8187; // @[decode.scala 431:29 330:31]
  wire  _GEN_8508 = 3'h2 == branchTracker ? reservedValidList4_46 : _GEN_8188; // @[decode.scala 431:29 330:31]
  wire  _GEN_8509 = 3'h2 == branchTracker ? reservedValidList4_47 : _GEN_8189; // @[decode.scala 431:29 330:31]
  wire  _GEN_8510 = 3'h2 == branchTracker ? reservedValidList4_48 : _GEN_8190; // @[decode.scala 431:29 330:31]
  wire  _GEN_8511 = 3'h2 == branchTracker ? reservedValidList4_49 : _GEN_8191; // @[decode.scala 431:29 330:31]
  wire  _GEN_8512 = 3'h2 == branchTracker ? reservedValidList4_50 : _GEN_8192; // @[decode.scala 431:29 330:31]
  wire  _GEN_8513 = 3'h2 == branchTracker ? reservedValidList4_51 : _GEN_8193; // @[decode.scala 431:29 330:31]
  wire  _GEN_8514 = 3'h2 == branchTracker ? reservedValidList4_52 : _GEN_8194; // @[decode.scala 431:29 330:31]
  wire  _GEN_8515 = 3'h2 == branchTracker ? reservedValidList4_53 : _GEN_8195; // @[decode.scala 431:29 330:31]
  wire  _GEN_8516 = 3'h2 == branchTracker ? reservedValidList4_54 : _GEN_8196; // @[decode.scala 431:29 330:31]
  wire  _GEN_8517 = 3'h2 == branchTracker ? reservedValidList4_55 : _GEN_8197; // @[decode.scala 431:29 330:31]
  wire  _GEN_8518 = 3'h2 == branchTracker ? reservedValidList4_56 : _GEN_8198; // @[decode.scala 431:29 330:31]
  wire  _GEN_8519 = 3'h2 == branchTracker ? reservedValidList4_57 : _GEN_8199; // @[decode.scala 431:29 330:31]
  wire  _GEN_8520 = 3'h2 == branchTracker ? reservedValidList4_58 : _GEN_8200; // @[decode.scala 431:29 330:31]
  wire  _GEN_8521 = 3'h2 == branchTracker ? reservedValidList4_59 : _GEN_8201; // @[decode.scala 431:29 330:31]
  wire  _GEN_8522 = 3'h2 == branchTracker ? reservedValidList4_60 : _GEN_8202; // @[decode.scala 431:29 330:31]
  wire  _GEN_8523 = 3'h2 == branchTracker ? reservedValidList4_61 : _GEN_8203; // @[decode.scala 431:29 330:31]
  wire  _GEN_8524 = 3'h2 == branchTracker ? reservedValidList4_62 : _GEN_8204; // @[decode.scala 431:29 330:31]
  wire  _GEN_8525 = 3'h2 == branchTracker ? reservedValidList4_63 : _GEN_8205; // @[decode.scala 431:29 330:31]
  wire  _GEN_8558 = 3'h1 == branchTracker ? _GEN_6958 : _GEN_6437; // @[decode.scala 431:29]
  wire  _GEN_8559 = 3'h1 == branchTracker ? _GEN_6959 : _GEN_6438; // @[decode.scala 431:29]
  wire  _GEN_8560 = 3'h1 == branchTracker ? _GEN_6960 : _GEN_6439; // @[decode.scala 431:29]
  wire  _GEN_8561 = 3'h1 == branchTracker ? _GEN_6961 : _GEN_6440; // @[decode.scala 431:29]
  wire  _GEN_8562 = 3'h1 == branchTracker ? _GEN_6962 : _GEN_6441; // @[decode.scala 431:29]
  wire  _GEN_8563 = 3'h1 == branchTracker ? _GEN_6963 : _GEN_6442; // @[decode.scala 431:29]
  wire  _GEN_8564 = 3'h1 == branchTracker ? _GEN_6964 : _GEN_6443; // @[decode.scala 431:29]
  wire  _GEN_8565 = 3'h1 == branchTracker ? _GEN_6965 : _GEN_6444; // @[decode.scala 431:29]
  wire  _GEN_8566 = 3'h1 == branchTracker ? _GEN_6966 : _GEN_6445; // @[decode.scala 431:29]
  wire  _GEN_8567 = 3'h1 == branchTracker ? _GEN_6967 : _GEN_6446; // @[decode.scala 431:29]
  wire  _GEN_8568 = 3'h1 == branchTracker ? _GEN_6968 : _GEN_6447; // @[decode.scala 431:29]
  wire  _GEN_8569 = 3'h1 == branchTracker ? _GEN_6969 : _GEN_6448; // @[decode.scala 431:29]
  wire  _GEN_8570 = 3'h1 == branchTracker ? _GEN_6970 : _GEN_6449; // @[decode.scala 431:29]
  wire  _GEN_8571 = 3'h1 == branchTracker ? _GEN_6971 : _GEN_6450; // @[decode.scala 431:29]
  wire  _GEN_8572 = 3'h1 == branchTracker ? _GEN_6972 : _GEN_6451; // @[decode.scala 431:29]
  wire  _GEN_8573 = 3'h1 == branchTracker ? _GEN_6973 : _GEN_6452; // @[decode.scala 431:29]
  wire  _GEN_8574 = 3'h1 == branchTracker ? _GEN_6974 : _GEN_6453; // @[decode.scala 431:29]
  wire  _GEN_8575 = 3'h1 == branchTracker ? _GEN_6975 : _GEN_6454; // @[decode.scala 431:29]
  wire  _GEN_8576 = 3'h1 == branchTracker ? _GEN_6976 : _GEN_6455; // @[decode.scala 431:29]
  wire  _GEN_8577 = 3'h1 == branchTracker ? _GEN_6977 : _GEN_6456; // @[decode.scala 431:29]
  wire  _GEN_8578 = 3'h1 == branchTracker ? _GEN_6978 : _GEN_6457; // @[decode.scala 431:29]
  wire  _GEN_8579 = 3'h1 == branchTracker ? _GEN_6979 : _GEN_6458; // @[decode.scala 431:29]
  wire  _GEN_8580 = 3'h1 == branchTracker ? _GEN_6980 : _GEN_6459; // @[decode.scala 431:29]
  wire  _GEN_8581 = 3'h1 == branchTracker ? _GEN_6981 : _GEN_6460; // @[decode.scala 431:29]
  wire  _GEN_8582 = 3'h1 == branchTracker ? _GEN_6982 : _GEN_6461; // @[decode.scala 431:29]
  wire  _GEN_8583 = 3'h1 == branchTracker ? _GEN_6983 : _GEN_6462; // @[decode.scala 431:29]
  wire  _GEN_8584 = 3'h1 == branchTracker ? _GEN_6984 : _GEN_6463; // @[decode.scala 431:29]
  wire  _GEN_8585 = 3'h1 == branchTracker ? _GEN_6985 : _GEN_6464; // @[decode.scala 431:29]
  wire  _GEN_8586 = 3'h1 == branchTracker ? _GEN_6986 : _GEN_6465; // @[decode.scala 431:29]
  wire  _GEN_8587 = 3'h1 == branchTracker ? _GEN_6987 : _GEN_6466; // @[decode.scala 431:29]
  wire  _GEN_8588 = 3'h1 == branchTracker ? _GEN_6988 : _GEN_6467; // @[decode.scala 431:29]
  wire  _GEN_8589 = 3'h1 == branchTracker ? _GEN_6989 : _GEN_6468; // @[decode.scala 431:29]
  wire  _GEN_8590 = 3'h1 == branchTracker ? _GEN_6990 : _GEN_6469; // @[decode.scala 431:29]
  wire  _GEN_8591 = 3'h1 == branchTracker ? _GEN_6991 : _GEN_6470; // @[decode.scala 431:29]
  wire  _GEN_8592 = 3'h1 == branchTracker ? _GEN_6992 : _GEN_6471; // @[decode.scala 431:29]
  wire  _GEN_8593 = 3'h1 == branchTracker ? _GEN_6993 : _GEN_6472; // @[decode.scala 431:29]
  wire  _GEN_8594 = 3'h1 == branchTracker ? _GEN_6994 : _GEN_6473; // @[decode.scala 431:29]
  wire  _GEN_8595 = 3'h1 == branchTracker ? _GEN_6995 : _GEN_6474; // @[decode.scala 431:29]
  wire  _GEN_8596 = 3'h1 == branchTracker ? _GEN_6996 : _GEN_6475; // @[decode.scala 431:29]
  wire  _GEN_8597 = 3'h1 == branchTracker ? _GEN_6997 : _GEN_6476; // @[decode.scala 431:29]
  wire  _GEN_8598 = 3'h1 == branchTracker ? _GEN_6998 : _GEN_6477; // @[decode.scala 431:29]
  wire  _GEN_8599 = 3'h1 == branchTracker ? _GEN_6999 : _GEN_6478; // @[decode.scala 431:29]
  wire  _GEN_8600 = 3'h1 == branchTracker ? _GEN_7000 : _GEN_6479; // @[decode.scala 431:29]
  wire  _GEN_8601 = 3'h1 == branchTracker ? _GEN_7001 : _GEN_6480; // @[decode.scala 431:29]
  wire  _GEN_8602 = 3'h1 == branchTracker ? _GEN_7002 : _GEN_6481; // @[decode.scala 431:29]
  wire  _GEN_8603 = 3'h1 == branchTracker ? _GEN_7003 : _GEN_6482; // @[decode.scala 431:29]
  wire  _GEN_8604 = 3'h1 == branchTracker ? _GEN_7004 : _GEN_6483; // @[decode.scala 431:29]
  wire  _GEN_8605 = 3'h1 == branchTracker ? _GEN_7005 : _GEN_6484; // @[decode.scala 431:29]
  wire  _GEN_8606 = 3'h1 == branchTracker ? _GEN_7006 : _GEN_6485; // @[decode.scala 431:29]
  wire  _GEN_8607 = 3'h1 == branchTracker ? _GEN_7007 : _GEN_6486; // @[decode.scala 431:29]
  wire  _GEN_8608 = 3'h1 == branchTracker ? _GEN_7008 : _GEN_6487; // @[decode.scala 431:29]
  wire  _GEN_8609 = 3'h1 == branchTracker ? _GEN_7009 : _GEN_6488; // @[decode.scala 431:29]
  wire  _GEN_8610 = 3'h1 == branchTracker ? _GEN_7010 : _GEN_6489; // @[decode.scala 431:29]
  wire  _GEN_8611 = 3'h1 == branchTracker ? _GEN_7011 : _GEN_6490; // @[decode.scala 431:29]
  wire  _GEN_8612 = 3'h1 == branchTracker ? _GEN_7012 : _GEN_6491; // @[decode.scala 431:29]
  wire  _GEN_8613 = 3'h1 == branchTracker ? _GEN_7013 : _GEN_6492; // @[decode.scala 431:29]
  wire  _GEN_8614 = 3'h1 == branchTracker ? _GEN_7014 : _GEN_6493; // @[decode.scala 431:29]
  wire  _GEN_8615 = 3'h1 == branchTracker ? _GEN_7015 : _GEN_6494; // @[decode.scala 431:29]
  wire  _GEN_8616 = 3'h1 == branchTracker ? _GEN_7016 : _GEN_6495; // @[decode.scala 431:29]
  wire  _GEN_8617 = 3'h1 == branchTracker ? _GEN_7017 : _GEN_6496; // @[decode.scala 431:29]
  wire  _GEN_8618 = 3'h1 == branchTracker ? _GEN_7018 : _GEN_6497; // @[decode.scala 431:29]
  wire  _GEN_8619 = 3'h1 == branchTracker ? _GEN_7019 : _GEN_6498; // @[decode.scala 431:29]
  wire  _GEN_8620 = 3'h1 == branchTracker ? _GEN_7020 : _GEN_6499; // @[decode.scala 431:29]
  wire  _GEN_8718 = 3'h1 == branchTracker ? _GEN_6501 : _GEN_8238; // @[decode.scala 431:29]
  wire  _GEN_8719 = 3'h1 == branchTracker ? _GEN_6502 : _GEN_8239; // @[decode.scala 431:29]
  wire  _GEN_8720 = 3'h1 == branchTracker ? _GEN_6503 : _GEN_8240; // @[decode.scala 431:29]
  wire  _GEN_8721 = 3'h1 == branchTracker ? _GEN_6504 : _GEN_8241; // @[decode.scala 431:29]
  wire  _GEN_8722 = 3'h1 == branchTracker ? _GEN_6505 : _GEN_8242; // @[decode.scala 431:29]
  wire  _GEN_8723 = 3'h1 == branchTracker ? _GEN_6506 : _GEN_8243; // @[decode.scala 431:29]
  wire  _GEN_8724 = 3'h1 == branchTracker ? _GEN_6507 : _GEN_8244; // @[decode.scala 431:29]
  wire  _GEN_8725 = 3'h1 == branchTracker ? _GEN_6508 : _GEN_8245; // @[decode.scala 431:29]
  wire  _GEN_8726 = 3'h1 == branchTracker ? _GEN_6509 : _GEN_8246; // @[decode.scala 431:29]
  wire  _GEN_8727 = 3'h1 == branchTracker ? _GEN_6510 : _GEN_8247; // @[decode.scala 431:29]
  wire  _GEN_8728 = 3'h1 == branchTracker ? _GEN_6511 : _GEN_8248; // @[decode.scala 431:29]
  wire  _GEN_8729 = 3'h1 == branchTracker ? _GEN_6512 : _GEN_8249; // @[decode.scala 431:29]
  wire  _GEN_8730 = 3'h1 == branchTracker ? _GEN_6513 : _GEN_8250; // @[decode.scala 431:29]
  wire  _GEN_8731 = 3'h1 == branchTracker ? _GEN_6514 : _GEN_8251; // @[decode.scala 431:29]
  wire  _GEN_8732 = 3'h1 == branchTracker ? _GEN_6515 : _GEN_8252; // @[decode.scala 431:29]
  wire  _GEN_8733 = 3'h1 == branchTracker ? _GEN_6516 : _GEN_8253; // @[decode.scala 431:29]
  wire  _GEN_8734 = 3'h1 == branchTracker ? _GEN_6517 : _GEN_8254; // @[decode.scala 431:29]
  wire  _GEN_8735 = 3'h1 == branchTracker ? _GEN_6518 : _GEN_8255; // @[decode.scala 431:29]
  wire  _GEN_8736 = 3'h1 == branchTracker ? _GEN_6519 : _GEN_8256; // @[decode.scala 431:29]
  wire  _GEN_8737 = 3'h1 == branchTracker ? _GEN_6520 : _GEN_8257; // @[decode.scala 431:29]
  wire  _GEN_8738 = 3'h1 == branchTracker ? _GEN_6521 : _GEN_8258; // @[decode.scala 431:29]
  wire  _GEN_8739 = 3'h1 == branchTracker ? _GEN_6522 : _GEN_8259; // @[decode.scala 431:29]
  wire  _GEN_8740 = 3'h1 == branchTracker ? _GEN_6523 : _GEN_8260; // @[decode.scala 431:29]
  wire  _GEN_8741 = 3'h1 == branchTracker ? _GEN_6524 : _GEN_8261; // @[decode.scala 431:29]
  wire  _GEN_8742 = 3'h1 == branchTracker ? _GEN_6525 : _GEN_8262; // @[decode.scala 431:29]
  wire  _GEN_8743 = 3'h1 == branchTracker ? _GEN_6526 : _GEN_8263; // @[decode.scala 431:29]
  wire  _GEN_8744 = 3'h1 == branchTracker ? _GEN_6527 : _GEN_8264; // @[decode.scala 431:29]
  wire  _GEN_8745 = 3'h1 == branchTracker ? _GEN_6528 : _GEN_8265; // @[decode.scala 431:29]
  wire  _GEN_8746 = 3'h1 == branchTracker ? _GEN_6529 : _GEN_8266; // @[decode.scala 431:29]
  wire  _GEN_8747 = 3'h1 == branchTracker ? _GEN_6530 : _GEN_8267; // @[decode.scala 431:29]
  wire  _GEN_8748 = 3'h1 == branchTracker ? _GEN_6531 : _GEN_8268; // @[decode.scala 431:29]
  wire  _GEN_8749 = 3'h1 == branchTracker ? _GEN_6532 : _GEN_8269; // @[decode.scala 431:29]
  wire  _GEN_8750 = 3'h1 == branchTracker ? _GEN_6533 : _GEN_8270; // @[decode.scala 431:29]
  wire  _GEN_8751 = 3'h1 == branchTracker ? _GEN_6534 : _GEN_8271; // @[decode.scala 431:29]
  wire  _GEN_8752 = 3'h1 == branchTracker ? _GEN_6535 : _GEN_8272; // @[decode.scala 431:29]
  wire  _GEN_8753 = 3'h1 == branchTracker ? _GEN_6536 : _GEN_8273; // @[decode.scala 431:29]
  wire  _GEN_8754 = 3'h1 == branchTracker ? _GEN_6537 : _GEN_8274; // @[decode.scala 431:29]
  wire  _GEN_8755 = 3'h1 == branchTracker ? _GEN_6538 : _GEN_8275; // @[decode.scala 431:29]
  wire  _GEN_8756 = 3'h1 == branchTracker ? _GEN_6539 : _GEN_8276; // @[decode.scala 431:29]
  wire  _GEN_8757 = 3'h1 == branchTracker ? _GEN_6540 : _GEN_8277; // @[decode.scala 431:29]
  wire  _GEN_8758 = 3'h1 == branchTracker ? _GEN_6541 : _GEN_8278; // @[decode.scala 431:29]
  wire  _GEN_8759 = 3'h1 == branchTracker ? _GEN_6542 : _GEN_8279; // @[decode.scala 431:29]
  wire  _GEN_8760 = 3'h1 == branchTracker ? _GEN_6543 : _GEN_8280; // @[decode.scala 431:29]
  wire  _GEN_8761 = 3'h1 == branchTracker ? _GEN_6544 : _GEN_8281; // @[decode.scala 431:29]
  wire  _GEN_8762 = 3'h1 == branchTracker ? _GEN_6545 : _GEN_8282; // @[decode.scala 431:29]
  wire  _GEN_8763 = 3'h1 == branchTracker ? _GEN_6546 : _GEN_8283; // @[decode.scala 431:29]
  wire  _GEN_8764 = 3'h1 == branchTracker ? _GEN_6547 : _GEN_8284; // @[decode.scala 431:29]
  wire  _GEN_8765 = 3'h1 == branchTracker ? _GEN_6548 : _GEN_8285; // @[decode.scala 431:29]
  wire  _GEN_8766 = 3'h1 == branchTracker ? _GEN_6549 : _GEN_8286; // @[decode.scala 431:29]
  wire  _GEN_8767 = 3'h1 == branchTracker ? _GEN_6550 : _GEN_8287; // @[decode.scala 431:29]
  wire  _GEN_8768 = 3'h1 == branchTracker ? _GEN_6551 : _GEN_8288; // @[decode.scala 431:29]
  wire  _GEN_8769 = 3'h1 == branchTracker ? _GEN_6552 : _GEN_8289; // @[decode.scala 431:29]
  wire  _GEN_8770 = 3'h1 == branchTracker ? _GEN_6553 : _GEN_8290; // @[decode.scala 431:29]
  wire  _GEN_8771 = 3'h1 == branchTracker ? _GEN_6554 : _GEN_8291; // @[decode.scala 431:29]
  wire  _GEN_8772 = 3'h1 == branchTracker ? _GEN_6555 : _GEN_8292; // @[decode.scala 431:29]
  wire  _GEN_8773 = 3'h1 == branchTracker ? _GEN_6556 : _GEN_8293; // @[decode.scala 431:29]
  wire  _GEN_8774 = 3'h1 == branchTracker ? _GEN_6557 : _GEN_8294; // @[decode.scala 431:29]
  wire  _GEN_8775 = 3'h1 == branchTracker ? _GEN_6558 : _GEN_8295; // @[decode.scala 431:29]
  wire  _GEN_8776 = 3'h1 == branchTracker ? _GEN_6559 : _GEN_8296; // @[decode.scala 431:29]
  wire  _GEN_8777 = 3'h1 == branchTracker ? _GEN_6560 : _GEN_8297; // @[decode.scala 431:29]
  wire  _GEN_8778 = 3'h1 == branchTracker ? _GEN_6561 : _GEN_8298; // @[decode.scala 431:29]
  wire  _GEN_8779 = 3'h1 == branchTracker ? _GEN_6562 : _GEN_8299; // @[decode.scala 431:29]
  wire  _GEN_8780 = 3'h1 == branchTracker ? _GEN_6563 : _GEN_8300; // @[decode.scala 431:29]
  wire  _GEN_8878 = 3'h1 == branchTracker ? reservedFreeList4_0 : _GEN_8398; // @[decode.scala 431:29 325:30]
  wire  _GEN_8879 = 3'h1 == branchTracker ? reservedFreeList4_1 : _GEN_8399; // @[decode.scala 431:29 325:30]
  wire  _GEN_8880 = 3'h1 == branchTracker ? reservedFreeList4_2 : _GEN_8400; // @[decode.scala 431:29 325:30]
  wire  _GEN_8881 = 3'h1 == branchTracker ? reservedFreeList4_3 : _GEN_8401; // @[decode.scala 431:29 325:30]
  wire  _GEN_8882 = 3'h1 == branchTracker ? reservedFreeList4_4 : _GEN_8402; // @[decode.scala 431:29 325:30]
  wire  _GEN_8883 = 3'h1 == branchTracker ? reservedFreeList4_5 : _GEN_8403; // @[decode.scala 431:29 325:30]
  wire  _GEN_8884 = 3'h1 == branchTracker ? reservedFreeList4_6 : _GEN_8404; // @[decode.scala 431:29 325:30]
  wire  _GEN_8885 = 3'h1 == branchTracker ? reservedFreeList4_7 : _GEN_8405; // @[decode.scala 431:29 325:30]
  wire  _GEN_8886 = 3'h1 == branchTracker ? reservedFreeList4_8 : _GEN_8406; // @[decode.scala 431:29 325:30]
  wire  _GEN_8887 = 3'h1 == branchTracker ? reservedFreeList4_9 : _GEN_8407; // @[decode.scala 431:29 325:30]
  wire  _GEN_8888 = 3'h1 == branchTracker ? reservedFreeList4_10 : _GEN_8408; // @[decode.scala 431:29 325:30]
  wire  _GEN_8889 = 3'h1 == branchTracker ? reservedFreeList4_11 : _GEN_8409; // @[decode.scala 431:29 325:30]
  wire  _GEN_8890 = 3'h1 == branchTracker ? reservedFreeList4_12 : _GEN_8410; // @[decode.scala 431:29 325:30]
  wire  _GEN_8891 = 3'h1 == branchTracker ? reservedFreeList4_13 : _GEN_8411; // @[decode.scala 431:29 325:30]
  wire  _GEN_8892 = 3'h1 == branchTracker ? reservedFreeList4_14 : _GEN_8412; // @[decode.scala 431:29 325:30]
  wire  _GEN_8893 = 3'h1 == branchTracker ? reservedFreeList4_15 : _GEN_8413; // @[decode.scala 431:29 325:30]
  wire  _GEN_8894 = 3'h1 == branchTracker ? reservedFreeList4_16 : _GEN_8414; // @[decode.scala 431:29 325:30]
  wire  _GEN_8895 = 3'h1 == branchTracker ? reservedFreeList4_17 : _GEN_8415; // @[decode.scala 431:29 325:30]
  wire  _GEN_8896 = 3'h1 == branchTracker ? reservedFreeList4_18 : _GEN_8416; // @[decode.scala 431:29 325:30]
  wire  _GEN_8897 = 3'h1 == branchTracker ? reservedFreeList4_19 : _GEN_8417; // @[decode.scala 431:29 325:30]
  wire  _GEN_8898 = 3'h1 == branchTracker ? reservedFreeList4_20 : _GEN_8418; // @[decode.scala 431:29 325:30]
  wire  _GEN_8899 = 3'h1 == branchTracker ? reservedFreeList4_21 : _GEN_8419; // @[decode.scala 431:29 325:30]
  wire  _GEN_8900 = 3'h1 == branchTracker ? reservedFreeList4_22 : _GEN_8420; // @[decode.scala 431:29 325:30]
  wire  _GEN_8901 = 3'h1 == branchTracker ? reservedFreeList4_23 : _GEN_8421; // @[decode.scala 431:29 325:30]
  wire  _GEN_8902 = 3'h1 == branchTracker ? reservedFreeList4_24 : _GEN_8422; // @[decode.scala 431:29 325:30]
  wire  _GEN_8903 = 3'h1 == branchTracker ? reservedFreeList4_25 : _GEN_8423; // @[decode.scala 431:29 325:30]
  wire  _GEN_8904 = 3'h1 == branchTracker ? reservedFreeList4_26 : _GEN_8424; // @[decode.scala 431:29 325:30]
  wire  _GEN_8905 = 3'h1 == branchTracker ? reservedFreeList4_27 : _GEN_8425; // @[decode.scala 431:29 325:30]
  wire  _GEN_8906 = 3'h1 == branchTracker ? reservedFreeList4_28 : _GEN_8426; // @[decode.scala 431:29 325:30]
  wire  _GEN_8907 = 3'h1 == branchTracker ? reservedFreeList4_29 : _GEN_8427; // @[decode.scala 431:29 325:30]
  wire  _GEN_8908 = 3'h1 == branchTracker ? reservedFreeList4_30 : _GEN_8428; // @[decode.scala 431:29 325:30]
  wire  _GEN_8909 = 3'h1 == branchTracker ? reservedFreeList4_31 : _GEN_8429; // @[decode.scala 431:29 325:30]
  wire  _GEN_8910 = 3'h1 == branchTracker ? reservedFreeList4_32 : _GEN_8430; // @[decode.scala 431:29 325:30]
  wire  _GEN_8911 = 3'h1 == branchTracker ? reservedFreeList4_33 : _GEN_8431; // @[decode.scala 431:29 325:30]
  wire  _GEN_8912 = 3'h1 == branchTracker ? reservedFreeList4_34 : _GEN_8432; // @[decode.scala 431:29 325:30]
  wire  _GEN_8913 = 3'h1 == branchTracker ? reservedFreeList4_35 : _GEN_8433; // @[decode.scala 431:29 325:30]
  wire  _GEN_8914 = 3'h1 == branchTracker ? reservedFreeList4_36 : _GEN_8434; // @[decode.scala 431:29 325:30]
  wire  _GEN_8915 = 3'h1 == branchTracker ? reservedFreeList4_37 : _GEN_8435; // @[decode.scala 431:29 325:30]
  wire  _GEN_8916 = 3'h1 == branchTracker ? reservedFreeList4_38 : _GEN_8436; // @[decode.scala 431:29 325:30]
  wire  _GEN_8917 = 3'h1 == branchTracker ? reservedFreeList4_39 : _GEN_8437; // @[decode.scala 431:29 325:30]
  wire  _GEN_8918 = 3'h1 == branchTracker ? reservedFreeList4_40 : _GEN_8438; // @[decode.scala 431:29 325:30]
  wire  _GEN_8919 = 3'h1 == branchTracker ? reservedFreeList4_41 : _GEN_8439; // @[decode.scala 431:29 325:30]
  wire  _GEN_8920 = 3'h1 == branchTracker ? reservedFreeList4_42 : _GEN_8440; // @[decode.scala 431:29 325:30]
  wire  _GEN_8921 = 3'h1 == branchTracker ? reservedFreeList4_43 : _GEN_8441; // @[decode.scala 431:29 325:30]
  wire  _GEN_8922 = 3'h1 == branchTracker ? reservedFreeList4_44 : _GEN_8442; // @[decode.scala 431:29 325:30]
  wire  _GEN_8923 = 3'h1 == branchTracker ? reservedFreeList4_45 : _GEN_8443; // @[decode.scala 431:29 325:30]
  wire  _GEN_8924 = 3'h1 == branchTracker ? reservedFreeList4_46 : _GEN_8444; // @[decode.scala 431:29 325:30]
  wire  _GEN_8925 = 3'h1 == branchTracker ? reservedFreeList4_47 : _GEN_8445; // @[decode.scala 431:29 325:30]
  wire  _GEN_8926 = 3'h1 == branchTracker ? reservedFreeList4_48 : _GEN_8446; // @[decode.scala 431:29 325:30]
  wire  _GEN_8927 = 3'h1 == branchTracker ? reservedFreeList4_49 : _GEN_8447; // @[decode.scala 431:29 325:30]
  wire  _GEN_8928 = 3'h1 == branchTracker ? reservedFreeList4_50 : _GEN_8448; // @[decode.scala 431:29 325:30]
  wire  _GEN_8929 = 3'h1 == branchTracker ? reservedFreeList4_51 : _GEN_8449; // @[decode.scala 431:29 325:30]
  wire  _GEN_8930 = 3'h1 == branchTracker ? reservedFreeList4_52 : _GEN_8450; // @[decode.scala 431:29 325:30]
  wire  _GEN_8931 = 3'h1 == branchTracker ? reservedFreeList4_53 : _GEN_8451; // @[decode.scala 431:29 325:30]
  wire  _GEN_8932 = 3'h1 == branchTracker ? reservedFreeList4_54 : _GEN_8452; // @[decode.scala 431:29 325:30]
  wire  _GEN_8933 = 3'h1 == branchTracker ? reservedFreeList4_55 : _GEN_8453; // @[decode.scala 431:29 325:30]
  wire  _GEN_8934 = 3'h1 == branchTracker ? reservedFreeList4_56 : _GEN_8454; // @[decode.scala 431:29 325:30]
  wire  _GEN_8935 = 3'h1 == branchTracker ? reservedFreeList4_57 : _GEN_8455; // @[decode.scala 431:29 325:30]
  wire  _GEN_8936 = 3'h1 == branchTracker ? reservedFreeList4_58 : _GEN_8456; // @[decode.scala 431:29 325:30]
  wire  _GEN_8937 = 3'h1 == branchTracker ? reservedFreeList4_59 : _GEN_8457; // @[decode.scala 431:29 325:30]
  wire  _GEN_8938 = 3'h1 == branchTracker ? reservedFreeList4_60 : _GEN_8458; // @[decode.scala 431:29 325:30]
  wire  _GEN_8939 = 3'h1 == branchTracker ? reservedFreeList4_61 : _GEN_8459; // @[decode.scala 431:29 325:30]
  wire  _GEN_8940 = 3'h1 == branchTracker ? reservedFreeList4_62 : _GEN_8460; // @[decode.scala 431:29 325:30]
  wire  _GEN_9038 = 3'h0 == branchTracker ? _GEN_6958 : _GEN_6373; // @[decode.scala 431:29]
  wire  _GEN_9039 = 3'h0 == branchTracker ? _GEN_6959 : _GEN_6374; // @[decode.scala 431:29]
  wire  _GEN_9040 = 3'h0 == branchTracker ? _GEN_6960 : _GEN_6375; // @[decode.scala 431:29]
  wire  _GEN_9041 = 3'h0 == branchTracker ? _GEN_6961 : _GEN_6376; // @[decode.scala 431:29]
  wire  _GEN_9042 = 3'h0 == branchTracker ? _GEN_6962 : _GEN_6377; // @[decode.scala 431:29]
  wire  _GEN_9043 = 3'h0 == branchTracker ? _GEN_6963 : _GEN_6378; // @[decode.scala 431:29]
  wire  _GEN_9044 = 3'h0 == branchTracker ? _GEN_6964 : _GEN_6379; // @[decode.scala 431:29]
  wire  _GEN_9045 = 3'h0 == branchTracker ? _GEN_6965 : _GEN_6380; // @[decode.scala 431:29]
  wire  _GEN_9046 = 3'h0 == branchTracker ? _GEN_6966 : _GEN_6381; // @[decode.scala 431:29]
  wire  _GEN_9047 = 3'h0 == branchTracker ? _GEN_6967 : _GEN_6382; // @[decode.scala 431:29]
  wire  _GEN_9048 = 3'h0 == branchTracker ? _GEN_6968 : _GEN_6383; // @[decode.scala 431:29]
  wire  _GEN_9049 = 3'h0 == branchTracker ? _GEN_6969 : _GEN_6384; // @[decode.scala 431:29]
  wire  _GEN_9050 = 3'h0 == branchTracker ? _GEN_6970 : _GEN_6385; // @[decode.scala 431:29]
  wire  _GEN_9051 = 3'h0 == branchTracker ? _GEN_6971 : _GEN_6386; // @[decode.scala 431:29]
  wire  _GEN_9052 = 3'h0 == branchTracker ? _GEN_6972 : _GEN_6387; // @[decode.scala 431:29]
  wire  _GEN_9053 = 3'h0 == branchTracker ? _GEN_6973 : _GEN_6388; // @[decode.scala 431:29]
  wire  _GEN_9054 = 3'h0 == branchTracker ? _GEN_6974 : _GEN_6389; // @[decode.scala 431:29]
  wire  _GEN_9055 = 3'h0 == branchTracker ? _GEN_6975 : _GEN_6390; // @[decode.scala 431:29]
  wire  _GEN_9056 = 3'h0 == branchTracker ? _GEN_6976 : _GEN_6391; // @[decode.scala 431:29]
  wire  _GEN_9057 = 3'h0 == branchTracker ? _GEN_6977 : _GEN_6392; // @[decode.scala 431:29]
  wire  _GEN_9058 = 3'h0 == branchTracker ? _GEN_6978 : _GEN_6393; // @[decode.scala 431:29]
  wire  _GEN_9059 = 3'h0 == branchTracker ? _GEN_6979 : _GEN_6394; // @[decode.scala 431:29]
  wire  _GEN_9060 = 3'h0 == branchTracker ? _GEN_6980 : _GEN_6395; // @[decode.scala 431:29]
  wire  _GEN_9061 = 3'h0 == branchTracker ? _GEN_6981 : _GEN_6396; // @[decode.scala 431:29]
  wire  _GEN_9062 = 3'h0 == branchTracker ? _GEN_6982 : _GEN_6397; // @[decode.scala 431:29]
  wire  _GEN_9063 = 3'h0 == branchTracker ? _GEN_6983 : _GEN_6398; // @[decode.scala 431:29]
  wire  _GEN_9064 = 3'h0 == branchTracker ? _GEN_6984 : _GEN_6399; // @[decode.scala 431:29]
  wire  _GEN_9065 = 3'h0 == branchTracker ? _GEN_6985 : _GEN_6400; // @[decode.scala 431:29]
  wire  _GEN_9066 = 3'h0 == branchTracker ? _GEN_6986 : _GEN_6401; // @[decode.scala 431:29]
  wire  _GEN_9067 = 3'h0 == branchTracker ? _GEN_6987 : _GEN_6402; // @[decode.scala 431:29]
  wire  _GEN_9068 = 3'h0 == branchTracker ? _GEN_6988 : _GEN_6403; // @[decode.scala 431:29]
  wire  _GEN_9069 = 3'h0 == branchTracker ? _GEN_6989 : _GEN_6404; // @[decode.scala 431:29]
  wire  _GEN_9070 = 3'h0 == branchTracker ? _GEN_6990 : _GEN_6405; // @[decode.scala 431:29]
  wire  _GEN_9071 = 3'h0 == branchTracker ? _GEN_6991 : _GEN_6406; // @[decode.scala 431:29]
  wire  _GEN_9072 = 3'h0 == branchTracker ? _GEN_6992 : _GEN_6407; // @[decode.scala 431:29]
  wire  _GEN_9073 = 3'h0 == branchTracker ? _GEN_6993 : _GEN_6408; // @[decode.scala 431:29]
  wire  _GEN_9074 = 3'h0 == branchTracker ? _GEN_6994 : _GEN_6409; // @[decode.scala 431:29]
  wire  _GEN_9075 = 3'h0 == branchTracker ? _GEN_6995 : _GEN_6410; // @[decode.scala 431:29]
  wire  _GEN_9076 = 3'h0 == branchTracker ? _GEN_6996 : _GEN_6411; // @[decode.scala 431:29]
  wire  _GEN_9077 = 3'h0 == branchTracker ? _GEN_6997 : _GEN_6412; // @[decode.scala 431:29]
  wire  _GEN_9078 = 3'h0 == branchTracker ? _GEN_6998 : _GEN_6413; // @[decode.scala 431:29]
  wire  _GEN_9079 = 3'h0 == branchTracker ? _GEN_6999 : _GEN_6414; // @[decode.scala 431:29]
  wire  _GEN_9080 = 3'h0 == branchTracker ? _GEN_7000 : _GEN_6415; // @[decode.scala 431:29]
  wire  _GEN_9081 = 3'h0 == branchTracker ? _GEN_7001 : _GEN_6416; // @[decode.scala 431:29]
  wire  _GEN_9082 = 3'h0 == branchTracker ? _GEN_7002 : _GEN_6417; // @[decode.scala 431:29]
  wire  _GEN_9083 = 3'h0 == branchTracker ? _GEN_7003 : _GEN_6418; // @[decode.scala 431:29]
  wire  _GEN_9084 = 3'h0 == branchTracker ? _GEN_7004 : _GEN_6419; // @[decode.scala 431:29]
  wire  _GEN_9085 = 3'h0 == branchTracker ? _GEN_7005 : _GEN_6420; // @[decode.scala 431:29]
  wire  _GEN_9086 = 3'h0 == branchTracker ? _GEN_7006 : _GEN_6421; // @[decode.scala 431:29]
  wire  _GEN_9087 = 3'h0 == branchTracker ? _GEN_7007 : _GEN_6422; // @[decode.scala 431:29]
  wire  _GEN_9088 = 3'h0 == branchTracker ? _GEN_7008 : _GEN_6423; // @[decode.scala 431:29]
  wire  _GEN_9089 = 3'h0 == branchTracker ? _GEN_7009 : _GEN_6424; // @[decode.scala 431:29]
  wire  _GEN_9090 = 3'h0 == branchTracker ? _GEN_7010 : _GEN_6425; // @[decode.scala 431:29]
  wire  _GEN_9091 = 3'h0 == branchTracker ? _GEN_7011 : _GEN_6426; // @[decode.scala 431:29]
  wire  _GEN_9092 = 3'h0 == branchTracker ? _GEN_7012 : _GEN_6427; // @[decode.scala 431:29]
  wire  _GEN_9093 = 3'h0 == branchTracker ? _GEN_7013 : _GEN_6428; // @[decode.scala 431:29]
  wire  _GEN_9094 = 3'h0 == branchTracker ? _GEN_7014 : _GEN_6429; // @[decode.scala 431:29]
  wire  _GEN_9095 = 3'h0 == branchTracker ? _GEN_7015 : _GEN_6430; // @[decode.scala 431:29]
  wire  _GEN_9096 = 3'h0 == branchTracker ? _GEN_7016 : _GEN_6431; // @[decode.scala 431:29]
  wire  _GEN_9097 = 3'h0 == branchTracker ? _GEN_7017 : _GEN_6432; // @[decode.scala 431:29]
  wire  _GEN_9098 = 3'h0 == branchTracker ? _GEN_7018 : _GEN_6433; // @[decode.scala 431:29]
  wire  _GEN_9099 = 3'h0 == branchTracker ? _GEN_7019 : _GEN_6434; // @[decode.scala 431:29]
  wire  _GEN_9100 = 3'h0 == branchTracker ? _GEN_7020 : _GEN_6435; // @[decode.scala 431:29]
  wire  _GEN_9198 = 3'h0 == branchTracker ? _GEN_6437 : _GEN_8558; // @[decode.scala 431:29]
  wire  _GEN_9199 = 3'h0 == branchTracker ? _GEN_6438 : _GEN_8559; // @[decode.scala 431:29]
  wire  _GEN_9200 = 3'h0 == branchTracker ? _GEN_6439 : _GEN_8560; // @[decode.scala 431:29]
  wire  _GEN_9201 = 3'h0 == branchTracker ? _GEN_6440 : _GEN_8561; // @[decode.scala 431:29]
  wire  _GEN_9202 = 3'h0 == branchTracker ? _GEN_6441 : _GEN_8562; // @[decode.scala 431:29]
  wire  _GEN_9203 = 3'h0 == branchTracker ? _GEN_6442 : _GEN_8563; // @[decode.scala 431:29]
  wire  _GEN_9204 = 3'h0 == branchTracker ? _GEN_6443 : _GEN_8564; // @[decode.scala 431:29]
  wire  _GEN_9205 = 3'h0 == branchTracker ? _GEN_6444 : _GEN_8565; // @[decode.scala 431:29]
  wire  _GEN_9206 = 3'h0 == branchTracker ? _GEN_6445 : _GEN_8566; // @[decode.scala 431:29]
  wire  _GEN_9207 = 3'h0 == branchTracker ? _GEN_6446 : _GEN_8567; // @[decode.scala 431:29]
  wire  _GEN_9208 = 3'h0 == branchTracker ? _GEN_6447 : _GEN_8568; // @[decode.scala 431:29]
  wire  _GEN_9209 = 3'h0 == branchTracker ? _GEN_6448 : _GEN_8569; // @[decode.scala 431:29]
  wire  _GEN_9210 = 3'h0 == branchTracker ? _GEN_6449 : _GEN_8570; // @[decode.scala 431:29]
  wire  _GEN_9211 = 3'h0 == branchTracker ? _GEN_6450 : _GEN_8571; // @[decode.scala 431:29]
  wire  _GEN_9212 = 3'h0 == branchTracker ? _GEN_6451 : _GEN_8572; // @[decode.scala 431:29]
  wire  _GEN_9213 = 3'h0 == branchTracker ? _GEN_6452 : _GEN_8573; // @[decode.scala 431:29]
  wire  _GEN_9214 = 3'h0 == branchTracker ? _GEN_6453 : _GEN_8574; // @[decode.scala 431:29]
  wire  _GEN_9215 = 3'h0 == branchTracker ? _GEN_6454 : _GEN_8575; // @[decode.scala 431:29]
  wire  _GEN_9216 = 3'h0 == branchTracker ? _GEN_6455 : _GEN_8576; // @[decode.scala 431:29]
  wire  _GEN_9217 = 3'h0 == branchTracker ? _GEN_6456 : _GEN_8577; // @[decode.scala 431:29]
  wire  _GEN_9218 = 3'h0 == branchTracker ? _GEN_6457 : _GEN_8578; // @[decode.scala 431:29]
  wire  _GEN_9219 = 3'h0 == branchTracker ? _GEN_6458 : _GEN_8579; // @[decode.scala 431:29]
  wire  _GEN_9220 = 3'h0 == branchTracker ? _GEN_6459 : _GEN_8580; // @[decode.scala 431:29]
  wire  _GEN_9221 = 3'h0 == branchTracker ? _GEN_6460 : _GEN_8581; // @[decode.scala 431:29]
  wire  _GEN_9222 = 3'h0 == branchTracker ? _GEN_6461 : _GEN_8582; // @[decode.scala 431:29]
  wire  _GEN_9223 = 3'h0 == branchTracker ? _GEN_6462 : _GEN_8583; // @[decode.scala 431:29]
  wire  _GEN_9224 = 3'h0 == branchTracker ? _GEN_6463 : _GEN_8584; // @[decode.scala 431:29]
  wire  _GEN_9225 = 3'h0 == branchTracker ? _GEN_6464 : _GEN_8585; // @[decode.scala 431:29]
  wire  _GEN_9226 = 3'h0 == branchTracker ? _GEN_6465 : _GEN_8586; // @[decode.scala 431:29]
  wire  _GEN_9227 = 3'h0 == branchTracker ? _GEN_6466 : _GEN_8587; // @[decode.scala 431:29]
  wire  _GEN_9228 = 3'h0 == branchTracker ? _GEN_6467 : _GEN_8588; // @[decode.scala 431:29]
  wire  _GEN_9229 = 3'h0 == branchTracker ? _GEN_6468 : _GEN_8589; // @[decode.scala 431:29]
  wire  _GEN_9230 = 3'h0 == branchTracker ? _GEN_6469 : _GEN_8590; // @[decode.scala 431:29]
  wire  _GEN_9231 = 3'h0 == branchTracker ? _GEN_6470 : _GEN_8591; // @[decode.scala 431:29]
  wire  _GEN_9232 = 3'h0 == branchTracker ? _GEN_6471 : _GEN_8592; // @[decode.scala 431:29]
  wire  _GEN_9233 = 3'h0 == branchTracker ? _GEN_6472 : _GEN_8593; // @[decode.scala 431:29]
  wire  _GEN_9234 = 3'h0 == branchTracker ? _GEN_6473 : _GEN_8594; // @[decode.scala 431:29]
  wire  _GEN_9235 = 3'h0 == branchTracker ? _GEN_6474 : _GEN_8595; // @[decode.scala 431:29]
  wire  _GEN_9236 = 3'h0 == branchTracker ? _GEN_6475 : _GEN_8596; // @[decode.scala 431:29]
  wire  _GEN_9237 = 3'h0 == branchTracker ? _GEN_6476 : _GEN_8597; // @[decode.scala 431:29]
  wire  _GEN_9238 = 3'h0 == branchTracker ? _GEN_6477 : _GEN_8598; // @[decode.scala 431:29]
  wire  _GEN_9239 = 3'h0 == branchTracker ? _GEN_6478 : _GEN_8599; // @[decode.scala 431:29]
  wire  _GEN_9240 = 3'h0 == branchTracker ? _GEN_6479 : _GEN_8600; // @[decode.scala 431:29]
  wire  _GEN_9241 = 3'h0 == branchTracker ? _GEN_6480 : _GEN_8601; // @[decode.scala 431:29]
  wire  _GEN_9242 = 3'h0 == branchTracker ? _GEN_6481 : _GEN_8602; // @[decode.scala 431:29]
  wire  _GEN_9243 = 3'h0 == branchTracker ? _GEN_6482 : _GEN_8603; // @[decode.scala 431:29]
  wire  _GEN_9244 = 3'h0 == branchTracker ? _GEN_6483 : _GEN_8604; // @[decode.scala 431:29]
  wire  _GEN_9245 = 3'h0 == branchTracker ? _GEN_6484 : _GEN_8605; // @[decode.scala 431:29]
  wire  _GEN_9246 = 3'h0 == branchTracker ? _GEN_6485 : _GEN_8606; // @[decode.scala 431:29]
  wire  _GEN_9247 = 3'h0 == branchTracker ? _GEN_6486 : _GEN_8607; // @[decode.scala 431:29]
  wire  _GEN_9248 = 3'h0 == branchTracker ? _GEN_6487 : _GEN_8608; // @[decode.scala 431:29]
  wire  _GEN_9249 = 3'h0 == branchTracker ? _GEN_6488 : _GEN_8609; // @[decode.scala 431:29]
  wire  _GEN_9250 = 3'h0 == branchTracker ? _GEN_6489 : _GEN_8610; // @[decode.scala 431:29]
  wire  _GEN_9251 = 3'h0 == branchTracker ? _GEN_6490 : _GEN_8611; // @[decode.scala 431:29]
  wire  _GEN_9252 = 3'h0 == branchTracker ? _GEN_6491 : _GEN_8612; // @[decode.scala 431:29]
  wire  _GEN_9253 = 3'h0 == branchTracker ? _GEN_6492 : _GEN_8613; // @[decode.scala 431:29]
  wire  _GEN_9254 = 3'h0 == branchTracker ? _GEN_6493 : _GEN_8614; // @[decode.scala 431:29]
  wire  _GEN_9255 = 3'h0 == branchTracker ? _GEN_6494 : _GEN_8615; // @[decode.scala 431:29]
  wire  _GEN_9256 = 3'h0 == branchTracker ? _GEN_6495 : _GEN_8616; // @[decode.scala 431:29]
  wire  _GEN_9257 = 3'h0 == branchTracker ? _GEN_6496 : _GEN_8617; // @[decode.scala 431:29]
  wire  _GEN_9258 = 3'h0 == branchTracker ? _GEN_6497 : _GEN_8618; // @[decode.scala 431:29]
  wire  _GEN_9259 = 3'h0 == branchTracker ? _GEN_6498 : _GEN_8619; // @[decode.scala 431:29]
  wire  _GEN_9260 = 3'h0 == branchTracker ? _GEN_6499 : _GEN_8620; // @[decode.scala 431:29]
  wire  _GEN_9358 = 3'h0 == branchTracker ? _GEN_6501 : _GEN_8718; // @[decode.scala 431:29]
  wire  _GEN_9359 = 3'h0 == branchTracker ? _GEN_6502 : _GEN_8719; // @[decode.scala 431:29]
  wire  _GEN_9360 = 3'h0 == branchTracker ? _GEN_6503 : _GEN_8720; // @[decode.scala 431:29]
  wire  _GEN_9361 = 3'h0 == branchTracker ? _GEN_6504 : _GEN_8721; // @[decode.scala 431:29]
  wire  _GEN_9362 = 3'h0 == branchTracker ? _GEN_6505 : _GEN_8722; // @[decode.scala 431:29]
  wire  _GEN_9363 = 3'h0 == branchTracker ? _GEN_6506 : _GEN_8723; // @[decode.scala 431:29]
  wire  _GEN_9364 = 3'h0 == branchTracker ? _GEN_6507 : _GEN_8724; // @[decode.scala 431:29]
  wire  _GEN_9365 = 3'h0 == branchTracker ? _GEN_6508 : _GEN_8725; // @[decode.scala 431:29]
  wire  _GEN_9366 = 3'h0 == branchTracker ? _GEN_6509 : _GEN_8726; // @[decode.scala 431:29]
  wire  _GEN_9367 = 3'h0 == branchTracker ? _GEN_6510 : _GEN_8727; // @[decode.scala 431:29]
  wire  _GEN_9368 = 3'h0 == branchTracker ? _GEN_6511 : _GEN_8728; // @[decode.scala 431:29]
  wire  _GEN_9369 = 3'h0 == branchTracker ? _GEN_6512 : _GEN_8729; // @[decode.scala 431:29]
  wire  _GEN_9370 = 3'h0 == branchTracker ? _GEN_6513 : _GEN_8730; // @[decode.scala 431:29]
  wire  _GEN_9371 = 3'h0 == branchTracker ? _GEN_6514 : _GEN_8731; // @[decode.scala 431:29]
  wire  _GEN_9372 = 3'h0 == branchTracker ? _GEN_6515 : _GEN_8732; // @[decode.scala 431:29]
  wire  _GEN_9373 = 3'h0 == branchTracker ? _GEN_6516 : _GEN_8733; // @[decode.scala 431:29]
  wire  _GEN_9374 = 3'h0 == branchTracker ? _GEN_6517 : _GEN_8734; // @[decode.scala 431:29]
  wire  _GEN_9375 = 3'h0 == branchTracker ? _GEN_6518 : _GEN_8735; // @[decode.scala 431:29]
  wire  _GEN_9376 = 3'h0 == branchTracker ? _GEN_6519 : _GEN_8736; // @[decode.scala 431:29]
  wire  _GEN_9377 = 3'h0 == branchTracker ? _GEN_6520 : _GEN_8737; // @[decode.scala 431:29]
  wire  _GEN_9378 = 3'h0 == branchTracker ? _GEN_6521 : _GEN_8738; // @[decode.scala 431:29]
  wire  _GEN_9379 = 3'h0 == branchTracker ? _GEN_6522 : _GEN_8739; // @[decode.scala 431:29]
  wire  _GEN_9380 = 3'h0 == branchTracker ? _GEN_6523 : _GEN_8740; // @[decode.scala 431:29]
  wire  _GEN_9381 = 3'h0 == branchTracker ? _GEN_6524 : _GEN_8741; // @[decode.scala 431:29]
  wire  _GEN_9382 = 3'h0 == branchTracker ? _GEN_6525 : _GEN_8742; // @[decode.scala 431:29]
  wire  _GEN_9383 = 3'h0 == branchTracker ? _GEN_6526 : _GEN_8743; // @[decode.scala 431:29]
  wire  _GEN_9384 = 3'h0 == branchTracker ? _GEN_6527 : _GEN_8744; // @[decode.scala 431:29]
  wire  _GEN_9385 = 3'h0 == branchTracker ? _GEN_6528 : _GEN_8745; // @[decode.scala 431:29]
  wire  _GEN_9386 = 3'h0 == branchTracker ? _GEN_6529 : _GEN_8746; // @[decode.scala 431:29]
  wire  _GEN_9387 = 3'h0 == branchTracker ? _GEN_6530 : _GEN_8747; // @[decode.scala 431:29]
  wire  _GEN_9388 = 3'h0 == branchTracker ? _GEN_6531 : _GEN_8748; // @[decode.scala 431:29]
  wire  _GEN_9389 = 3'h0 == branchTracker ? _GEN_6532 : _GEN_8749; // @[decode.scala 431:29]
  wire  _GEN_9390 = 3'h0 == branchTracker ? _GEN_6533 : _GEN_8750; // @[decode.scala 431:29]
  wire  _GEN_9391 = 3'h0 == branchTracker ? _GEN_6534 : _GEN_8751; // @[decode.scala 431:29]
  wire  _GEN_9392 = 3'h0 == branchTracker ? _GEN_6535 : _GEN_8752; // @[decode.scala 431:29]
  wire  _GEN_9393 = 3'h0 == branchTracker ? _GEN_6536 : _GEN_8753; // @[decode.scala 431:29]
  wire  _GEN_9394 = 3'h0 == branchTracker ? _GEN_6537 : _GEN_8754; // @[decode.scala 431:29]
  wire  _GEN_9395 = 3'h0 == branchTracker ? _GEN_6538 : _GEN_8755; // @[decode.scala 431:29]
  wire  _GEN_9396 = 3'h0 == branchTracker ? _GEN_6539 : _GEN_8756; // @[decode.scala 431:29]
  wire  _GEN_9397 = 3'h0 == branchTracker ? _GEN_6540 : _GEN_8757; // @[decode.scala 431:29]
  wire  _GEN_9398 = 3'h0 == branchTracker ? _GEN_6541 : _GEN_8758; // @[decode.scala 431:29]
  wire  _GEN_9399 = 3'h0 == branchTracker ? _GEN_6542 : _GEN_8759; // @[decode.scala 431:29]
  wire  _GEN_9400 = 3'h0 == branchTracker ? _GEN_6543 : _GEN_8760; // @[decode.scala 431:29]
  wire  _GEN_9401 = 3'h0 == branchTracker ? _GEN_6544 : _GEN_8761; // @[decode.scala 431:29]
  wire  _GEN_9402 = 3'h0 == branchTracker ? _GEN_6545 : _GEN_8762; // @[decode.scala 431:29]
  wire  _GEN_9403 = 3'h0 == branchTracker ? _GEN_6546 : _GEN_8763; // @[decode.scala 431:29]
  wire  _GEN_9404 = 3'h0 == branchTracker ? _GEN_6547 : _GEN_8764; // @[decode.scala 431:29]
  wire  _GEN_9405 = 3'h0 == branchTracker ? _GEN_6548 : _GEN_8765; // @[decode.scala 431:29]
  wire  _GEN_9406 = 3'h0 == branchTracker ? _GEN_6549 : _GEN_8766; // @[decode.scala 431:29]
  wire  _GEN_9407 = 3'h0 == branchTracker ? _GEN_6550 : _GEN_8767; // @[decode.scala 431:29]
  wire  _GEN_9408 = 3'h0 == branchTracker ? _GEN_6551 : _GEN_8768; // @[decode.scala 431:29]
  wire  _GEN_9409 = 3'h0 == branchTracker ? _GEN_6552 : _GEN_8769; // @[decode.scala 431:29]
  wire  _GEN_9410 = 3'h0 == branchTracker ? _GEN_6553 : _GEN_8770; // @[decode.scala 431:29]
  wire  _GEN_9411 = 3'h0 == branchTracker ? _GEN_6554 : _GEN_8771; // @[decode.scala 431:29]
  wire  _GEN_9412 = 3'h0 == branchTracker ? _GEN_6555 : _GEN_8772; // @[decode.scala 431:29]
  wire  _GEN_9413 = 3'h0 == branchTracker ? _GEN_6556 : _GEN_8773; // @[decode.scala 431:29]
  wire  _GEN_9414 = 3'h0 == branchTracker ? _GEN_6557 : _GEN_8774; // @[decode.scala 431:29]
  wire  _GEN_9415 = 3'h0 == branchTracker ? _GEN_6558 : _GEN_8775; // @[decode.scala 431:29]
  wire  _GEN_9416 = 3'h0 == branchTracker ? _GEN_6559 : _GEN_8776; // @[decode.scala 431:29]
  wire  _GEN_9417 = 3'h0 == branchTracker ? _GEN_6560 : _GEN_8777; // @[decode.scala 431:29]
  wire  _GEN_9418 = 3'h0 == branchTracker ? _GEN_6561 : _GEN_8778; // @[decode.scala 431:29]
  wire  _GEN_9419 = 3'h0 == branchTracker ? _GEN_6562 : _GEN_8779; // @[decode.scala 431:29]
  wire  _GEN_9420 = 3'h0 == branchTracker ? _GEN_6563 : _GEN_8780; // @[decode.scala 431:29]
  wire  _GEN_9518 = 3'h0 == branchTracker ? reservedFreeList4_0 : _GEN_8878; // @[decode.scala 431:29 325:30]
  wire  _GEN_9519 = 3'h0 == branchTracker ? reservedFreeList4_1 : _GEN_8879; // @[decode.scala 431:29 325:30]
  wire  _GEN_9520 = 3'h0 == branchTracker ? reservedFreeList4_2 : _GEN_8880; // @[decode.scala 431:29 325:30]
  wire  _GEN_9521 = 3'h0 == branchTracker ? reservedFreeList4_3 : _GEN_8881; // @[decode.scala 431:29 325:30]
  wire  _GEN_9522 = 3'h0 == branchTracker ? reservedFreeList4_4 : _GEN_8882; // @[decode.scala 431:29 325:30]
  wire  _GEN_9523 = 3'h0 == branchTracker ? reservedFreeList4_5 : _GEN_8883; // @[decode.scala 431:29 325:30]
  wire  _GEN_9524 = 3'h0 == branchTracker ? reservedFreeList4_6 : _GEN_8884; // @[decode.scala 431:29 325:30]
  wire  _GEN_9525 = 3'h0 == branchTracker ? reservedFreeList4_7 : _GEN_8885; // @[decode.scala 431:29 325:30]
  wire  _GEN_9526 = 3'h0 == branchTracker ? reservedFreeList4_8 : _GEN_8886; // @[decode.scala 431:29 325:30]
  wire  _GEN_9527 = 3'h0 == branchTracker ? reservedFreeList4_9 : _GEN_8887; // @[decode.scala 431:29 325:30]
  wire  _GEN_9528 = 3'h0 == branchTracker ? reservedFreeList4_10 : _GEN_8888; // @[decode.scala 431:29 325:30]
  wire  _GEN_9529 = 3'h0 == branchTracker ? reservedFreeList4_11 : _GEN_8889; // @[decode.scala 431:29 325:30]
  wire  _GEN_9530 = 3'h0 == branchTracker ? reservedFreeList4_12 : _GEN_8890; // @[decode.scala 431:29 325:30]
  wire  _GEN_9531 = 3'h0 == branchTracker ? reservedFreeList4_13 : _GEN_8891; // @[decode.scala 431:29 325:30]
  wire  _GEN_9532 = 3'h0 == branchTracker ? reservedFreeList4_14 : _GEN_8892; // @[decode.scala 431:29 325:30]
  wire  _GEN_9533 = 3'h0 == branchTracker ? reservedFreeList4_15 : _GEN_8893; // @[decode.scala 431:29 325:30]
  wire  _GEN_9534 = 3'h0 == branchTracker ? reservedFreeList4_16 : _GEN_8894; // @[decode.scala 431:29 325:30]
  wire  _GEN_9535 = 3'h0 == branchTracker ? reservedFreeList4_17 : _GEN_8895; // @[decode.scala 431:29 325:30]
  wire  _GEN_9536 = 3'h0 == branchTracker ? reservedFreeList4_18 : _GEN_8896; // @[decode.scala 431:29 325:30]
  wire  _GEN_9537 = 3'h0 == branchTracker ? reservedFreeList4_19 : _GEN_8897; // @[decode.scala 431:29 325:30]
  wire  _GEN_9538 = 3'h0 == branchTracker ? reservedFreeList4_20 : _GEN_8898; // @[decode.scala 431:29 325:30]
  wire  _GEN_9539 = 3'h0 == branchTracker ? reservedFreeList4_21 : _GEN_8899; // @[decode.scala 431:29 325:30]
  wire  _GEN_9540 = 3'h0 == branchTracker ? reservedFreeList4_22 : _GEN_8900; // @[decode.scala 431:29 325:30]
  wire  _GEN_9541 = 3'h0 == branchTracker ? reservedFreeList4_23 : _GEN_8901; // @[decode.scala 431:29 325:30]
  wire  _GEN_9542 = 3'h0 == branchTracker ? reservedFreeList4_24 : _GEN_8902; // @[decode.scala 431:29 325:30]
  wire  _GEN_9543 = 3'h0 == branchTracker ? reservedFreeList4_25 : _GEN_8903; // @[decode.scala 431:29 325:30]
  wire  _GEN_9544 = 3'h0 == branchTracker ? reservedFreeList4_26 : _GEN_8904; // @[decode.scala 431:29 325:30]
  wire  _GEN_9545 = 3'h0 == branchTracker ? reservedFreeList4_27 : _GEN_8905; // @[decode.scala 431:29 325:30]
  wire  _GEN_9546 = 3'h0 == branchTracker ? reservedFreeList4_28 : _GEN_8906; // @[decode.scala 431:29 325:30]
  wire  _GEN_9547 = 3'h0 == branchTracker ? reservedFreeList4_29 : _GEN_8907; // @[decode.scala 431:29 325:30]
  wire  _GEN_9548 = 3'h0 == branchTracker ? reservedFreeList4_30 : _GEN_8908; // @[decode.scala 431:29 325:30]
  wire  _GEN_9549 = 3'h0 == branchTracker ? reservedFreeList4_31 : _GEN_8909; // @[decode.scala 431:29 325:30]
  wire  _GEN_9550 = 3'h0 == branchTracker ? reservedFreeList4_32 : _GEN_8910; // @[decode.scala 431:29 325:30]
  wire  _GEN_9551 = 3'h0 == branchTracker ? reservedFreeList4_33 : _GEN_8911; // @[decode.scala 431:29 325:30]
  wire  _GEN_9552 = 3'h0 == branchTracker ? reservedFreeList4_34 : _GEN_8912; // @[decode.scala 431:29 325:30]
  wire  _GEN_9553 = 3'h0 == branchTracker ? reservedFreeList4_35 : _GEN_8913; // @[decode.scala 431:29 325:30]
  wire  _GEN_9554 = 3'h0 == branchTracker ? reservedFreeList4_36 : _GEN_8914; // @[decode.scala 431:29 325:30]
  wire  _GEN_9555 = 3'h0 == branchTracker ? reservedFreeList4_37 : _GEN_8915; // @[decode.scala 431:29 325:30]
  wire  _GEN_9556 = 3'h0 == branchTracker ? reservedFreeList4_38 : _GEN_8916; // @[decode.scala 431:29 325:30]
  wire  _GEN_9557 = 3'h0 == branchTracker ? reservedFreeList4_39 : _GEN_8917; // @[decode.scala 431:29 325:30]
  wire  _GEN_9558 = 3'h0 == branchTracker ? reservedFreeList4_40 : _GEN_8918; // @[decode.scala 431:29 325:30]
  wire  _GEN_9559 = 3'h0 == branchTracker ? reservedFreeList4_41 : _GEN_8919; // @[decode.scala 431:29 325:30]
  wire  _GEN_9560 = 3'h0 == branchTracker ? reservedFreeList4_42 : _GEN_8920; // @[decode.scala 431:29 325:30]
  wire  _GEN_9561 = 3'h0 == branchTracker ? reservedFreeList4_43 : _GEN_8921; // @[decode.scala 431:29 325:30]
  wire  _GEN_9562 = 3'h0 == branchTracker ? reservedFreeList4_44 : _GEN_8922; // @[decode.scala 431:29 325:30]
  wire  _GEN_9563 = 3'h0 == branchTracker ? reservedFreeList4_45 : _GEN_8923; // @[decode.scala 431:29 325:30]
  wire  _GEN_9564 = 3'h0 == branchTracker ? reservedFreeList4_46 : _GEN_8924; // @[decode.scala 431:29 325:30]
  wire  _GEN_9565 = 3'h0 == branchTracker ? reservedFreeList4_47 : _GEN_8925; // @[decode.scala 431:29 325:30]
  wire  _GEN_9566 = 3'h0 == branchTracker ? reservedFreeList4_48 : _GEN_8926; // @[decode.scala 431:29 325:30]
  wire  _GEN_9567 = 3'h0 == branchTracker ? reservedFreeList4_49 : _GEN_8927; // @[decode.scala 431:29 325:30]
  wire  _GEN_9568 = 3'h0 == branchTracker ? reservedFreeList4_50 : _GEN_8928; // @[decode.scala 431:29 325:30]
  wire  _GEN_9569 = 3'h0 == branchTracker ? reservedFreeList4_51 : _GEN_8929; // @[decode.scala 431:29 325:30]
  wire  _GEN_9570 = 3'h0 == branchTracker ? reservedFreeList4_52 : _GEN_8930; // @[decode.scala 431:29 325:30]
  wire  _GEN_9571 = 3'h0 == branchTracker ? reservedFreeList4_53 : _GEN_8931; // @[decode.scala 431:29 325:30]
  wire  _GEN_9572 = 3'h0 == branchTracker ? reservedFreeList4_54 : _GEN_8932; // @[decode.scala 431:29 325:30]
  wire  _GEN_9573 = 3'h0 == branchTracker ? reservedFreeList4_55 : _GEN_8933; // @[decode.scala 431:29 325:30]
  wire  _GEN_9574 = 3'h0 == branchTracker ? reservedFreeList4_56 : _GEN_8934; // @[decode.scala 431:29 325:30]
  wire  _GEN_9575 = 3'h0 == branchTracker ? reservedFreeList4_57 : _GEN_8935; // @[decode.scala 431:29 325:30]
  wire  _GEN_9576 = 3'h0 == branchTracker ? reservedFreeList4_58 : _GEN_8936; // @[decode.scala 431:29 325:30]
  wire  _GEN_9577 = 3'h0 == branchTracker ? reservedFreeList4_59 : _GEN_8937; // @[decode.scala 431:29 325:30]
  wire  _GEN_9578 = 3'h0 == branchTracker ? reservedFreeList4_60 : _GEN_8938; // @[decode.scala 431:29 325:30]
  wire  _GEN_9579 = 3'h0 == branchTracker ? reservedFreeList4_61 : _GEN_8939; // @[decode.scala 431:29 325:30]
  wire  _GEN_9580 = 3'h0 == branchTracker ? reservedFreeList4_62 : _GEN_8940; // @[decode.scala 431:29 325:30]
  wire [2:0] _branchTracker_T_3 = branchTracker + 3'h1; // @[decode.scala 473:38]
  wire  _GEN_9652 = _T_442 | _T_444 | _T_441 ? _GEN_6761 : _GEN_6113; // @[decode.scala 420:73]
  wire  _GEN_9686 = _T_442 | _T_444 | _T_441 ? _GEN_9038 : _GEN_6373; // @[decode.scala 420:73]
  wire  _GEN_9687 = _T_442 | _T_444 | _T_441 ? _GEN_9039 : _GEN_6374; // @[decode.scala 420:73]
  wire  _GEN_9688 = _T_442 | _T_444 | _T_441 ? _GEN_9040 : _GEN_6375; // @[decode.scala 420:73]
  wire  _GEN_9689 = _T_442 | _T_444 | _T_441 ? _GEN_9041 : _GEN_6376; // @[decode.scala 420:73]
  wire  _GEN_9690 = _T_442 | _T_444 | _T_441 ? _GEN_9042 : _GEN_6377; // @[decode.scala 420:73]
  wire  _GEN_9691 = _T_442 | _T_444 | _T_441 ? _GEN_9043 : _GEN_6378; // @[decode.scala 420:73]
  wire  _GEN_9692 = _T_442 | _T_444 | _T_441 ? _GEN_9044 : _GEN_6379; // @[decode.scala 420:73]
  wire  _GEN_9693 = _T_442 | _T_444 | _T_441 ? _GEN_9045 : _GEN_6380; // @[decode.scala 420:73]
  wire  _GEN_9694 = _T_442 | _T_444 | _T_441 ? _GEN_9046 : _GEN_6381; // @[decode.scala 420:73]
  wire  _GEN_9695 = _T_442 | _T_444 | _T_441 ? _GEN_9047 : _GEN_6382; // @[decode.scala 420:73]
  wire  _GEN_9696 = _T_442 | _T_444 | _T_441 ? _GEN_9048 : _GEN_6383; // @[decode.scala 420:73]
  wire  _GEN_9697 = _T_442 | _T_444 | _T_441 ? _GEN_9049 : _GEN_6384; // @[decode.scala 420:73]
  wire  _GEN_9698 = _T_442 | _T_444 | _T_441 ? _GEN_9050 : _GEN_6385; // @[decode.scala 420:73]
  wire  _GEN_9699 = _T_442 | _T_444 | _T_441 ? _GEN_9051 : _GEN_6386; // @[decode.scala 420:73]
  wire  _GEN_9700 = _T_442 | _T_444 | _T_441 ? _GEN_9052 : _GEN_6387; // @[decode.scala 420:73]
  wire  _GEN_9701 = _T_442 | _T_444 | _T_441 ? _GEN_9053 : _GEN_6388; // @[decode.scala 420:73]
  wire  _GEN_9702 = _T_442 | _T_444 | _T_441 ? _GEN_9054 : _GEN_6389; // @[decode.scala 420:73]
  wire  _GEN_9703 = _T_442 | _T_444 | _T_441 ? _GEN_9055 : _GEN_6390; // @[decode.scala 420:73]
  wire  _GEN_9704 = _T_442 | _T_444 | _T_441 ? _GEN_9056 : _GEN_6391; // @[decode.scala 420:73]
  wire  _GEN_9705 = _T_442 | _T_444 | _T_441 ? _GEN_9057 : _GEN_6392; // @[decode.scala 420:73]
  wire  _GEN_9706 = _T_442 | _T_444 | _T_441 ? _GEN_9058 : _GEN_6393; // @[decode.scala 420:73]
  wire  _GEN_9707 = _T_442 | _T_444 | _T_441 ? _GEN_9059 : _GEN_6394; // @[decode.scala 420:73]
  wire  _GEN_9708 = _T_442 | _T_444 | _T_441 ? _GEN_9060 : _GEN_6395; // @[decode.scala 420:73]
  wire  _GEN_9709 = _T_442 | _T_444 | _T_441 ? _GEN_9061 : _GEN_6396; // @[decode.scala 420:73]
  wire  _GEN_9710 = _T_442 | _T_444 | _T_441 ? _GEN_9062 : _GEN_6397; // @[decode.scala 420:73]
  wire  _GEN_9711 = _T_442 | _T_444 | _T_441 ? _GEN_9063 : _GEN_6398; // @[decode.scala 420:73]
  wire  _GEN_9712 = _T_442 | _T_444 | _T_441 ? _GEN_9064 : _GEN_6399; // @[decode.scala 420:73]
  wire  _GEN_9713 = _T_442 | _T_444 | _T_441 ? _GEN_9065 : _GEN_6400; // @[decode.scala 420:73]
  wire  _GEN_9714 = _T_442 | _T_444 | _T_441 ? _GEN_9066 : _GEN_6401; // @[decode.scala 420:73]
  wire  _GEN_9715 = _T_442 | _T_444 | _T_441 ? _GEN_9067 : _GEN_6402; // @[decode.scala 420:73]
  wire  _GEN_9716 = _T_442 | _T_444 | _T_441 ? _GEN_9068 : _GEN_6403; // @[decode.scala 420:73]
  wire  _GEN_9717 = _T_442 | _T_444 | _T_441 ? _GEN_9069 : _GEN_6404; // @[decode.scala 420:73]
  wire  _GEN_9718 = _T_442 | _T_444 | _T_441 ? _GEN_9070 : _GEN_6405; // @[decode.scala 420:73]
  wire  _GEN_9719 = _T_442 | _T_444 | _T_441 ? _GEN_9071 : _GEN_6406; // @[decode.scala 420:73]
  wire  _GEN_9720 = _T_442 | _T_444 | _T_441 ? _GEN_9072 : _GEN_6407; // @[decode.scala 420:73]
  wire  _GEN_9721 = _T_442 | _T_444 | _T_441 ? _GEN_9073 : _GEN_6408; // @[decode.scala 420:73]
  wire  _GEN_9722 = _T_442 | _T_444 | _T_441 ? _GEN_9074 : _GEN_6409; // @[decode.scala 420:73]
  wire  _GEN_9723 = _T_442 | _T_444 | _T_441 ? _GEN_9075 : _GEN_6410; // @[decode.scala 420:73]
  wire  _GEN_9724 = _T_442 | _T_444 | _T_441 ? _GEN_9076 : _GEN_6411; // @[decode.scala 420:73]
  wire  _GEN_9725 = _T_442 | _T_444 | _T_441 ? _GEN_9077 : _GEN_6412; // @[decode.scala 420:73]
  wire  _GEN_9726 = _T_442 | _T_444 | _T_441 ? _GEN_9078 : _GEN_6413; // @[decode.scala 420:73]
  wire  _GEN_9727 = _T_442 | _T_444 | _T_441 ? _GEN_9079 : _GEN_6414; // @[decode.scala 420:73]
  wire  _GEN_9728 = _T_442 | _T_444 | _T_441 ? _GEN_9080 : _GEN_6415; // @[decode.scala 420:73]
  wire  _GEN_9729 = _T_442 | _T_444 | _T_441 ? _GEN_9081 : _GEN_6416; // @[decode.scala 420:73]
  wire  _GEN_9730 = _T_442 | _T_444 | _T_441 ? _GEN_9082 : _GEN_6417; // @[decode.scala 420:73]
  wire  _GEN_9731 = _T_442 | _T_444 | _T_441 ? _GEN_9083 : _GEN_6418; // @[decode.scala 420:73]
  wire  _GEN_9732 = _T_442 | _T_444 | _T_441 ? _GEN_9084 : _GEN_6419; // @[decode.scala 420:73]
  wire  _GEN_9733 = _T_442 | _T_444 | _T_441 ? _GEN_9085 : _GEN_6420; // @[decode.scala 420:73]
  wire  _GEN_9734 = _T_442 | _T_444 | _T_441 ? _GEN_9086 : _GEN_6421; // @[decode.scala 420:73]
  wire  _GEN_9735 = _T_442 | _T_444 | _T_441 ? _GEN_9087 : _GEN_6422; // @[decode.scala 420:73]
  wire  _GEN_9736 = _T_442 | _T_444 | _T_441 ? _GEN_9088 : _GEN_6423; // @[decode.scala 420:73]
  wire  _GEN_9737 = _T_442 | _T_444 | _T_441 ? _GEN_9089 : _GEN_6424; // @[decode.scala 420:73]
  wire  _GEN_9738 = _T_442 | _T_444 | _T_441 ? _GEN_9090 : _GEN_6425; // @[decode.scala 420:73]
  wire  _GEN_9739 = _T_442 | _T_444 | _T_441 ? _GEN_9091 : _GEN_6426; // @[decode.scala 420:73]
  wire  _GEN_9740 = _T_442 | _T_444 | _T_441 ? _GEN_9092 : _GEN_6427; // @[decode.scala 420:73]
  wire  _GEN_9741 = _T_442 | _T_444 | _T_441 ? _GEN_9093 : _GEN_6428; // @[decode.scala 420:73]
  wire  _GEN_9742 = _T_442 | _T_444 | _T_441 ? _GEN_9094 : _GEN_6429; // @[decode.scala 420:73]
  wire  _GEN_9743 = _T_442 | _T_444 | _T_441 ? _GEN_9095 : _GEN_6430; // @[decode.scala 420:73]
  wire  _GEN_9744 = _T_442 | _T_444 | _T_441 ? _GEN_9096 : _GEN_6431; // @[decode.scala 420:73]
  wire  _GEN_9745 = _T_442 | _T_444 | _T_441 ? _GEN_9097 : _GEN_6432; // @[decode.scala 420:73]
  wire  _GEN_9746 = _T_442 | _T_444 | _T_441 ? _GEN_9098 : _GEN_6433; // @[decode.scala 420:73]
  wire  _GEN_9747 = _T_442 | _T_444 | _T_441 ? _GEN_9099 : _GEN_6434; // @[decode.scala 420:73]
  wire  _GEN_9748 = _T_442 | _T_444 | _T_441 ? _GEN_9100 : _GEN_6435; // @[decode.scala 420:73]
  wire  _GEN_9846 = _T_442 | _T_444 | _T_441 ? _GEN_9198 : _GEN_6437; // @[decode.scala 420:73]
  wire  _GEN_9847 = _T_442 | _T_444 | _T_441 ? _GEN_9199 : _GEN_6438; // @[decode.scala 420:73]
  wire  _GEN_9848 = _T_442 | _T_444 | _T_441 ? _GEN_9200 : _GEN_6439; // @[decode.scala 420:73]
  wire  _GEN_9849 = _T_442 | _T_444 | _T_441 ? _GEN_9201 : _GEN_6440; // @[decode.scala 420:73]
  wire  _GEN_9850 = _T_442 | _T_444 | _T_441 ? _GEN_9202 : _GEN_6441; // @[decode.scala 420:73]
  wire  _GEN_9851 = _T_442 | _T_444 | _T_441 ? _GEN_9203 : _GEN_6442; // @[decode.scala 420:73]
  wire  _GEN_9852 = _T_442 | _T_444 | _T_441 ? _GEN_9204 : _GEN_6443; // @[decode.scala 420:73]
  wire  _GEN_9853 = _T_442 | _T_444 | _T_441 ? _GEN_9205 : _GEN_6444; // @[decode.scala 420:73]
  wire  _GEN_9854 = _T_442 | _T_444 | _T_441 ? _GEN_9206 : _GEN_6445; // @[decode.scala 420:73]
  wire  _GEN_9855 = _T_442 | _T_444 | _T_441 ? _GEN_9207 : _GEN_6446; // @[decode.scala 420:73]
  wire  _GEN_9856 = _T_442 | _T_444 | _T_441 ? _GEN_9208 : _GEN_6447; // @[decode.scala 420:73]
  wire  _GEN_9857 = _T_442 | _T_444 | _T_441 ? _GEN_9209 : _GEN_6448; // @[decode.scala 420:73]
  wire  _GEN_9858 = _T_442 | _T_444 | _T_441 ? _GEN_9210 : _GEN_6449; // @[decode.scala 420:73]
  wire  _GEN_9859 = _T_442 | _T_444 | _T_441 ? _GEN_9211 : _GEN_6450; // @[decode.scala 420:73]
  wire  _GEN_9860 = _T_442 | _T_444 | _T_441 ? _GEN_9212 : _GEN_6451; // @[decode.scala 420:73]
  wire  _GEN_9861 = _T_442 | _T_444 | _T_441 ? _GEN_9213 : _GEN_6452; // @[decode.scala 420:73]
  wire  _GEN_9862 = _T_442 | _T_444 | _T_441 ? _GEN_9214 : _GEN_6453; // @[decode.scala 420:73]
  wire  _GEN_9863 = _T_442 | _T_444 | _T_441 ? _GEN_9215 : _GEN_6454; // @[decode.scala 420:73]
  wire  _GEN_9864 = _T_442 | _T_444 | _T_441 ? _GEN_9216 : _GEN_6455; // @[decode.scala 420:73]
  wire  _GEN_9865 = _T_442 | _T_444 | _T_441 ? _GEN_9217 : _GEN_6456; // @[decode.scala 420:73]
  wire  _GEN_9866 = _T_442 | _T_444 | _T_441 ? _GEN_9218 : _GEN_6457; // @[decode.scala 420:73]
  wire  _GEN_9867 = _T_442 | _T_444 | _T_441 ? _GEN_9219 : _GEN_6458; // @[decode.scala 420:73]
  wire  _GEN_9868 = _T_442 | _T_444 | _T_441 ? _GEN_9220 : _GEN_6459; // @[decode.scala 420:73]
  wire  _GEN_9869 = _T_442 | _T_444 | _T_441 ? _GEN_9221 : _GEN_6460; // @[decode.scala 420:73]
  wire  _GEN_9870 = _T_442 | _T_444 | _T_441 ? _GEN_9222 : _GEN_6461; // @[decode.scala 420:73]
  wire  _GEN_9871 = _T_442 | _T_444 | _T_441 ? _GEN_9223 : _GEN_6462; // @[decode.scala 420:73]
  wire  _GEN_9872 = _T_442 | _T_444 | _T_441 ? _GEN_9224 : _GEN_6463; // @[decode.scala 420:73]
  wire  _GEN_9873 = _T_442 | _T_444 | _T_441 ? _GEN_9225 : _GEN_6464; // @[decode.scala 420:73]
  wire  _GEN_9874 = _T_442 | _T_444 | _T_441 ? _GEN_9226 : _GEN_6465; // @[decode.scala 420:73]
  wire  _GEN_9875 = _T_442 | _T_444 | _T_441 ? _GEN_9227 : _GEN_6466; // @[decode.scala 420:73]
  wire  _GEN_9876 = _T_442 | _T_444 | _T_441 ? _GEN_9228 : _GEN_6467; // @[decode.scala 420:73]
  wire  _GEN_9877 = _T_442 | _T_444 | _T_441 ? _GEN_9229 : _GEN_6468; // @[decode.scala 420:73]
  wire  _GEN_9878 = _T_442 | _T_444 | _T_441 ? _GEN_9230 : _GEN_6469; // @[decode.scala 420:73]
  wire  _GEN_9879 = _T_442 | _T_444 | _T_441 ? _GEN_9231 : _GEN_6470; // @[decode.scala 420:73]
  wire  _GEN_9880 = _T_442 | _T_444 | _T_441 ? _GEN_9232 : _GEN_6471; // @[decode.scala 420:73]
  wire  _GEN_9881 = _T_442 | _T_444 | _T_441 ? _GEN_9233 : _GEN_6472; // @[decode.scala 420:73]
  wire  _GEN_9882 = _T_442 | _T_444 | _T_441 ? _GEN_9234 : _GEN_6473; // @[decode.scala 420:73]
  wire  _GEN_9883 = _T_442 | _T_444 | _T_441 ? _GEN_9235 : _GEN_6474; // @[decode.scala 420:73]
  wire  _GEN_9884 = _T_442 | _T_444 | _T_441 ? _GEN_9236 : _GEN_6475; // @[decode.scala 420:73]
  wire  _GEN_9885 = _T_442 | _T_444 | _T_441 ? _GEN_9237 : _GEN_6476; // @[decode.scala 420:73]
  wire  _GEN_9886 = _T_442 | _T_444 | _T_441 ? _GEN_9238 : _GEN_6477; // @[decode.scala 420:73]
  wire  _GEN_9887 = _T_442 | _T_444 | _T_441 ? _GEN_9239 : _GEN_6478; // @[decode.scala 420:73]
  wire  _GEN_9888 = _T_442 | _T_444 | _T_441 ? _GEN_9240 : _GEN_6479; // @[decode.scala 420:73]
  wire  _GEN_9889 = _T_442 | _T_444 | _T_441 ? _GEN_9241 : _GEN_6480; // @[decode.scala 420:73]
  wire  _GEN_9890 = _T_442 | _T_444 | _T_441 ? _GEN_9242 : _GEN_6481; // @[decode.scala 420:73]
  wire  _GEN_9891 = _T_442 | _T_444 | _T_441 ? _GEN_9243 : _GEN_6482; // @[decode.scala 420:73]
  wire  _GEN_9892 = _T_442 | _T_444 | _T_441 ? _GEN_9244 : _GEN_6483; // @[decode.scala 420:73]
  wire  _GEN_9893 = _T_442 | _T_444 | _T_441 ? _GEN_9245 : _GEN_6484; // @[decode.scala 420:73]
  wire  _GEN_9894 = _T_442 | _T_444 | _T_441 ? _GEN_9246 : _GEN_6485; // @[decode.scala 420:73]
  wire  _GEN_9895 = _T_442 | _T_444 | _T_441 ? _GEN_9247 : _GEN_6486; // @[decode.scala 420:73]
  wire  _GEN_9896 = _T_442 | _T_444 | _T_441 ? _GEN_9248 : _GEN_6487; // @[decode.scala 420:73]
  wire  _GEN_9897 = _T_442 | _T_444 | _T_441 ? _GEN_9249 : _GEN_6488; // @[decode.scala 420:73]
  wire  _GEN_9898 = _T_442 | _T_444 | _T_441 ? _GEN_9250 : _GEN_6489; // @[decode.scala 420:73]
  wire  _GEN_9899 = _T_442 | _T_444 | _T_441 ? _GEN_9251 : _GEN_6490; // @[decode.scala 420:73]
  wire  _GEN_9900 = _T_442 | _T_444 | _T_441 ? _GEN_9252 : _GEN_6491; // @[decode.scala 420:73]
  wire  _GEN_9901 = _T_442 | _T_444 | _T_441 ? _GEN_9253 : _GEN_6492; // @[decode.scala 420:73]
  wire  _GEN_9902 = _T_442 | _T_444 | _T_441 ? _GEN_9254 : _GEN_6493; // @[decode.scala 420:73]
  wire  _GEN_9903 = _T_442 | _T_444 | _T_441 ? _GEN_9255 : _GEN_6494; // @[decode.scala 420:73]
  wire  _GEN_9904 = _T_442 | _T_444 | _T_441 ? _GEN_9256 : _GEN_6495; // @[decode.scala 420:73]
  wire  _GEN_9905 = _T_442 | _T_444 | _T_441 ? _GEN_9257 : _GEN_6496; // @[decode.scala 420:73]
  wire  _GEN_9906 = _T_442 | _T_444 | _T_441 ? _GEN_9258 : _GEN_6497; // @[decode.scala 420:73]
  wire  _GEN_9907 = _T_442 | _T_444 | _T_441 ? _GEN_9259 : _GEN_6498; // @[decode.scala 420:73]
  wire  _GEN_9908 = _T_442 | _T_444 | _T_441 ? _GEN_9260 : _GEN_6499; // @[decode.scala 420:73]
  wire  _GEN_10006 = _T_442 | _T_444 | _T_441 ? _GEN_9358 : _GEN_6501; // @[decode.scala 420:73]
  wire  _GEN_10007 = _T_442 | _T_444 | _T_441 ? _GEN_9359 : _GEN_6502; // @[decode.scala 420:73]
  wire  _GEN_10008 = _T_442 | _T_444 | _T_441 ? _GEN_9360 : _GEN_6503; // @[decode.scala 420:73]
  wire  _GEN_10009 = _T_442 | _T_444 | _T_441 ? _GEN_9361 : _GEN_6504; // @[decode.scala 420:73]
  wire  _GEN_10010 = _T_442 | _T_444 | _T_441 ? _GEN_9362 : _GEN_6505; // @[decode.scala 420:73]
  wire  _GEN_10011 = _T_442 | _T_444 | _T_441 ? _GEN_9363 : _GEN_6506; // @[decode.scala 420:73]
  wire  _GEN_10012 = _T_442 | _T_444 | _T_441 ? _GEN_9364 : _GEN_6507; // @[decode.scala 420:73]
  wire  _GEN_10013 = _T_442 | _T_444 | _T_441 ? _GEN_9365 : _GEN_6508; // @[decode.scala 420:73]
  wire  _GEN_10014 = _T_442 | _T_444 | _T_441 ? _GEN_9366 : _GEN_6509; // @[decode.scala 420:73]
  wire  _GEN_10015 = _T_442 | _T_444 | _T_441 ? _GEN_9367 : _GEN_6510; // @[decode.scala 420:73]
  wire  _GEN_10016 = _T_442 | _T_444 | _T_441 ? _GEN_9368 : _GEN_6511; // @[decode.scala 420:73]
  wire  _GEN_10017 = _T_442 | _T_444 | _T_441 ? _GEN_9369 : _GEN_6512; // @[decode.scala 420:73]
  wire  _GEN_10018 = _T_442 | _T_444 | _T_441 ? _GEN_9370 : _GEN_6513; // @[decode.scala 420:73]
  wire  _GEN_10019 = _T_442 | _T_444 | _T_441 ? _GEN_9371 : _GEN_6514; // @[decode.scala 420:73]
  wire  _GEN_10020 = _T_442 | _T_444 | _T_441 ? _GEN_9372 : _GEN_6515; // @[decode.scala 420:73]
  wire  _GEN_10021 = _T_442 | _T_444 | _T_441 ? _GEN_9373 : _GEN_6516; // @[decode.scala 420:73]
  wire  _GEN_10022 = _T_442 | _T_444 | _T_441 ? _GEN_9374 : _GEN_6517; // @[decode.scala 420:73]
  wire  _GEN_10023 = _T_442 | _T_444 | _T_441 ? _GEN_9375 : _GEN_6518; // @[decode.scala 420:73]
  wire  _GEN_10024 = _T_442 | _T_444 | _T_441 ? _GEN_9376 : _GEN_6519; // @[decode.scala 420:73]
  wire  _GEN_10025 = _T_442 | _T_444 | _T_441 ? _GEN_9377 : _GEN_6520; // @[decode.scala 420:73]
  wire  _GEN_10026 = _T_442 | _T_444 | _T_441 ? _GEN_9378 : _GEN_6521; // @[decode.scala 420:73]
  wire  _GEN_10027 = _T_442 | _T_444 | _T_441 ? _GEN_9379 : _GEN_6522; // @[decode.scala 420:73]
  wire  _GEN_10028 = _T_442 | _T_444 | _T_441 ? _GEN_9380 : _GEN_6523; // @[decode.scala 420:73]
  wire  _GEN_10029 = _T_442 | _T_444 | _T_441 ? _GEN_9381 : _GEN_6524; // @[decode.scala 420:73]
  wire  _GEN_10030 = _T_442 | _T_444 | _T_441 ? _GEN_9382 : _GEN_6525; // @[decode.scala 420:73]
  wire  _GEN_10031 = _T_442 | _T_444 | _T_441 ? _GEN_9383 : _GEN_6526; // @[decode.scala 420:73]
  wire  _GEN_10032 = _T_442 | _T_444 | _T_441 ? _GEN_9384 : _GEN_6527; // @[decode.scala 420:73]
  wire  _GEN_10033 = _T_442 | _T_444 | _T_441 ? _GEN_9385 : _GEN_6528; // @[decode.scala 420:73]
  wire  _GEN_10034 = _T_442 | _T_444 | _T_441 ? _GEN_9386 : _GEN_6529; // @[decode.scala 420:73]
  wire  _GEN_10035 = _T_442 | _T_444 | _T_441 ? _GEN_9387 : _GEN_6530; // @[decode.scala 420:73]
  wire  _GEN_10036 = _T_442 | _T_444 | _T_441 ? _GEN_9388 : _GEN_6531; // @[decode.scala 420:73]
  wire  _GEN_10037 = _T_442 | _T_444 | _T_441 ? _GEN_9389 : _GEN_6532; // @[decode.scala 420:73]
  wire  _GEN_10038 = _T_442 | _T_444 | _T_441 ? _GEN_9390 : _GEN_6533; // @[decode.scala 420:73]
  wire  _GEN_10039 = _T_442 | _T_444 | _T_441 ? _GEN_9391 : _GEN_6534; // @[decode.scala 420:73]
  wire  _GEN_10040 = _T_442 | _T_444 | _T_441 ? _GEN_9392 : _GEN_6535; // @[decode.scala 420:73]
  wire  _GEN_10041 = _T_442 | _T_444 | _T_441 ? _GEN_9393 : _GEN_6536; // @[decode.scala 420:73]
  wire  _GEN_10042 = _T_442 | _T_444 | _T_441 ? _GEN_9394 : _GEN_6537; // @[decode.scala 420:73]
  wire  _GEN_10043 = _T_442 | _T_444 | _T_441 ? _GEN_9395 : _GEN_6538; // @[decode.scala 420:73]
  wire  _GEN_10044 = _T_442 | _T_444 | _T_441 ? _GEN_9396 : _GEN_6539; // @[decode.scala 420:73]
  wire  _GEN_10045 = _T_442 | _T_444 | _T_441 ? _GEN_9397 : _GEN_6540; // @[decode.scala 420:73]
  wire  _GEN_10046 = _T_442 | _T_444 | _T_441 ? _GEN_9398 : _GEN_6541; // @[decode.scala 420:73]
  wire  _GEN_10047 = _T_442 | _T_444 | _T_441 ? _GEN_9399 : _GEN_6542; // @[decode.scala 420:73]
  wire  _GEN_10048 = _T_442 | _T_444 | _T_441 ? _GEN_9400 : _GEN_6543; // @[decode.scala 420:73]
  wire  _GEN_10049 = _T_442 | _T_444 | _T_441 ? _GEN_9401 : _GEN_6544; // @[decode.scala 420:73]
  wire  _GEN_10050 = _T_442 | _T_444 | _T_441 ? _GEN_9402 : _GEN_6545; // @[decode.scala 420:73]
  wire  _GEN_10051 = _T_442 | _T_444 | _T_441 ? _GEN_9403 : _GEN_6546; // @[decode.scala 420:73]
  wire  _GEN_10052 = _T_442 | _T_444 | _T_441 ? _GEN_9404 : _GEN_6547; // @[decode.scala 420:73]
  wire  _GEN_10053 = _T_442 | _T_444 | _T_441 ? _GEN_9405 : _GEN_6548; // @[decode.scala 420:73]
  wire  _GEN_10054 = _T_442 | _T_444 | _T_441 ? _GEN_9406 : _GEN_6549; // @[decode.scala 420:73]
  wire  _GEN_10055 = _T_442 | _T_444 | _T_441 ? _GEN_9407 : _GEN_6550; // @[decode.scala 420:73]
  wire  _GEN_10056 = _T_442 | _T_444 | _T_441 ? _GEN_9408 : _GEN_6551; // @[decode.scala 420:73]
  wire  _GEN_10057 = _T_442 | _T_444 | _T_441 ? _GEN_9409 : _GEN_6552; // @[decode.scala 420:73]
  wire  _GEN_10058 = _T_442 | _T_444 | _T_441 ? _GEN_9410 : _GEN_6553; // @[decode.scala 420:73]
  wire  _GEN_10059 = _T_442 | _T_444 | _T_441 ? _GEN_9411 : _GEN_6554; // @[decode.scala 420:73]
  wire  _GEN_10060 = _T_442 | _T_444 | _T_441 ? _GEN_9412 : _GEN_6555; // @[decode.scala 420:73]
  wire  _GEN_10061 = _T_442 | _T_444 | _T_441 ? _GEN_9413 : _GEN_6556; // @[decode.scala 420:73]
  wire  _GEN_10062 = _T_442 | _T_444 | _T_441 ? _GEN_9414 : _GEN_6557; // @[decode.scala 420:73]
  wire  _GEN_10063 = _T_442 | _T_444 | _T_441 ? _GEN_9415 : _GEN_6558; // @[decode.scala 420:73]
  wire  _GEN_10064 = _T_442 | _T_444 | _T_441 ? _GEN_9416 : _GEN_6559; // @[decode.scala 420:73]
  wire  _GEN_10065 = _T_442 | _T_444 | _T_441 ? _GEN_9417 : _GEN_6560; // @[decode.scala 420:73]
  wire  _GEN_10066 = _T_442 | _T_444 | _T_441 ? _GEN_9418 : _GEN_6561; // @[decode.scala 420:73]
  wire  _GEN_10067 = _T_442 | _T_444 | _T_441 ? _GEN_9419 : _GEN_6562; // @[decode.scala 420:73]
  wire  _GEN_10068 = _T_442 | _T_444 | _T_441 ? _GEN_9420 : _GEN_6563; // @[decode.scala 420:73]
  wire  _GEN_10166 = _T_442 | _T_444 | _T_441 ? _GEN_9518 : reservedFreeList4_0; // @[decode.scala 325:30 420:73]
  wire  _GEN_10167 = _T_442 | _T_444 | _T_441 ? _GEN_9519 : reservedFreeList4_1; // @[decode.scala 325:30 420:73]
  wire  _GEN_10168 = _T_442 | _T_444 | _T_441 ? _GEN_9520 : reservedFreeList4_2; // @[decode.scala 325:30 420:73]
  wire  _GEN_10169 = _T_442 | _T_444 | _T_441 ? _GEN_9521 : reservedFreeList4_3; // @[decode.scala 325:30 420:73]
  wire  _GEN_10170 = _T_442 | _T_444 | _T_441 ? _GEN_9522 : reservedFreeList4_4; // @[decode.scala 325:30 420:73]
  wire  _GEN_10171 = _T_442 | _T_444 | _T_441 ? _GEN_9523 : reservedFreeList4_5; // @[decode.scala 325:30 420:73]
  wire  _GEN_10172 = _T_442 | _T_444 | _T_441 ? _GEN_9524 : reservedFreeList4_6; // @[decode.scala 325:30 420:73]
  wire  _GEN_10173 = _T_442 | _T_444 | _T_441 ? _GEN_9525 : reservedFreeList4_7; // @[decode.scala 325:30 420:73]
  wire  _GEN_10174 = _T_442 | _T_444 | _T_441 ? _GEN_9526 : reservedFreeList4_8; // @[decode.scala 325:30 420:73]
  wire  _GEN_10175 = _T_442 | _T_444 | _T_441 ? _GEN_9527 : reservedFreeList4_9; // @[decode.scala 325:30 420:73]
  wire  _GEN_10176 = _T_442 | _T_444 | _T_441 ? _GEN_9528 : reservedFreeList4_10; // @[decode.scala 325:30 420:73]
  wire  _GEN_10177 = _T_442 | _T_444 | _T_441 ? _GEN_9529 : reservedFreeList4_11; // @[decode.scala 325:30 420:73]
  wire  _GEN_10178 = _T_442 | _T_444 | _T_441 ? _GEN_9530 : reservedFreeList4_12; // @[decode.scala 325:30 420:73]
  wire  _GEN_10179 = _T_442 | _T_444 | _T_441 ? _GEN_9531 : reservedFreeList4_13; // @[decode.scala 325:30 420:73]
  wire  _GEN_10180 = _T_442 | _T_444 | _T_441 ? _GEN_9532 : reservedFreeList4_14; // @[decode.scala 325:30 420:73]
  wire  _GEN_10181 = _T_442 | _T_444 | _T_441 ? _GEN_9533 : reservedFreeList4_15; // @[decode.scala 325:30 420:73]
  wire  _GEN_10182 = _T_442 | _T_444 | _T_441 ? _GEN_9534 : reservedFreeList4_16; // @[decode.scala 325:30 420:73]
  wire  _GEN_10183 = _T_442 | _T_444 | _T_441 ? _GEN_9535 : reservedFreeList4_17; // @[decode.scala 325:30 420:73]
  wire  _GEN_10184 = _T_442 | _T_444 | _T_441 ? _GEN_9536 : reservedFreeList4_18; // @[decode.scala 325:30 420:73]
  wire  _GEN_10185 = _T_442 | _T_444 | _T_441 ? _GEN_9537 : reservedFreeList4_19; // @[decode.scala 325:30 420:73]
  wire  _GEN_10186 = _T_442 | _T_444 | _T_441 ? _GEN_9538 : reservedFreeList4_20; // @[decode.scala 325:30 420:73]
  wire  _GEN_10187 = _T_442 | _T_444 | _T_441 ? _GEN_9539 : reservedFreeList4_21; // @[decode.scala 325:30 420:73]
  wire  _GEN_10188 = _T_442 | _T_444 | _T_441 ? _GEN_9540 : reservedFreeList4_22; // @[decode.scala 325:30 420:73]
  wire  _GEN_10189 = _T_442 | _T_444 | _T_441 ? _GEN_9541 : reservedFreeList4_23; // @[decode.scala 325:30 420:73]
  wire  _GEN_10190 = _T_442 | _T_444 | _T_441 ? _GEN_9542 : reservedFreeList4_24; // @[decode.scala 325:30 420:73]
  wire  _GEN_10191 = _T_442 | _T_444 | _T_441 ? _GEN_9543 : reservedFreeList4_25; // @[decode.scala 325:30 420:73]
  wire  _GEN_10192 = _T_442 | _T_444 | _T_441 ? _GEN_9544 : reservedFreeList4_26; // @[decode.scala 325:30 420:73]
  wire  _GEN_10193 = _T_442 | _T_444 | _T_441 ? _GEN_9545 : reservedFreeList4_27; // @[decode.scala 325:30 420:73]
  wire  _GEN_10194 = _T_442 | _T_444 | _T_441 ? _GEN_9546 : reservedFreeList4_28; // @[decode.scala 325:30 420:73]
  wire  _GEN_10195 = _T_442 | _T_444 | _T_441 ? _GEN_9547 : reservedFreeList4_29; // @[decode.scala 325:30 420:73]
  wire  _GEN_10196 = _T_442 | _T_444 | _T_441 ? _GEN_9548 : reservedFreeList4_30; // @[decode.scala 325:30 420:73]
  wire  _GEN_10197 = _T_442 | _T_444 | _T_441 ? _GEN_9549 : reservedFreeList4_31; // @[decode.scala 325:30 420:73]
  wire  _GEN_10198 = _T_442 | _T_444 | _T_441 ? _GEN_9550 : reservedFreeList4_32; // @[decode.scala 325:30 420:73]
  wire  _GEN_10199 = _T_442 | _T_444 | _T_441 ? _GEN_9551 : reservedFreeList4_33; // @[decode.scala 325:30 420:73]
  wire  _GEN_10200 = _T_442 | _T_444 | _T_441 ? _GEN_9552 : reservedFreeList4_34; // @[decode.scala 325:30 420:73]
  wire  _GEN_10201 = _T_442 | _T_444 | _T_441 ? _GEN_9553 : reservedFreeList4_35; // @[decode.scala 325:30 420:73]
  wire  _GEN_10202 = _T_442 | _T_444 | _T_441 ? _GEN_9554 : reservedFreeList4_36; // @[decode.scala 325:30 420:73]
  wire  _GEN_10203 = _T_442 | _T_444 | _T_441 ? _GEN_9555 : reservedFreeList4_37; // @[decode.scala 325:30 420:73]
  wire  _GEN_10204 = _T_442 | _T_444 | _T_441 ? _GEN_9556 : reservedFreeList4_38; // @[decode.scala 325:30 420:73]
  wire  _GEN_10205 = _T_442 | _T_444 | _T_441 ? _GEN_9557 : reservedFreeList4_39; // @[decode.scala 325:30 420:73]
  wire  _GEN_10206 = _T_442 | _T_444 | _T_441 ? _GEN_9558 : reservedFreeList4_40; // @[decode.scala 325:30 420:73]
  wire  _GEN_10207 = _T_442 | _T_444 | _T_441 ? _GEN_9559 : reservedFreeList4_41; // @[decode.scala 325:30 420:73]
  wire  _GEN_10208 = _T_442 | _T_444 | _T_441 ? _GEN_9560 : reservedFreeList4_42; // @[decode.scala 325:30 420:73]
  wire  _GEN_10209 = _T_442 | _T_444 | _T_441 ? _GEN_9561 : reservedFreeList4_43; // @[decode.scala 325:30 420:73]
  wire  _GEN_10210 = _T_442 | _T_444 | _T_441 ? _GEN_9562 : reservedFreeList4_44; // @[decode.scala 325:30 420:73]
  wire  _GEN_10211 = _T_442 | _T_444 | _T_441 ? _GEN_9563 : reservedFreeList4_45; // @[decode.scala 325:30 420:73]
  wire  _GEN_10212 = _T_442 | _T_444 | _T_441 ? _GEN_9564 : reservedFreeList4_46; // @[decode.scala 325:30 420:73]
  wire  _GEN_10213 = _T_442 | _T_444 | _T_441 ? _GEN_9565 : reservedFreeList4_47; // @[decode.scala 325:30 420:73]
  wire  _GEN_10214 = _T_442 | _T_444 | _T_441 ? _GEN_9566 : reservedFreeList4_48; // @[decode.scala 325:30 420:73]
  wire  _GEN_10215 = _T_442 | _T_444 | _T_441 ? _GEN_9567 : reservedFreeList4_49; // @[decode.scala 325:30 420:73]
  wire  _GEN_10216 = _T_442 | _T_444 | _T_441 ? _GEN_9568 : reservedFreeList4_50; // @[decode.scala 325:30 420:73]
  wire  _GEN_10217 = _T_442 | _T_444 | _T_441 ? _GEN_9569 : reservedFreeList4_51; // @[decode.scala 325:30 420:73]
  wire  _GEN_10218 = _T_442 | _T_444 | _T_441 ? _GEN_9570 : reservedFreeList4_52; // @[decode.scala 325:30 420:73]
  wire  _GEN_10219 = _T_442 | _T_444 | _T_441 ? _GEN_9571 : reservedFreeList4_53; // @[decode.scala 325:30 420:73]
  wire  _GEN_10220 = _T_442 | _T_444 | _T_441 ? _GEN_9572 : reservedFreeList4_54; // @[decode.scala 325:30 420:73]
  wire  _GEN_10221 = _T_442 | _T_444 | _T_441 ? _GEN_9573 : reservedFreeList4_55; // @[decode.scala 325:30 420:73]
  wire  _GEN_10222 = _T_442 | _T_444 | _T_441 ? _GEN_9574 : reservedFreeList4_56; // @[decode.scala 325:30 420:73]
  wire  _GEN_10223 = _T_442 | _T_444 | _T_441 ? _GEN_9575 : reservedFreeList4_57; // @[decode.scala 325:30 420:73]
  wire  _GEN_10224 = _T_442 | _T_444 | _T_441 ? _GEN_9576 : reservedFreeList4_58; // @[decode.scala 325:30 420:73]
  wire  _GEN_10225 = _T_442 | _T_444 | _T_441 ? _GEN_9577 : reservedFreeList4_59; // @[decode.scala 325:30 420:73]
  wire  _GEN_10226 = _T_442 | _T_444 | _T_441 ? _GEN_9578 : reservedFreeList4_60; // @[decode.scala 325:30 420:73]
  wire  _GEN_10227 = _T_442 | _T_444 | _T_441 ? _GEN_9579 : reservedFreeList4_61; // @[decode.scala 325:30 420:73]
  wire  _GEN_10228 = _T_442 | _T_444 | _T_441 ? _GEN_9580 : reservedFreeList4_62; // @[decode.scala 325:30 420:73]
  wire  _GEN_10301 = _T_3 ? _GEN_9652 : _GEN_6113; // @[decode.scala 419:41]
  wire  _GEN_10335 = _T_3 ? _GEN_9686 : _GEN_6373; // @[decode.scala 419:41]
  wire  _GEN_10336 = _T_3 ? _GEN_9687 : _GEN_6374; // @[decode.scala 419:41]
  wire  _GEN_10337 = _T_3 ? _GEN_9688 : _GEN_6375; // @[decode.scala 419:41]
  wire  _GEN_10338 = _T_3 ? _GEN_9689 : _GEN_6376; // @[decode.scala 419:41]
  wire  _GEN_10339 = _T_3 ? _GEN_9690 : _GEN_6377; // @[decode.scala 419:41]
  wire  _GEN_10340 = _T_3 ? _GEN_9691 : _GEN_6378; // @[decode.scala 419:41]
  wire  _GEN_10341 = _T_3 ? _GEN_9692 : _GEN_6379; // @[decode.scala 419:41]
  wire  _GEN_10342 = _T_3 ? _GEN_9693 : _GEN_6380; // @[decode.scala 419:41]
  wire  _GEN_10343 = _T_3 ? _GEN_9694 : _GEN_6381; // @[decode.scala 419:41]
  wire  _GEN_10344 = _T_3 ? _GEN_9695 : _GEN_6382; // @[decode.scala 419:41]
  wire  _GEN_10345 = _T_3 ? _GEN_9696 : _GEN_6383; // @[decode.scala 419:41]
  wire  _GEN_10346 = _T_3 ? _GEN_9697 : _GEN_6384; // @[decode.scala 419:41]
  wire  _GEN_10347 = _T_3 ? _GEN_9698 : _GEN_6385; // @[decode.scala 419:41]
  wire  _GEN_10348 = _T_3 ? _GEN_9699 : _GEN_6386; // @[decode.scala 419:41]
  wire  _GEN_10349 = _T_3 ? _GEN_9700 : _GEN_6387; // @[decode.scala 419:41]
  wire  _GEN_10350 = _T_3 ? _GEN_9701 : _GEN_6388; // @[decode.scala 419:41]
  wire  _GEN_10351 = _T_3 ? _GEN_9702 : _GEN_6389; // @[decode.scala 419:41]
  wire  _GEN_10352 = _T_3 ? _GEN_9703 : _GEN_6390; // @[decode.scala 419:41]
  wire  _GEN_10353 = _T_3 ? _GEN_9704 : _GEN_6391; // @[decode.scala 419:41]
  wire  _GEN_10354 = _T_3 ? _GEN_9705 : _GEN_6392; // @[decode.scala 419:41]
  wire  _GEN_10355 = _T_3 ? _GEN_9706 : _GEN_6393; // @[decode.scala 419:41]
  wire  _GEN_10356 = _T_3 ? _GEN_9707 : _GEN_6394; // @[decode.scala 419:41]
  wire  _GEN_10357 = _T_3 ? _GEN_9708 : _GEN_6395; // @[decode.scala 419:41]
  wire  _GEN_10358 = _T_3 ? _GEN_9709 : _GEN_6396; // @[decode.scala 419:41]
  wire  _GEN_10359 = _T_3 ? _GEN_9710 : _GEN_6397; // @[decode.scala 419:41]
  wire  _GEN_10360 = _T_3 ? _GEN_9711 : _GEN_6398; // @[decode.scala 419:41]
  wire  _GEN_10361 = _T_3 ? _GEN_9712 : _GEN_6399; // @[decode.scala 419:41]
  wire  _GEN_10362 = _T_3 ? _GEN_9713 : _GEN_6400; // @[decode.scala 419:41]
  wire  _GEN_10363 = _T_3 ? _GEN_9714 : _GEN_6401; // @[decode.scala 419:41]
  wire  _GEN_10364 = _T_3 ? _GEN_9715 : _GEN_6402; // @[decode.scala 419:41]
  wire  _GEN_10365 = _T_3 ? _GEN_9716 : _GEN_6403; // @[decode.scala 419:41]
  wire  _GEN_10366 = _T_3 ? _GEN_9717 : _GEN_6404; // @[decode.scala 419:41]
  wire  _GEN_10367 = _T_3 ? _GEN_9718 : _GEN_6405; // @[decode.scala 419:41]
  wire  _GEN_10368 = _T_3 ? _GEN_9719 : _GEN_6406; // @[decode.scala 419:41]
  wire  _GEN_10369 = _T_3 ? _GEN_9720 : _GEN_6407; // @[decode.scala 419:41]
  wire  _GEN_10370 = _T_3 ? _GEN_9721 : _GEN_6408; // @[decode.scala 419:41]
  wire  _GEN_10371 = _T_3 ? _GEN_9722 : _GEN_6409; // @[decode.scala 419:41]
  wire  _GEN_10372 = _T_3 ? _GEN_9723 : _GEN_6410; // @[decode.scala 419:41]
  wire  _GEN_10373 = _T_3 ? _GEN_9724 : _GEN_6411; // @[decode.scala 419:41]
  wire  _GEN_10374 = _T_3 ? _GEN_9725 : _GEN_6412; // @[decode.scala 419:41]
  wire  _GEN_10375 = _T_3 ? _GEN_9726 : _GEN_6413; // @[decode.scala 419:41]
  wire  _GEN_10376 = _T_3 ? _GEN_9727 : _GEN_6414; // @[decode.scala 419:41]
  wire  _GEN_10377 = _T_3 ? _GEN_9728 : _GEN_6415; // @[decode.scala 419:41]
  wire  _GEN_10378 = _T_3 ? _GEN_9729 : _GEN_6416; // @[decode.scala 419:41]
  wire  _GEN_10379 = _T_3 ? _GEN_9730 : _GEN_6417; // @[decode.scala 419:41]
  wire  _GEN_10380 = _T_3 ? _GEN_9731 : _GEN_6418; // @[decode.scala 419:41]
  wire  _GEN_10381 = _T_3 ? _GEN_9732 : _GEN_6419; // @[decode.scala 419:41]
  wire  _GEN_10382 = _T_3 ? _GEN_9733 : _GEN_6420; // @[decode.scala 419:41]
  wire  _GEN_10383 = _T_3 ? _GEN_9734 : _GEN_6421; // @[decode.scala 419:41]
  wire  _GEN_10384 = _T_3 ? _GEN_9735 : _GEN_6422; // @[decode.scala 419:41]
  wire  _GEN_10385 = _T_3 ? _GEN_9736 : _GEN_6423; // @[decode.scala 419:41]
  wire  _GEN_10386 = _T_3 ? _GEN_9737 : _GEN_6424; // @[decode.scala 419:41]
  wire  _GEN_10387 = _T_3 ? _GEN_9738 : _GEN_6425; // @[decode.scala 419:41]
  wire  _GEN_10388 = _T_3 ? _GEN_9739 : _GEN_6426; // @[decode.scala 419:41]
  wire  _GEN_10389 = _T_3 ? _GEN_9740 : _GEN_6427; // @[decode.scala 419:41]
  wire  _GEN_10390 = _T_3 ? _GEN_9741 : _GEN_6428; // @[decode.scala 419:41]
  wire  _GEN_10391 = _T_3 ? _GEN_9742 : _GEN_6429; // @[decode.scala 419:41]
  wire  _GEN_10392 = _T_3 ? _GEN_9743 : _GEN_6430; // @[decode.scala 419:41]
  wire  _GEN_10393 = _T_3 ? _GEN_9744 : _GEN_6431; // @[decode.scala 419:41]
  wire  _GEN_10394 = _T_3 ? _GEN_9745 : _GEN_6432; // @[decode.scala 419:41]
  wire  _GEN_10395 = _T_3 ? _GEN_9746 : _GEN_6433; // @[decode.scala 419:41]
  wire  _GEN_10396 = _T_3 ? _GEN_9747 : _GEN_6434; // @[decode.scala 419:41]
  wire  _GEN_10397 = _T_3 ? _GEN_9748 : _GEN_6435; // @[decode.scala 419:41]
  wire  _GEN_10495 = _T_3 ? _GEN_9846 : _GEN_6437; // @[decode.scala 419:41]
  wire  _GEN_10496 = _T_3 ? _GEN_9847 : _GEN_6438; // @[decode.scala 419:41]
  wire  _GEN_10497 = _T_3 ? _GEN_9848 : _GEN_6439; // @[decode.scala 419:41]
  wire  _GEN_10498 = _T_3 ? _GEN_9849 : _GEN_6440; // @[decode.scala 419:41]
  wire  _GEN_10499 = _T_3 ? _GEN_9850 : _GEN_6441; // @[decode.scala 419:41]
  wire  _GEN_10500 = _T_3 ? _GEN_9851 : _GEN_6442; // @[decode.scala 419:41]
  wire  _GEN_10501 = _T_3 ? _GEN_9852 : _GEN_6443; // @[decode.scala 419:41]
  wire  _GEN_10502 = _T_3 ? _GEN_9853 : _GEN_6444; // @[decode.scala 419:41]
  wire  _GEN_10503 = _T_3 ? _GEN_9854 : _GEN_6445; // @[decode.scala 419:41]
  wire  _GEN_10504 = _T_3 ? _GEN_9855 : _GEN_6446; // @[decode.scala 419:41]
  wire  _GEN_10505 = _T_3 ? _GEN_9856 : _GEN_6447; // @[decode.scala 419:41]
  wire  _GEN_10506 = _T_3 ? _GEN_9857 : _GEN_6448; // @[decode.scala 419:41]
  wire  _GEN_10507 = _T_3 ? _GEN_9858 : _GEN_6449; // @[decode.scala 419:41]
  wire  _GEN_10508 = _T_3 ? _GEN_9859 : _GEN_6450; // @[decode.scala 419:41]
  wire  _GEN_10509 = _T_3 ? _GEN_9860 : _GEN_6451; // @[decode.scala 419:41]
  wire  _GEN_10510 = _T_3 ? _GEN_9861 : _GEN_6452; // @[decode.scala 419:41]
  wire  _GEN_10511 = _T_3 ? _GEN_9862 : _GEN_6453; // @[decode.scala 419:41]
  wire  _GEN_10512 = _T_3 ? _GEN_9863 : _GEN_6454; // @[decode.scala 419:41]
  wire  _GEN_10513 = _T_3 ? _GEN_9864 : _GEN_6455; // @[decode.scala 419:41]
  wire  _GEN_10514 = _T_3 ? _GEN_9865 : _GEN_6456; // @[decode.scala 419:41]
  wire  _GEN_10515 = _T_3 ? _GEN_9866 : _GEN_6457; // @[decode.scala 419:41]
  wire  _GEN_10516 = _T_3 ? _GEN_9867 : _GEN_6458; // @[decode.scala 419:41]
  wire  _GEN_10517 = _T_3 ? _GEN_9868 : _GEN_6459; // @[decode.scala 419:41]
  wire  _GEN_10518 = _T_3 ? _GEN_9869 : _GEN_6460; // @[decode.scala 419:41]
  wire  _GEN_10519 = _T_3 ? _GEN_9870 : _GEN_6461; // @[decode.scala 419:41]
  wire  _GEN_10520 = _T_3 ? _GEN_9871 : _GEN_6462; // @[decode.scala 419:41]
  wire  _GEN_10521 = _T_3 ? _GEN_9872 : _GEN_6463; // @[decode.scala 419:41]
  wire  _GEN_10522 = _T_3 ? _GEN_9873 : _GEN_6464; // @[decode.scala 419:41]
  wire  _GEN_10523 = _T_3 ? _GEN_9874 : _GEN_6465; // @[decode.scala 419:41]
  wire  _GEN_10524 = _T_3 ? _GEN_9875 : _GEN_6466; // @[decode.scala 419:41]
  wire  _GEN_10525 = _T_3 ? _GEN_9876 : _GEN_6467; // @[decode.scala 419:41]
  wire  _GEN_10526 = _T_3 ? _GEN_9877 : _GEN_6468; // @[decode.scala 419:41]
  wire  _GEN_10527 = _T_3 ? _GEN_9878 : _GEN_6469; // @[decode.scala 419:41]
  wire  _GEN_10528 = _T_3 ? _GEN_9879 : _GEN_6470; // @[decode.scala 419:41]
  wire  _GEN_10529 = _T_3 ? _GEN_9880 : _GEN_6471; // @[decode.scala 419:41]
  wire  _GEN_10530 = _T_3 ? _GEN_9881 : _GEN_6472; // @[decode.scala 419:41]
  wire  _GEN_10531 = _T_3 ? _GEN_9882 : _GEN_6473; // @[decode.scala 419:41]
  wire  _GEN_10532 = _T_3 ? _GEN_9883 : _GEN_6474; // @[decode.scala 419:41]
  wire  _GEN_10533 = _T_3 ? _GEN_9884 : _GEN_6475; // @[decode.scala 419:41]
  wire  _GEN_10534 = _T_3 ? _GEN_9885 : _GEN_6476; // @[decode.scala 419:41]
  wire  _GEN_10535 = _T_3 ? _GEN_9886 : _GEN_6477; // @[decode.scala 419:41]
  wire  _GEN_10536 = _T_3 ? _GEN_9887 : _GEN_6478; // @[decode.scala 419:41]
  wire  _GEN_10537 = _T_3 ? _GEN_9888 : _GEN_6479; // @[decode.scala 419:41]
  wire  _GEN_10538 = _T_3 ? _GEN_9889 : _GEN_6480; // @[decode.scala 419:41]
  wire  _GEN_10539 = _T_3 ? _GEN_9890 : _GEN_6481; // @[decode.scala 419:41]
  wire  _GEN_10540 = _T_3 ? _GEN_9891 : _GEN_6482; // @[decode.scala 419:41]
  wire  _GEN_10541 = _T_3 ? _GEN_9892 : _GEN_6483; // @[decode.scala 419:41]
  wire  _GEN_10542 = _T_3 ? _GEN_9893 : _GEN_6484; // @[decode.scala 419:41]
  wire  _GEN_10543 = _T_3 ? _GEN_9894 : _GEN_6485; // @[decode.scala 419:41]
  wire  _GEN_10544 = _T_3 ? _GEN_9895 : _GEN_6486; // @[decode.scala 419:41]
  wire  _GEN_10545 = _T_3 ? _GEN_9896 : _GEN_6487; // @[decode.scala 419:41]
  wire  _GEN_10546 = _T_3 ? _GEN_9897 : _GEN_6488; // @[decode.scala 419:41]
  wire  _GEN_10547 = _T_3 ? _GEN_9898 : _GEN_6489; // @[decode.scala 419:41]
  wire  _GEN_10548 = _T_3 ? _GEN_9899 : _GEN_6490; // @[decode.scala 419:41]
  wire  _GEN_10549 = _T_3 ? _GEN_9900 : _GEN_6491; // @[decode.scala 419:41]
  wire  _GEN_10550 = _T_3 ? _GEN_9901 : _GEN_6492; // @[decode.scala 419:41]
  wire  _GEN_10551 = _T_3 ? _GEN_9902 : _GEN_6493; // @[decode.scala 419:41]
  wire  _GEN_10552 = _T_3 ? _GEN_9903 : _GEN_6494; // @[decode.scala 419:41]
  wire  _GEN_10553 = _T_3 ? _GEN_9904 : _GEN_6495; // @[decode.scala 419:41]
  wire  _GEN_10554 = _T_3 ? _GEN_9905 : _GEN_6496; // @[decode.scala 419:41]
  wire  _GEN_10555 = _T_3 ? _GEN_9906 : _GEN_6497; // @[decode.scala 419:41]
  wire  _GEN_10556 = _T_3 ? _GEN_9907 : _GEN_6498; // @[decode.scala 419:41]
  wire  _GEN_10557 = _T_3 ? _GEN_9908 : _GEN_6499; // @[decode.scala 419:41]
  wire  _GEN_10655 = _T_3 ? _GEN_10006 : _GEN_6501; // @[decode.scala 419:41]
  wire  _GEN_10656 = _T_3 ? _GEN_10007 : _GEN_6502; // @[decode.scala 419:41]
  wire  _GEN_10657 = _T_3 ? _GEN_10008 : _GEN_6503; // @[decode.scala 419:41]
  wire  _GEN_10658 = _T_3 ? _GEN_10009 : _GEN_6504; // @[decode.scala 419:41]
  wire  _GEN_10659 = _T_3 ? _GEN_10010 : _GEN_6505; // @[decode.scala 419:41]
  wire  _GEN_10660 = _T_3 ? _GEN_10011 : _GEN_6506; // @[decode.scala 419:41]
  wire  _GEN_10661 = _T_3 ? _GEN_10012 : _GEN_6507; // @[decode.scala 419:41]
  wire  _GEN_10662 = _T_3 ? _GEN_10013 : _GEN_6508; // @[decode.scala 419:41]
  wire  _GEN_10663 = _T_3 ? _GEN_10014 : _GEN_6509; // @[decode.scala 419:41]
  wire  _GEN_10664 = _T_3 ? _GEN_10015 : _GEN_6510; // @[decode.scala 419:41]
  wire  _GEN_10665 = _T_3 ? _GEN_10016 : _GEN_6511; // @[decode.scala 419:41]
  wire  _GEN_10666 = _T_3 ? _GEN_10017 : _GEN_6512; // @[decode.scala 419:41]
  wire  _GEN_10667 = _T_3 ? _GEN_10018 : _GEN_6513; // @[decode.scala 419:41]
  wire  _GEN_10668 = _T_3 ? _GEN_10019 : _GEN_6514; // @[decode.scala 419:41]
  wire  _GEN_10669 = _T_3 ? _GEN_10020 : _GEN_6515; // @[decode.scala 419:41]
  wire  _GEN_10670 = _T_3 ? _GEN_10021 : _GEN_6516; // @[decode.scala 419:41]
  wire  _GEN_10671 = _T_3 ? _GEN_10022 : _GEN_6517; // @[decode.scala 419:41]
  wire  _GEN_10672 = _T_3 ? _GEN_10023 : _GEN_6518; // @[decode.scala 419:41]
  wire  _GEN_10673 = _T_3 ? _GEN_10024 : _GEN_6519; // @[decode.scala 419:41]
  wire  _GEN_10674 = _T_3 ? _GEN_10025 : _GEN_6520; // @[decode.scala 419:41]
  wire  _GEN_10675 = _T_3 ? _GEN_10026 : _GEN_6521; // @[decode.scala 419:41]
  wire  _GEN_10676 = _T_3 ? _GEN_10027 : _GEN_6522; // @[decode.scala 419:41]
  wire  _GEN_10677 = _T_3 ? _GEN_10028 : _GEN_6523; // @[decode.scala 419:41]
  wire  _GEN_10678 = _T_3 ? _GEN_10029 : _GEN_6524; // @[decode.scala 419:41]
  wire  _GEN_10679 = _T_3 ? _GEN_10030 : _GEN_6525; // @[decode.scala 419:41]
  wire  _GEN_10680 = _T_3 ? _GEN_10031 : _GEN_6526; // @[decode.scala 419:41]
  wire  _GEN_10681 = _T_3 ? _GEN_10032 : _GEN_6527; // @[decode.scala 419:41]
  wire  _GEN_10682 = _T_3 ? _GEN_10033 : _GEN_6528; // @[decode.scala 419:41]
  wire  _GEN_10683 = _T_3 ? _GEN_10034 : _GEN_6529; // @[decode.scala 419:41]
  wire  _GEN_10684 = _T_3 ? _GEN_10035 : _GEN_6530; // @[decode.scala 419:41]
  wire  _GEN_10685 = _T_3 ? _GEN_10036 : _GEN_6531; // @[decode.scala 419:41]
  wire  _GEN_10686 = _T_3 ? _GEN_10037 : _GEN_6532; // @[decode.scala 419:41]
  wire  _GEN_10687 = _T_3 ? _GEN_10038 : _GEN_6533; // @[decode.scala 419:41]
  wire  _GEN_10688 = _T_3 ? _GEN_10039 : _GEN_6534; // @[decode.scala 419:41]
  wire  _GEN_10689 = _T_3 ? _GEN_10040 : _GEN_6535; // @[decode.scala 419:41]
  wire  _GEN_10690 = _T_3 ? _GEN_10041 : _GEN_6536; // @[decode.scala 419:41]
  wire  _GEN_10691 = _T_3 ? _GEN_10042 : _GEN_6537; // @[decode.scala 419:41]
  wire  _GEN_10692 = _T_3 ? _GEN_10043 : _GEN_6538; // @[decode.scala 419:41]
  wire  _GEN_10693 = _T_3 ? _GEN_10044 : _GEN_6539; // @[decode.scala 419:41]
  wire  _GEN_10694 = _T_3 ? _GEN_10045 : _GEN_6540; // @[decode.scala 419:41]
  wire  _GEN_10695 = _T_3 ? _GEN_10046 : _GEN_6541; // @[decode.scala 419:41]
  wire  _GEN_10696 = _T_3 ? _GEN_10047 : _GEN_6542; // @[decode.scala 419:41]
  wire  _GEN_10697 = _T_3 ? _GEN_10048 : _GEN_6543; // @[decode.scala 419:41]
  wire  _GEN_10698 = _T_3 ? _GEN_10049 : _GEN_6544; // @[decode.scala 419:41]
  wire  _GEN_10699 = _T_3 ? _GEN_10050 : _GEN_6545; // @[decode.scala 419:41]
  wire  _GEN_10700 = _T_3 ? _GEN_10051 : _GEN_6546; // @[decode.scala 419:41]
  wire  _GEN_10701 = _T_3 ? _GEN_10052 : _GEN_6547; // @[decode.scala 419:41]
  wire  _GEN_10702 = _T_3 ? _GEN_10053 : _GEN_6548; // @[decode.scala 419:41]
  wire  _GEN_10703 = _T_3 ? _GEN_10054 : _GEN_6549; // @[decode.scala 419:41]
  wire  _GEN_10704 = _T_3 ? _GEN_10055 : _GEN_6550; // @[decode.scala 419:41]
  wire  _GEN_10705 = _T_3 ? _GEN_10056 : _GEN_6551; // @[decode.scala 419:41]
  wire  _GEN_10706 = _T_3 ? _GEN_10057 : _GEN_6552; // @[decode.scala 419:41]
  wire  _GEN_10707 = _T_3 ? _GEN_10058 : _GEN_6553; // @[decode.scala 419:41]
  wire  _GEN_10708 = _T_3 ? _GEN_10059 : _GEN_6554; // @[decode.scala 419:41]
  wire  _GEN_10709 = _T_3 ? _GEN_10060 : _GEN_6555; // @[decode.scala 419:41]
  wire  _GEN_10710 = _T_3 ? _GEN_10061 : _GEN_6556; // @[decode.scala 419:41]
  wire  _GEN_10711 = _T_3 ? _GEN_10062 : _GEN_6557; // @[decode.scala 419:41]
  wire  _GEN_10712 = _T_3 ? _GEN_10063 : _GEN_6558; // @[decode.scala 419:41]
  wire  _GEN_10713 = _T_3 ? _GEN_10064 : _GEN_6559; // @[decode.scala 419:41]
  wire  _GEN_10714 = _T_3 ? _GEN_10065 : _GEN_6560; // @[decode.scala 419:41]
  wire  _GEN_10715 = _T_3 ? _GEN_10066 : _GEN_6561; // @[decode.scala 419:41]
  wire  _GEN_10716 = _T_3 ? _GEN_10067 : _GEN_6562; // @[decode.scala 419:41]
  wire  _GEN_10717 = _T_3 ? _GEN_10068 : _GEN_6563; // @[decode.scala 419:41]
  wire  _GEN_10815 = _T_3 ? _GEN_10166 : reservedFreeList4_0; // @[decode.scala 325:30 419:41]
  wire  _GEN_10816 = _T_3 ? _GEN_10167 : reservedFreeList4_1; // @[decode.scala 325:30 419:41]
  wire  _GEN_10817 = _T_3 ? _GEN_10168 : reservedFreeList4_2; // @[decode.scala 325:30 419:41]
  wire  _GEN_10818 = _T_3 ? _GEN_10169 : reservedFreeList4_3; // @[decode.scala 325:30 419:41]
  wire  _GEN_10819 = _T_3 ? _GEN_10170 : reservedFreeList4_4; // @[decode.scala 325:30 419:41]
  wire  _GEN_10820 = _T_3 ? _GEN_10171 : reservedFreeList4_5; // @[decode.scala 325:30 419:41]
  wire  _GEN_10821 = _T_3 ? _GEN_10172 : reservedFreeList4_6; // @[decode.scala 325:30 419:41]
  wire  _GEN_10822 = _T_3 ? _GEN_10173 : reservedFreeList4_7; // @[decode.scala 325:30 419:41]
  wire  _GEN_10823 = _T_3 ? _GEN_10174 : reservedFreeList4_8; // @[decode.scala 325:30 419:41]
  wire  _GEN_10824 = _T_3 ? _GEN_10175 : reservedFreeList4_9; // @[decode.scala 325:30 419:41]
  wire  _GEN_10825 = _T_3 ? _GEN_10176 : reservedFreeList4_10; // @[decode.scala 325:30 419:41]
  wire  _GEN_10826 = _T_3 ? _GEN_10177 : reservedFreeList4_11; // @[decode.scala 325:30 419:41]
  wire  _GEN_10827 = _T_3 ? _GEN_10178 : reservedFreeList4_12; // @[decode.scala 325:30 419:41]
  wire  _GEN_10828 = _T_3 ? _GEN_10179 : reservedFreeList4_13; // @[decode.scala 325:30 419:41]
  wire  _GEN_10829 = _T_3 ? _GEN_10180 : reservedFreeList4_14; // @[decode.scala 325:30 419:41]
  wire  _GEN_10830 = _T_3 ? _GEN_10181 : reservedFreeList4_15; // @[decode.scala 325:30 419:41]
  wire  _GEN_10831 = _T_3 ? _GEN_10182 : reservedFreeList4_16; // @[decode.scala 325:30 419:41]
  wire  _GEN_10832 = _T_3 ? _GEN_10183 : reservedFreeList4_17; // @[decode.scala 325:30 419:41]
  wire  _GEN_10833 = _T_3 ? _GEN_10184 : reservedFreeList4_18; // @[decode.scala 325:30 419:41]
  wire  _GEN_10834 = _T_3 ? _GEN_10185 : reservedFreeList4_19; // @[decode.scala 325:30 419:41]
  wire  _GEN_10835 = _T_3 ? _GEN_10186 : reservedFreeList4_20; // @[decode.scala 325:30 419:41]
  wire  _GEN_10836 = _T_3 ? _GEN_10187 : reservedFreeList4_21; // @[decode.scala 325:30 419:41]
  wire  _GEN_10837 = _T_3 ? _GEN_10188 : reservedFreeList4_22; // @[decode.scala 325:30 419:41]
  wire  _GEN_10838 = _T_3 ? _GEN_10189 : reservedFreeList4_23; // @[decode.scala 325:30 419:41]
  wire  _GEN_10839 = _T_3 ? _GEN_10190 : reservedFreeList4_24; // @[decode.scala 325:30 419:41]
  wire  _GEN_10840 = _T_3 ? _GEN_10191 : reservedFreeList4_25; // @[decode.scala 325:30 419:41]
  wire  _GEN_10841 = _T_3 ? _GEN_10192 : reservedFreeList4_26; // @[decode.scala 325:30 419:41]
  wire  _GEN_10842 = _T_3 ? _GEN_10193 : reservedFreeList4_27; // @[decode.scala 325:30 419:41]
  wire  _GEN_10843 = _T_3 ? _GEN_10194 : reservedFreeList4_28; // @[decode.scala 325:30 419:41]
  wire  _GEN_10844 = _T_3 ? _GEN_10195 : reservedFreeList4_29; // @[decode.scala 325:30 419:41]
  wire  _GEN_10845 = _T_3 ? _GEN_10196 : reservedFreeList4_30; // @[decode.scala 325:30 419:41]
  wire  _GEN_10846 = _T_3 ? _GEN_10197 : reservedFreeList4_31; // @[decode.scala 325:30 419:41]
  wire  _GEN_10847 = _T_3 ? _GEN_10198 : reservedFreeList4_32; // @[decode.scala 325:30 419:41]
  wire  _GEN_10848 = _T_3 ? _GEN_10199 : reservedFreeList4_33; // @[decode.scala 325:30 419:41]
  wire  _GEN_10849 = _T_3 ? _GEN_10200 : reservedFreeList4_34; // @[decode.scala 325:30 419:41]
  wire  _GEN_10850 = _T_3 ? _GEN_10201 : reservedFreeList4_35; // @[decode.scala 325:30 419:41]
  wire  _GEN_10851 = _T_3 ? _GEN_10202 : reservedFreeList4_36; // @[decode.scala 325:30 419:41]
  wire  _GEN_10852 = _T_3 ? _GEN_10203 : reservedFreeList4_37; // @[decode.scala 325:30 419:41]
  wire  _GEN_10853 = _T_3 ? _GEN_10204 : reservedFreeList4_38; // @[decode.scala 325:30 419:41]
  wire  _GEN_10854 = _T_3 ? _GEN_10205 : reservedFreeList4_39; // @[decode.scala 325:30 419:41]
  wire  _GEN_10855 = _T_3 ? _GEN_10206 : reservedFreeList4_40; // @[decode.scala 325:30 419:41]
  wire  _GEN_10856 = _T_3 ? _GEN_10207 : reservedFreeList4_41; // @[decode.scala 325:30 419:41]
  wire  _GEN_10857 = _T_3 ? _GEN_10208 : reservedFreeList4_42; // @[decode.scala 325:30 419:41]
  wire  _GEN_10858 = _T_3 ? _GEN_10209 : reservedFreeList4_43; // @[decode.scala 325:30 419:41]
  wire  _GEN_10859 = _T_3 ? _GEN_10210 : reservedFreeList4_44; // @[decode.scala 325:30 419:41]
  wire  _GEN_10860 = _T_3 ? _GEN_10211 : reservedFreeList4_45; // @[decode.scala 325:30 419:41]
  wire  _GEN_10861 = _T_3 ? _GEN_10212 : reservedFreeList4_46; // @[decode.scala 325:30 419:41]
  wire  _GEN_10862 = _T_3 ? _GEN_10213 : reservedFreeList4_47; // @[decode.scala 325:30 419:41]
  wire  _GEN_10863 = _T_3 ? _GEN_10214 : reservedFreeList4_48; // @[decode.scala 325:30 419:41]
  wire  _GEN_10864 = _T_3 ? _GEN_10215 : reservedFreeList4_49; // @[decode.scala 325:30 419:41]
  wire  _GEN_10865 = _T_3 ? _GEN_10216 : reservedFreeList4_50; // @[decode.scala 325:30 419:41]
  wire  _GEN_10866 = _T_3 ? _GEN_10217 : reservedFreeList4_51; // @[decode.scala 325:30 419:41]
  wire  _GEN_10867 = _T_3 ? _GEN_10218 : reservedFreeList4_52; // @[decode.scala 325:30 419:41]
  wire  _GEN_10868 = _T_3 ? _GEN_10219 : reservedFreeList4_53; // @[decode.scala 325:30 419:41]
  wire  _GEN_10869 = _T_3 ? _GEN_10220 : reservedFreeList4_54; // @[decode.scala 325:30 419:41]
  wire  _GEN_10870 = _T_3 ? _GEN_10221 : reservedFreeList4_55; // @[decode.scala 325:30 419:41]
  wire  _GEN_10871 = _T_3 ? _GEN_10222 : reservedFreeList4_56; // @[decode.scala 325:30 419:41]
  wire  _GEN_10872 = _T_3 ? _GEN_10223 : reservedFreeList4_57; // @[decode.scala 325:30 419:41]
  wire  _GEN_10873 = _T_3 ? _GEN_10224 : reservedFreeList4_58; // @[decode.scala 325:30 419:41]
  wire  _GEN_10874 = _T_3 ? _GEN_10225 : reservedFreeList4_59; // @[decode.scala 325:30 419:41]
  wire  _GEN_10875 = _T_3 ? _GEN_10226 : reservedFreeList4_60; // @[decode.scala 325:30 419:41]
  wire  _GEN_10876 = _T_3 ? _GEN_10227 : reservedFreeList4_61; // @[decode.scala 325:30 419:41]
  wire  _GEN_10877 = _T_3 ? _GEN_10228 : reservedFreeList4_62; // @[decode.scala 325:30 419:41]
  wire  _T_222 = fromFetch_expected_pc == fromFetch_pc; // @[decode.scala 487:71]
  wire [63:0] _GEN_10945 = _fromFetch_expected_valid_T & fromFetch_fired & fromFetch_expected_pc == fromFetch_pc ? 64'h0
     : _GEN_6115; // @[decode.scala 487:89 488:16]
  wire  isCSR = csrIns & toExec_fired; // @[decode.scala 495:98]
  reg [63:0] ustatus; // @[decode.scala 497:28]
  reg [63:0] utvec; // @[decode.scala 498:28]
  reg [63:0] uepc; // @[decode.scala 499:28]
  reg [63:0] ucause; // @[decode.scala 500:28]
  reg [63:0] scounteren; // @[decode.scala 501:28]
  reg [63:0] satp; // @[decode.scala 502:28]
  reg [63:0] mstatus; // @[decode.scala 503:28]
  reg [63:0] misa; // @[decode.scala 504:28]
  reg [63:0] medeleg; // @[decode.scala 505:28]
  reg [63:0] mideleg; // @[decode.scala 506:28]
  reg [63:0] mie; // @[decode.scala 507:28]
  reg [63:0] mtvec; // @[decode.scala 508:28]
  reg [63:0] mcounteren; // @[decode.scala 509:28]
  reg [63:0] mscratch; // @[decode.scala 510:28]
  reg [63:0] mepc; // @[decode.scala 511:28]
  reg [63:0] mcause; // @[decode.scala 512:28]
  reg [63:0] mtval; // @[decode.scala 513:28]
  reg [63:0] mip; // @[decode.scala 514:28]
  reg [63:0] pmpcfg0; // @[decode.scala 515:28]
  reg [63:0] pmpaddr0; // @[decode.scala 516:28]
  reg [63:0] mvendorid; // @[decode.scala 517:28]
  reg [63:0] marchid; // @[decode.scala 518:28]
  reg [63:0] mimpid; // @[decode.scala 519:28]
  reg [63:0] mhartid; // @[decode.scala 520:28]
  wire [63:0] _mstatus_T = mstatus & 64'h1888; // @[decode.scala 522:23]
  wire [63:0] _mstatus_T_1 = _mstatus_T | 64'ha00000000; // @[decode.scala 522:48]
  wire [63:0] _GEN_10951 = isCSR ? outputBuffer_immediate : {{52'd0}, csrAddrReg}; // @[decode.scala 525:15 528:19 242:27]
  wire  _T_224 = opcode == 7'h73; // @[decode.scala 534:15]
  wire [63:0] _T_229 = immediate_immediate & 64'hfff; // @[decode.scala 535:22]
  wire [63:0] _GEN_10954 = 64'hf14 == _T_229 ? mhartid : csrReadDataReg; // @[decode.scala 240:31 535:34 559:37]
  wire [63:0] _GEN_10955 = 64'hf13 == _T_229 ? mimpid : _GEN_10954; // @[decode.scala 535:34 558:37]
  wire [63:0] _GEN_10956 = 64'hf12 == _T_229 ? marchid : _GEN_10955; // @[decode.scala 535:34 557:37]
  wire [63:0] _GEN_10957 = 64'hf11 == _T_229 ? mvendorid : _GEN_10956; // @[decode.scala 535:34 556:37]
  wire [63:0] _GEN_10958 = 64'h3b0 == _T_229 ? pmpaddr0 : _GEN_10957; // @[decode.scala 535:34 555:37]
  wire [63:0] _GEN_10959 = 64'h3a0 == _T_229 ? pmpcfg0 : _GEN_10958; // @[decode.scala 535:34 554:37]
  wire [63:0] _GEN_10960 = 64'h344 == _T_229 ? mip : _GEN_10959; // @[decode.scala 535:34 553:37]
  wire [63:0] _GEN_10961 = 64'h343 == _T_229 ? mtval : _GEN_10960; // @[decode.scala 535:34 552:37]
  wire [63:0] _GEN_10962 = 64'h342 == _T_229 ? mcause : _GEN_10961; // @[decode.scala 535:34 551:37]
  wire [63:0] _GEN_10963 = 64'h341 == _T_229 ? mepc : _GEN_10962; // @[decode.scala 535:34 550:37]
  wire [63:0] _GEN_10964 = 64'h340 == _T_229 ? mscratch : _GEN_10963; // @[decode.scala 535:34 549:37]
  wire [63:0] _GEN_10965 = 64'h306 == _T_229 ? mcounteren : _GEN_10964; // @[decode.scala 535:34 548:37]
  wire [63:0] _GEN_10966 = 64'h305 == _T_229 ? mtvec : _GEN_10965; // @[decode.scala 535:34 547:37]
  wire [63:0] _GEN_10967 = 64'h304 == _T_229 ? mie : _GEN_10966; // @[decode.scala 535:34 546:37]
  wire [63:0] _GEN_10968 = 64'h303 == _T_229 ? mideleg : _GEN_10967; // @[decode.scala 535:34 545:37]
  wire [63:0] _GEN_10969 = 64'h302 == _T_229 ? medeleg : _GEN_10968; // @[decode.scala 535:34 544:37]
  wire [63:0] _GEN_10970 = 64'h301 == _T_229 ? misa : _GEN_10969; // @[decode.scala 535:34 543:37]
  wire [63:0] _GEN_10971 = 64'h300 == _T_229 ? mstatus : _GEN_10970; // @[decode.scala 535:34 542:37]
  wire [63:0] _GEN_10972 = 64'h180 == _T_229 ? satp : _GEN_10971; // @[decode.scala 535:34 541:37]
  wire [63:0] _GEN_10973 = 64'h106 == _T_229 ? scounteren : _GEN_10972; // @[decode.scala 535:34 540:37]
  wire [63:0] _GEN_10974 = 64'h42 == _T_229 ? ucause : _GEN_10973; // @[decode.scala 535:34 539:37]
  wire [63:0] _GEN_10975 = 64'h41 == _T_229 ? uepc : _GEN_10974; // @[decode.scala 535:34 538:37]
  wire  _T_256 = writeBackResult_fired & writeBackResult_instruction[6:0] == 7'h73; // @[decode.scala 564:30]
  wire  _GEN_10979 = writeBackResult_fired & writeBackResult_instruction[6:0] == 7'h73 ? 1'h0 : _GEN_4; // @[decode.scala 564:80 565:14]
  wire  _T_266 = 12'h0 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_267 = 12'h5 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_268 = 12'h41 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_269 = 12'h42 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_270 = 12'h106 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_271 = 12'h180 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_272 = 12'h300 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_273 = 12'h301 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_274 = 12'h302 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_275 = 12'h303 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_276 = 12'h304 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_277 = 12'h305 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_278 = 12'h306 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_279 = 12'h340 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_280 = 12'h341 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_281 = 12'h342 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_282 = 12'h343 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_283 = 12'h344 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_284 = 12'h3a0 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_285 = 12'h3b0 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_286 = 12'hf11 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_287 = 12'hf12 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_288 = 12'hf13 == csrAddrReg; // @[decode.scala 573:39]
  wire  _T_289 = 12'hf14 == csrAddrReg; // @[decode.scala 573:39]
  wire [63:0] csrWriteData = _T_256 & writeBackResult_instruction[14:12] != 3'h0 ? writeBackResult_data : 64'h0; // @[decode.scala 568:126 570:18]
  wire [63:0] _GEN_10980 = 12'hf14 == csrAddrReg ? csrWriteData : mhartid; // @[decode.scala 520:28 573:39 597:37]
  wire [63:0] _GEN_10981 = 12'hf13 == csrAddrReg ? csrWriteData : mimpid; // @[decode.scala 519:28 573:39 596:37]
  wire [63:0] _GEN_10982 = 12'hf13 == csrAddrReg ? mhartid : _GEN_10980; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_10983 = 12'hf12 == csrAddrReg ? csrWriteData : marchid; // @[decode.scala 518:28 573:39 595:37]
  wire [63:0] _GEN_10984 = 12'hf12 == csrAddrReg ? mimpid : _GEN_10981; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_10985 = 12'hf12 == csrAddrReg ? mhartid : _GEN_10982; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_10986 = 12'hf11 == csrAddrReg ? csrWriteData : mvendorid; // @[decode.scala 517:28 573:39 594:37]
  wire [63:0] _GEN_10987 = 12'hf11 == csrAddrReg ? marchid : _GEN_10983; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_10988 = 12'hf11 == csrAddrReg ? mimpid : _GEN_10984; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_10989 = 12'hf11 == csrAddrReg ? mhartid : _GEN_10985; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_10990 = 12'h3b0 == csrAddrReg ? csrWriteData : pmpaddr0; // @[decode.scala 516:28 573:39 593:37]
  wire [63:0] _GEN_10991 = 12'h3b0 == csrAddrReg ? mvendorid : _GEN_10986; // @[decode.scala 517:28 573:39]
  wire [63:0] _GEN_10992 = 12'h3b0 == csrAddrReg ? marchid : _GEN_10987; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_10993 = 12'h3b0 == csrAddrReg ? mimpid : _GEN_10988; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_10994 = 12'h3b0 == csrAddrReg ? mhartid : _GEN_10989; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_10995 = 12'h3a0 == csrAddrReg ? csrWriteData : pmpcfg0; // @[decode.scala 515:28 573:39 592:37]
  wire [63:0] _GEN_10996 = 12'h3a0 == csrAddrReg ? pmpaddr0 : _GEN_10990; // @[decode.scala 516:28 573:39]
  wire [63:0] _GEN_10997 = 12'h3a0 == csrAddrReg ? mvendorid : _GEN_10991; // @[decode.scala 517:28 573:39]
  wire [63:0] _GEN_10998 = 12'h3a0 == csrAddrReg ? marchid : _GEN_10992; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_10999 = 12'h3a0 == csrAddrReg ? mimpid : _GEN_10993; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_11000 = 12'h3a0 == csrAddrReg ? mhartid : _GEN_10994; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_11001 = 12'h344 == csrAddrReg ? csrWriteData : mip; // @[decode.scala 514:28 573:39 591:37]
  wire [63:0] _GEN_11002 = 12'h344 == csrAddrReg ? pmpcfg0 : _GEN_10995; // @[decode.scala 515:28 573:39]
  wire [63:0] _GEN_11003 = 12'h344 == csrAddrReg ? pmpaddr0 : _GEN_10996; // @[decode.scala 516:28 573:39]
  wire [63:0] _GEN_11004 = 12'h344 == csrAddrReg ? mvendorid : _GEN_10997; // @[decode.scala 517:28 573:39]
  wire [63:0] _GEN_11005 = 12'h344 == csrAddrReg ? marchid : _GEN_10998; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_11006 = 12'h344 == csrAddrReg ? mimpid : _GEN_10999; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_11007 = 12'h344 == csrAddrReg ? mhartid : _GEN_11000; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_11008 = 12'h343 == csrAddrReg ? csrWriteData : mtval; // @[decode.scala 513:28 573:39 590:37]
  wire [63:0] _GEN_11009 = 12'h343 == csrAddrReg ? mip : _GEN_11001; // @[decode.scala 514:28 573:39]
  wire [63:0] _GEN_11010 = 12'h343 == csrAddrReg ? pmpcfg0 : _GEN_11002; // @[decode.scala 515:28 573:39]
  wire [63:0] _GEN_11011 = 12'h343 == csrAddrReg ? pmpaddr0 : _GEN_11003; // @[decode.scala 516:28 573:39]
  wire [63:0] _GEN_11012 = 12'h343 == csrAddrReg ? mvendorid : _GEN_11004; // @[decode.scala 517:28 573:39]
  wire [63:0] _GEN_11013 = 12'h343 == csrAddrReg ? marchid : _GEN_11005; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_11014 = 12'h343 == csrAddrReg ? mimpid : _GEN_11006; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_11015 = 12'h343 == csrAddrReg ? mhartid : _GEN_11007; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_11016 = 12'h342 == csrAddrReg ? csrWriteData : mcause; // @[decode.scala 512:28 573:39 589:37]
  wire [63:0] _GEN_11017 = 12'h342 == csrAddrReg ? mtval : _GEN_11008; // @[decode.scala 513:28 573:39]
  wire [63:0] _GEN_11018 = 12'h342 == csrAddrReg ? mip : _GEN_11009; // @[decode.scala 514:28 573:39]
  wire [63:0] _GEN_11019 = 12'h342 == csrAddrReg ? pmpcfg0 : _GEN_11010; // @[decode.scala 515:28 573:39]
  wire [63:0] _GEN_11020 = 12'h342 == csrAddrReg ? pmpaddr0 : _GEN_11011; // @[decode.scala 516:28 573:39]
  wire [63:0] _GEN_11021 = 12'h342 == csrAddrReg ? mvendorid : _GEN_11012; // @[decode.scala 517:28 573:39]
  wire [63:0] _GEN_11022 = 12'h342 == csrAddrReg ? marchid : _GEN_11013; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_11023 = 12'h342 == csrAddrReg ? mimpid : _GEN_11014; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_11024 = 12'h342 == csrAddrReg ? mhartid : _GEN_11015; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_11025 = 12'h341 == csrAddrReg ? csrWriteData : mepc; // @[decode.scala 511:28 573:39 588:37]
  wire [63:0] _GEN_11026 = 12'h341 == csrAddrReg ? mcause : _GEN_11016; // @[decode.scala 512:28 573:39]
  wire [63:0] _GEN_11027 = 12'h341 == csrAddrReg ? mtval : _GEN_11017; // @[decode.scala 513:28 573:39]
  wire [63:0] _GEN_11028 = 12'h341 == csrAddrReg ? mip : _GEN_11018; // @[decode.scala 514:28 573:39]
  wire [63:0] _GEN_11029 = 12'h341 == csrAddrReg ? pmpcfg0 : _GEN_11019; // @[decode.scala 515:28 573:39]
  wire [63:0] _GEN_11030 = 12'h341 == csrAddrReg ? pmpaddr0 : _GEN_11020; // @[decode.scala 516:28 573:39]
  wire [63:0] _GEN_11031 = 12'h341 == csrAddrReg ? mvendorid : _GEN_11021; // @[decode.scala 517:28 573:39]
  wire [63:0] _GEN_11032 = 12'h341 == csrAddrReg ? marchid : _GEN_11022; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_11033 = 12'h341 == csrAddrReg ? mimpid : _GEN_11023; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_11034 = 12'h341 == csrAddrReg ? mhartid : _GEN_11024; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_11035 = 12'h340 == csrAddrReg ? csrWriteData : mscratch; // @[decode.scala 510:28 573:39 587:37]
  wire [63:0] _GEN_11036 = 12'h340 == csrAddrReg ? mepc : _GEN_11025; // @[decode.scala 511:28 573:39]
  wire [63:0] _GEN_11037 = 12'h340 == csrAddrReg ? mcause : _GEN_11026; // @[decode.scala 512:28 573:39]
  wire [63:0] _GEN_11038 = 12'h340 == csrAddrReg ? mtval : _GEN_11027; // @[decode.scala 513:28 573:39]
  wire [63:0] _GEN_11039 = 12'h340 == csrAddrReg ? mip : _GEN_11028; // @[decode.scala 514:28 573:39]
  wire [63:0] _GEN_11040 = 12'h340 == csrAddrReg ? pmpcfg0 : _GEN_11029; // @[decode.scala 515:28 573:39]
  wire [63:0] _GEN_11041 = 12'h340 == csrAddrReg ? pmpaddr0 : _GEN_11030; // @[decode.scala 516:28 573:39]
  wire [63:0] _GEN_11042 = 12'h340 == csrAddrReg ? mvendorid : _GEN_11031; // @[decode.scala 517:28 573:39]
  wire [63:0] _GEN_11043 = 12'h340 == csrAddrReg ? marchid : _GEN_11032; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_11044 = 12'h340 == csrAddrReg ? mimpid : _GEN_11033; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_11045 = 12'h340 == csrAddrReg ? mhartid : _GEN_11034; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_11046 = 12'h306 == csrAddrReg ? csrWriteData : mcounteren; // @[decode.scala 509:28 573:39 586:37]
  wire [63:0] _GEN_11047 = 12'h306 == csrAddrReg ? mscratch : _GEN_11035; // @[decode.scala 510:28 573:39]
  wire [63:0] _GEN_11048 = 12'h306 == csrAddrReg ? mepc : _GEN_11036; // @[decode.scala 511:28 573:39]
  wire [63:0] _GEN_11049 = 12'h306 == csrAddrReg ? mcause : _GEN_11037; // @[decode.scala 512:28 573:39]
  wire [63:0] _GEN_11050 = 12'h306 == csrAddrReg ? mtval : _GEN_11038; // @[decode.scala 513:28 573:39]
  wire [63:0] _GEN_11051 = 12'h306 == csrAddrReg ? mip : _GEN_11039; // @[decode.scala 514:28 573:39]
  wire [63:0] _GEN_11052 = 12'h306 == csrAddrReg ? pmpcfg0 : _GEN_11040; // @[decode.scala 515:28 573:39]
  wire [63:0] _GEN_11053 = 12'h306 == csrAddrReg ? pmpaddr0 : _GEN_11041; // @[decode.scala 516:28 573:39]
  wire [63:0] _GEN_11054 = 12'h306 == csrAddrReg ? mvendorid : _GEN_11042; // @[decode.scala 517:28 573:39]
  wire [63:0] _GEN_11055 = 12'h306 == csrAddrReg ? marchid : _GEN_11043; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_11056 = 12'h306 == csrAddrReg ? mimpid : _GEN_11044; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_11057 = 12'h306 == csrAddrReg ? mhartid : _GEN_11045; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_11058 = 12'h305 == csrAddrReg ? csrWriteData : mtvec; // @[decode.scala 508:28 573:39 585:37]
  wire [63:0] _GEN_11059 = 12'h305 == csrAddrReg ? mcounteren : _GEN_11046; // @[decode.scala 509:28 573:39]
  wire [63:0] _GEN_11060 = 12'h305 == csrAddrReg ? mscratch : _GEN_11047; // @[decode.scala 510:28 573:39]
  wire [63:0] _GEN_11061 = 12'h305 == csrAddrReg ? mepc : _GEN_11048; // @[decode.scala 511:28 573:39]
  wire [63:0] _GEN_11062 = 12'h305 == csrAddrReg ? mcause : _GEN_11049; // @[decode.scala 512:28 573:39]
  wire [63:0] _GEN_11063 = 12'h305 == csrAddrReg ? mtval : _GEN_11050; // @[decode.scala 513:28 573:39]
  wire [63:0] _GEN_11064 = 12'h305 == csrAddrReg ? mip : _GEN_11051; // @[decode.scala 514:28 573:39]
  wire [63:0] _GEN_11065 = 12'h305 == csrAddrReg ? pmpcfg0 : _GEN_11052; // @[decode.scala 515:28 573:39]
  wire [63:0] _GEN_11066 = 12'h305 == csrAddrReg ? pmpaddr0 : _GEN_11053; // @[decode.scala 516:28 573:39]
  wire [63:0] _GEN_11067 = 12'h305 == csrAddrReg ? mvendorid : _GEN_11054; // @[decode.scala 517:28 573:39]
  wire [63:0] _GEN_11068 = 12'h305 == csrAddrReg ? marchid : _GEN_11055; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_11069 = 12'h305 == csrAddrReg ? mimpid : _GEN_11056; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_11070 = 12'h305 == csrAddrReg ? mhartid : _GEN_11057; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_11071 = 12'h304 == csrAddrReg ? csrWriteData : mie; // @[decode.scala 507:28 573:39 584:37]
  wire [63:0] _GEN_11072 = 12'h304 == csrAddrReg ? mtvec : _GEN_11058; // @[decode.scala 508:28 573:39]
  wire [63:0] _GEN_11073 = 12'h304 == csrAddrReg ? mcounteren : _GEN_11059; // @[decode.scala 509:28 573:39]
  wire [63:0] _GEN_11074 = 12'h304 == csrAddrReg ? mscratch : _GEN_11060; // @[decode.scala 510:28 573:39]
  wire [63:0] _GEN_11075 = 12'h304 == csrAddrReg ? mepc : _GEN_11061; // @[decode.scala 511:28 573:39]
  wire [63:0] _GEN_11076 = 12'h304 == csrAddrReg ? mcause : _GEN_11062; // @[decode.scala 512:28 573:39]
  wire [63:0] _GEN_11077 = 12'h304 == csrAddrReg ? mtval : _GEN_11063; // @[decode.scala 513:28 573:39]
  wire [63:0] _GEN_11078 = 12'h304 == csrAddrReg ? mip : _GEN_11064; // @[decode.scala 514:28 573:39]
  wire [63:0] _GEN_11079 = 12'h304 == csrAddrReg ? pmpcfg0 : _GEN_11065; // @[decode.scala 515:28 573:39]
  wire [63:0] _GEN_11080 = 12'h304 == csrAddrReg ? pmpaddr0 : _GEN_11066; // @[decode.scala 516:28 573:39]
  wire [63:0] _GEN_11081 = 12'h304 == csrAddrReg ? mvendorid : _GEN_11067; // @[decode.scala 517:28 573:39]
  wire [63:0] _GEN_11082 = 12'h304 == csrAddrReg ? marchid : _GEN_11068; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_11083 = 12'h304 == csrAddrReg ? mimpid : _GEN_11069; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_11084 = 12'h304 == csrAddrReg ? mhartid : _GEN_11070; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_11085 = 12'h303 == csrAddrReg ? csrWriteData : mideleg; // @[decode.scala 506:28 573:39 583:37]
  wire [63:0] _GEN_11086 = 12'h303 == csrAddrReg ? mie : _GEN_11071; // @[decode.scala 507:28 573:39]
  wire [63:0] _GEN_11087 = 12'h303 == csrAddrReg ? mtvec : _GEN_11072; // @[decode.scala 508:28 573:39]
  wire [63:0] _GEN_11088 = 12'h303 == csrAddrReg ? mcounteren : _GEN_11073; // @[decode.scala 509:28 573:39]
  wire [63:0] _GEN_11089 = 12'h303 == csrAddrReg ? mscratch : _GEN_11074; // @[decode.scala 510:28 573:39]
  wire [63:0] _GEN_11090 = 12'h303 == csrAddrReg ? mepc : _GEN_11075; // @[decode.scala 511:28 573:39]
  wire [63:0] _GEN_11091 = 12'h303 == csrAddrReg ? mcause : _GEN_11076; // @[decode.scala 512:28 573:39]
  wire [63:0] _GEN_11092 = 12'h303 == csrAddrReg ? mtval : _GEN_11077; // @[decode.scala 513:28 573:39]
  wire [63:0] _GEN_11093 = 12'h303 == csrAddrReg ? mip : _GEN_11078; // @[decode.scala 514:28 573:39]
  wire [63:0] _GEN_11094 = 12'h303 == csrAddrReg ? pmpcfg0 : _GEN_11079; // @[decode.scala 515:28 573:39]
  wire [63:0] _GEN_11095 = 12'h303 == csrAddrReg ? pmpaddr0 : _GEN_11080; // @[decode.scala 516:28 573:39]
  wire [63:0] _GEN_11096 = 12'h303 == csrAddrReg ? mvendorid : _GEN_11081; // @[decode.scala 517:28 573:39]
  wire [63:0] _GEN_11097 = 12'h303 == csrAddrReg ? marchid : _GEN_11082; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_11098 = 12'h303 == csrAddrReg ? mimpid : _GEN_11083; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_11099 = 12'h303 == csrAddrReg ? mhartid : _GEN_11084; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_11100 = 12'h302 == csrAddrReg ? csrWriteData : medeleg; // @[decode.scala 505:28 573:39 582:37]
  wire [63:0] _GEN_11101 = 12'h302 == csrAddrReg ? mideleg : _GEN_11085; // @[decode.scala 506:28 573:39]
  wire [63:0] _GEN_11102 = 12'h302 == csrAddrReg ? mie : _GEN_11086; // @[decode.scala 507:28 573:39]
  wire [63:0] _GEN_11103 = 12'h302 == csrAddrReg ? mtvec : _GEN_11087; // @[decode.scala 508:28 573:39]
  wire [63:0] _GEN_11104 = 12'h302 == csrAddrReg ? mcounteren : _GEN_11088; // @[decode.scala 509:28 573:39]
  wire [63:0] _GEN_11105 = 12'h302 == csrAddrReg ? mscratch : _GEN_11089; // @[decode.scala 510:28 573:39]
  wire [63:0] _GEN_11106 = 12'h302 == csrAddrReg ? mepc : _GEN_11090; // @[decode.scala 511:28 573:39]
  wire [63:0] _GEN_11107 = 12'h302 == csrAddrReg ? mcause : _GEN_11091; // @[decode.scala 512:28 573:39]
  wire [63:0] _GEN_11108 = 12'h302 == csrAddrReg ? mtval : _GEN_11092; // @[decode.scala 513:28 573:39]
  wire [63:0] _GEN_11109 = 12'h302 == csrAddrReg ? mip : _GEN_11093; // @[decode.scala 514:28 573:39]
  wire [63:0] _GEN_11110 = 12'h302 == csrAddrReg ? pmpcfg0 : _GEN_11094; // @[decode.scala 515:28 573:39]
  wire [63:0] _GEN_11111 = 12'h302 == csrAddrReg ? pmpaddr0 : _GEN_11095; // @[decode.scala 516:28 573:39]
  wire [63:0] _GEN_11112 = 12'h302 == csrAddrReg ? mvendorid : _GEN_11096; // @[decode.scala 517:28 573:39]
  wire [63:0] _GEN_11113 = 12'h302 == csrAddrReg ? marchid : _GEN_11097; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_11114 = 12'h302 == csrAddrReg ? mimpid : _GEN_11098; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_11115 = 12'h302 == csrAddrReg ? mhartid : _GEN_11099; // @[decode.scala 520:28 573:39]
  wire [126:0] _GEN_11116 = 12'h301 == csrAddrReg ? {{63'd0}, csrWriteData} : 127'h8000000000101101; // @[decode.scala 573:39 581:37 523:8]
  wire [63:0] _GEN_11117 = 12'h301 == csrAddrReg ? medeleg : _GEN_11100; // @[decode.scala 505:28 573:39]
  wire [63:0] _GEN_11118 = 12'h301 == csrAddrReg ? mideleg : _GEN_11101; // @[decode.scala 506:28 573:39]
  wire [63:0] _GEN_11119 = 12'h301 == csrAddrReg ? mie : _GEN_11102; // @[decode.scala 507:28 573:39]
  wire [63:0] _GEN_11120 = 12'h301 == csrAddrReg ? mtvec : _GEN_11103; // @[decode.scala 508:28 573:39]
  wire [63:0] _GEN_11121 = 12'h301 == csrAddrReg ? mcounteren : _GEN_11104; // @[decode.scala 509:28 573:39]
  wire [63:0] _GEN_11122 = 12'h301 == csrAddrReg ? mscratch : _GEN_11105; // @[decode.scala 510:28 573:39]
  wire [63:0] _GEN_11123 = 12'h301 == csrAddrReg ? mepc : _GEN_11106; // @[decode.scala 511:28 573:39]
  wire [63:0] _GEN_11124 = 12'h301 == csrAddrReg ? mcause : _GEN_11107; // @[decode.scala 512:28 573:39]
  wire [63:0] _GEN_11125 = 12'h301 == csrAddrReg ? mtval : _GEN_11108; // @[decode.scala 513:28 573:39]
  wire [63:0] _GEN_11126 = 12'h301 == csrAddrReg ? mip : _GEN_11109; // @[decode.scala 514:28 573:39]
  wire [63:0] _GEN_11127 = 12'h301 == csrAddrReg ? pmpcfg0 : _GEN_11110; // @[decode.scala 515:28 573:39]
  wire [63:0] _GEN_11128 = 12'h301 == csrAddrReg ? pmpaddr0 : _GEN_11111; // @[decode.scala 516:28 573:39]
  wire [63:0] _GEN_11129 = 12'h301 == csrAddrReg ? mvendorid : _GEN_11112; // @[decode.scala 517:28 573:39]
  wire [63:0] _GEN_11130 = 12'h301 == csrAddrReg ? marchid : _GEN_11113; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_11131 = 12'h301 == csrAddrReg ? mimpid : _GEN_11114; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_11132 = 12'h301 == csrAddrReg ? mhartid : _GEN_11115; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_11133 = 12'h300 == csrAddrReg ? csrWriteData : _mstatus_T_1; // @[decode.scala 522:11 573:39 580:37]
  wire [126:0] _GEN_11134 = 12'h300 == csrAddrReg ? 127'h8000000000101101 : _GEN_11116; // @[decode.scala 573:39 523:8]
  wire [63:0] _GEN_11135 = 12'h300 == csrAddrReg ? medeleg : _GEN_11117; // @[decode.scala 505:28 573:39]
  wire [63:0] _GEN_11136 = 12'h300 == csrAddrReg ? mideleg : _GEN_11118; // @[decode.scala 506:28 573:39]
  wire [63:0] _GEN_11137 = 12'h300 == csrAddrReg ? mie : _GEN_11119; // @[decode.scala 507:28 573:39]
  wire [63:0] _GEN_11138 = 12'h300 == csrAddrReg ? mtvec : _GEN_11120; // @[decode.scala 508:28 573:39]
  wire [63:0] _GEN_11139 = 12'h300 == csrAddrReg ? mcounteren : _GEN_11121; // @[decode.scala 509:28 573:39]
  wire [63:0] _GEN_11140 = 12'h300 == csrAddrReg ? mscratch : _GEN_11122; // @[decode.scala 510:28 573:39]
  wire [63:0] _GEN_11141 = 12'h300 == csrAddrReg ? mepc : _GEN_11123; // @[decode.scala 511:28 573:39]
  wire [63:0] _GEN_11142 = 12'h300 == csrAddrReg ? mcause : _GEN_11124; // @[decode.scala 512:28 573:39]
  wire [63:0] _GEN_11143 = 12'h300 == csrAddrReg ? mtval : _GEN_11125; // @[decode.scala 513:28 573:39]
  wire [63:0] _GEN_11144 = 12'h300 == csrAddrReg ? mip : _GEN_11126; // @[decode.scala 514:28 573:39]
  wire [63:0] _GEN_11145 = 12'h300 == csrAddrReg ? pmpcfg0 : _GEN_11127; // @[decode.scala 515:28 573:39]
  wire [63:0] _GEN_11146 = 12'h300 == csrAddrReg ? pmpaddr0 : _GEN_11128; // @[decode.scala 516:28 573:39]
  wire [63:0] _GEN_11147 = 12'h300 == csrAddrReg ? mvendorid : _GEN_11129; // @[decode.scala 517:28 573:39]
  wire [63:0] _GEN_11148 = 12'h300 == csrAddrReg ? marchid : _GEN_11130; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_11149 = 12'h300 == csrAddrReg ? mimpid : _GEN_11131; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_11150 = 12'h300 == csrAddrReg ? mhartid : _GEN_11132; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_11151 = 12'h180 == csrAddrReg ? csrWriteData : satp; // @[decode.scala 502:28 573:39 579:37]
  wire [63:0] _GEN_11152 = 12'h180 == csrAddrReg ? _mstatus_T_1 : _GEN_11133; // @[decode.scala 522:11 573:39]
  wire [126:0] _GEN_11153 = 12'h180 == csrAddrReg ? 127'h8000000000101101 : _GEN_11134; // @[decode.scala 573:39 523:8]
  wire [63:0] _GEN_11154 = 12'h180 == csrAddrReg ? medeleg : _GEN_11135; // @[decode.scala 505:28 573:39]
  wire [63:0] _GEN_11155 = 12'h180 == csrAddrReg ? mideleg : _GEN_11136; // @[decode.scala 506:28 573:39]
  wire [63:0] _GEN_11156 = 12'h180 == csrAddrReg ? mie : _GEN_11137; // @[decode.scala 507:28 573:39]
  wire [63:0] _GEN_11157 = 12'h180 == csrAddrReg ? mtvec : _GEN_11138; // @[decode.scala 508:28 573:39]
  wire [63:0] _GEN_11158 = 12'h180 == csrAddrReg ? mcounteren : _GEN_11139; // @[decode.scala 509:28 573:39]
  wire [63:0] _GEN_11159 = 12'h180 == csrAddrReg ? mscratch : _GEN_11140; // @[decode.scala 510:28 573:39]
  wire [63:0] _GEN_11160 = 12'h180 == csrAddrReg ? mepc : _GEN_11141; // @[decode.scala 511:28 573:39]
  wire [63:0] _GEN_11161 = 12'h180 == csrAddrReg ? mcause : _GEN_11142; // @[decode.scala 512:28 573:39]
  wire [63:0] _GEN_11162 = 12'h180 == csrAddrReg ? mtval : _GEN_11143; // @[decode.scala 513:28 573:39]
  wire [63:0] _GEN_11163 = 12'h180 == csrAddrReg ? mip : _GEN_11144; // @[decode.scala 514:28 573:39]
  wire [63:0] _GEN_11164 = 12'h180 == csrAddrReg ? pmpcfg0 : _GEN_11145; // @[decode.scala 515:28 573:39]
  wire [63:0] _GEN_11165 = 12'h180 == csrAddrReg ? pmpaddr0 : _GEN_11146; // @[decode.scala 516:28 573:39]
  wire [63:0] _GEN_11166 = 12'h180 == csrAddrReg ? mvendorid : _GEN_11147; // @[decode.scala 517:28 573:39]
  wire [63:0] _GEN_11167 = 12'h180 == csrAddrReg ? marchid : _GEN_11148; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_11168 = 12'h180 == csrAddrReg ? mimpid : _GEN_11149; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_11169 = 12'h180 == csrAddrReg ? mhartid : _GEN_11150; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_11170 = 12'h106 == csrAddrReg ? csrWriteData : scounteren; // @[decode.scala 501:28 573:39 578:37]
  wire [63:0] _GEN_11171 = 12'h106 == csrAddrReg ? satp : _GEN_11151; // @[decode.scala 502:28 573:39]
  wire [63:0] _GEN_11172 = 12'h106 == csrAddrReg ? _mstatus_T_1 : _GEN_11152; // @[decode.scala 522:11 573:39]
  wire [126:0] _GEN_11173 = 12'h106 == csrAddrReg ? 127'h8000000000101101 : _GEN_11153; // @[decode.scala 573:39 523:8]
  wire [63:0] _GEN_11174 = 12'h106 == csrAddrReg ? medeleg : _GEN_11154; // @[decode.scala 505:28 573:39]
  wire [63:0] _GEN_11175 = 12'h106 == csrAddrReg ? mideleg : _GEN_11155; // @[decode.scala 506:28 573:39]
  wire [63:0] _GEN_11176 = 12'h106 == csrAddrReg ? mie : _GEN_11156; // @[decode.scala 507:28 573:39]
  wire [63:0] _GEN_11177 = 12'h106 == csrAddrReg ? mtvec : _GEN_11157; // @[decode.scala 508:28 573:39]
  wire [63:0] _GEN_11178 = 12'h106 == csrAddrReg ? mcounteren : _GEN_11158; // @[decode.scala 509:28 573:39]
  wire [63:0] _GEN_11179 = 12'h106 == csrAddrReg ? mscratch : _GEN_11159; // @[decode.scala 510:28 573:39]
  wire [63:0] _GEN_11180 = 12'h106 == csrAddrReg ? mepc : _GEN_11160; // @[decode.scala 511:28 573:39]
  wire [63:0] _GEN_11181 = 12'h106 == csrAddrReg ? mcause : _GEN_11161; // @[decode.scala 512:28 573:39]
  wire [63:0] _GEN_11182 = 12'h106 == csrAddrReg ? mtval : _GEN_11162; // @[decode.scala 513:28 573:39]
  wire [63:0] _GEN_11183 = 12'h106 == csrAddrReg ? mip : _GEN_11163; // @[decode.scala 514:28 573:39]
  wire [63:0] _GEN_11184 = 12'h106 == csrAddrReg ? pmpcfg0 : _GEN_11164; // @[decode.scala 515:28 573:39]
  wire [63:0] _GEN_11185 = 12'h106 == csrAddrReg ? pmpaddr0 : _GEN_11165; // @[decode.scala 516:28 573:39]
  wire [63:0] _GEN_11186 = 12'h106 == csrAddrReg ? mvendorid : _GEN_11166; // @[decode.scala 517:28 573:39]
  wire [63:0] _GEN_11187 = 12'h106 == csrAddrReg ? marchid : _GEN_11167; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_11188 = 12'h106 == csrAddrReg ? mimpid : _GEN_11168; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_11189 = 12'h106 == csrAddrReg ? mhartid : _GEN_11169; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_11190 = 12'h42 == csrAddrReg ? csrWriteData : ucause; // @[decode.scala 500:28 573:39 577:37]
  wire [63:0] _GEN_11191 = 12'h42 == csrAddrReg ? scounteren : _GEN_11170; // @[decode.scala 501:28 573:39]
  wire [63:0] _GEN_11192 = 12'h42 == csrAddrReg ? satp : _GEN_11171; // @[decode.scala 502:28 573:39]
  wire [63:0] _GEN_11193 = 12'h42 == csrAddrReg ? _mstatus_T_1 : _GEN_11172; // @[decode.scala 522:11 573:39]
  wire [126:0] _GEN_11194 = 12'h42 == csrAddrReg ? 127'h8000000000101101 : _GEN_11173; // @[decode.scala 573:39 523:8]
  wire [63:0] _GEN_11195 = 12'h42 == csrAddrReg ? medeleg : _GEN_11174; // @[decode.scala 505:28 573:39]
  wire [63:0] _GEN_11196 = 12'h42 == csrAddrReg ? mideleg : _GEN_11175; // @[decode.scala 506:28 573:39]
  wire [63:0] _GEN_11197 = 12'h42 == csrAddrReg ? mie : _GEN_11176; // @[decode.scala 507:28 573:39]
  wire [63:0] _GEN_11198 = 12'h42 == csrAddrReg ? mtvec : _GEN_11177; // @[decode.scala 508:28 573:39]
  wire [63:0] _GEN_11199 = 12'h42 == csrAddrReg ? mcounteren : _GEN_11178; // @[decode.scala 509:28 573:39]
  wire [63:0] _GEN_11200 = 12'h42 == csrAddrReg ? mscratch : _GEN_11179; // @[decode.scala 510:28 573:39]
  wire [63:0] _GEN_11201 = 12'h42 == csrAddrReg ? mepc : _GEN_11180; // @[decode.scala 511:28 573:39]
  wire [63:0] _GEN_11202 = 12'h42 == csrAddrReg ? mcause : _GEN_11181; // @[decode.scala 512:28 573:39]
  wire [63:0] _GEN_11203 = 12'h42 == csrAddrReg ? mtval : _GEN_11182; // @[decode.scala 513:28 573:39]
  wire [63:0] _GEN_11204 = 12'h42 == csrAddrReg ? mip : _GEN_11183; // @[decode.scala 514:28 573:39]
  wire [63:0] _GEN_11205 = 12'h42 == csrAddrReg ? pmpcfg0 : _GEN_11184; // @[decode.scala 515:28 573:39]
  wire [63:0] _GEN_11206 = 12'h42 == csrAddrReg ? pmpaddr0 : _GEN_11185; // @[decode.scala 516:28 573:39]
  wire [63:0] _GEN_11207 = 12'h42 == csrAddrReg ? mvendorid : _GEN_11186; // @[decode.scala 517:28 573:39]
  wire [63:0] _GEN_11208 = 12'h42 == csrAddrReg ? marchid : _GEN_11187; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_11209 = 12'h42 == csrAddrReg ? mimpid : _GEN_11188; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_11210 = 12'h42 == csrAddrReg ? mhartid : _GEN_11189; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_11211 = 12'h41 == csrAddrReg ? csrWriteData : uepc; // @[decode.scala 499:28 573:39 576:37]
  wire [63:0] _GEN_11212 = 12'h41 == csrAddrReg ? ucause : _GEN_11190; // @[decode.scala 500:28 573:39]
  wire [63:0] _GEN_11213 = 12'h41 == csrAddrReg ? scounteren : _GEN_11191; // @[decode.scala 501:28 573:39]
  wire [63:0] _GEN_11214 = 12'h41 == csrAddrReg ? satp : _GEN_11192; // @[decode.scala 502:28 573:39]
  wire [63:0] _GEN_11215 = 12'h41 == csrAddrReg ? _mstatus_T_1 : _GEN_11193; // @[decode.scala 522:11 573:39]
  wire [126:0] _GEN_11216 = 12'h41 == csrAddrReg ? 127'h8000000000101101 : _GEN_11194; // @[decode.scala 573:39 523:8]
  wire [63:0] _GEN_11217 = 12'h41 == csrAddrReg ? medeleg : _GEN_11195; // @[decode.scala 505:28 573:39]
  wire [63:0] _GEN_11218 = 12'h41 == csrAddrReg ? mideleg : _GEN_11196; // @[decode.scala 506:28 573:39]
  wire [63:0] _GEN_11219 = 12'h41 == csrAddrReg ? mie : _GEN_11197; // @[decode.scala 507:28 573:39]
  wire [63:0] _GEN_11220 = 12'h41 == csrAddrReg ? mtvec : _GEN_11198; // @[decode.scala 508:28 573:39]
  wire [63:0] _GEN_11221 = 12'h41 == csrAddrReg ? mcounteren : _GEN_11199; // @[decode.scala 509:28 573:39]
  wire [63:0] _GEN_11222 = 12'h41 == csrAddrReg ? mscratch : _GEN_11200; // @[decode.scala 510:28 573:39]
  wire [63:0] _GEN_11223 = 12'h41 == csrAddrReg ? mepc : _GEN_11201; // @[decode.scala 511:28 573:39]
  wire [63:0] _GEN_11224 = 12'h41 == csrAddrReg ? mcause : _GEN_11202; // @[decode.scala 512:28 573:39]
  wire [63:0] _GEN_11225 = 12'h41 == csrAddrReg ? mtval : _GEN_11203; // @[decode.scala 513:28 573:39]
  wire [63:0] _GEN_11226 = 12'h41 == csrAddrReg ? mip : _GEN_11204; // @[decode.scala 514:28 573:39]
  wire [63:0] _GEN_11227 = 12'h41 == csrAddrReg ? pmpcfg0 : _GEN_11205; // @[decode.scala 515:28 573:39]
  wire [63:0] _GEN_11228 = 12'h41 == csrAddrReg ? pmpaddr0 : _GEN_11206; // @[decode.scala 516:28 573:39]
  wire [63:0] _GEN_11229 = 12'h41 == csrAddrReg ? mvendorid : _GEN_11207; // @[decode.scala 517:28 573:39]
  wire [63:0] _GEN_11230 = 12'h41 == csrAddrReg ? marchid : _GEN_11208; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_11231 = 12'h41 == csrAddrReg ? mimpid : _GEN_11209; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_11232 = 12'h41 == csrAddrReg ? mhartid : _GEN_11210; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_11233 = 12'h5 == csrAddrReg ? csrWriteData : utvec; // @[decode.scala 498:28 573:39 575:37]
  wire [63:0] _GEN_11234 = 12'h5 == csrAddrReg ? uepc : _GEN_11211; // @[decode.scala 499:28 573:39]
  wire [63:0] _GEN_11235 = 12'h5 == csrAddrReg ? ucause : _GEN_11212; // @[decode.scala 500:28 573:39]
  wire [63:0] _GEN_11236 = 12'h5 == csrAddrReg ? scounteren : _GEN_11213; // @[decode.scala 501:28 573:39]
  wire [63:0] _GEN_11237 = 12'h5 == csrAddrReg ? satp : _GEN_11214; // @[decode.scala 502:28 573:39]
  wire [63:0] _GEN_11238 = 12'h5 == csrAddrReg ? _mstatus_T_1 : _GEN_11215; // @[decode.scala 522:11 573:39]
  wire [126:0] _GEN_11239 = 12'h5 == csrAddrReg ? 127'h8000000000101101 : _GEN_11216; // @[decode.scala 573:39 523:8]
  wire [63:0] _GEN_11240 = 12'h5 == csrAddrReg ? medeleg : _GEN_11217; // @[decode.scala 505:28 573:39]
  wire [63:0] _GEN_11241 = 12'h5 == csrAddrReg ? mideleg : _GEN_11218; // @[decode.scala 506:28 573:39]
  wire [63:0] _GEN_11242 = 12'h5 == csrAddrReg ? mie : _GEN_11219; // @[decode.scala 507:28 573:39]
  wire [63:0] _GEN_11243 = 12'h5 == csrAddrReg ? mtvec : _GEN_11220; // @[decode.scala 508:28 573:39]
  wire [63:0] _GEN_11244 = 12'h5 == csrAddrReg ? mcounteren : _GEN_11221; // @[decode.scala 509:28 573:39]
  wire [63:0] _GEN_11245 = 12'h5 == csrAddrReg ? mscratch : _GEN_11222; // @[decode.scala 510:28 573:39]
  wire [63:0] _GEN_11246 = 12'h5 == csrAddrReg ? mepc : _GEN_11223; // @[decode.scala 511:28 573:39]
  wire [63:0] _GEN_11247 = 12'h5 == csrAddrReg ? mcause : _GEN_11224; // @[decode.scala 512:28 573:39]
  wire [63:0] _GEN_11248 = 12'h5 == csrAddrReg ? mtval : _GEN_11225; // @[decode.scala 513:28 573:39]
  wire [63:0] _GEN_11249 = 12'h5 == csrAddrReg ? mip : _GEN_11226; // @[decode.scala 514:28 573:39]
  wire [63:0] _GEN_11250 = 12'h5 == csrAddrReg ? pmpcfg0 : _GEN_11227; // @[decode.scala 515:28 573:39]
  wire [63:0] _GEN_11251 = 12'h5 == csrAddrReg ? pmpaddr0 : _GEN_11228; // @[decode.scala 516:28 573:39]
  wire [63:0] _GEN_11252 = 12'h5 == csrAddrReg ? mvendorid : _GEN_11229; // @[decode.scala 517:28 573:39]
  wire [63:0] _GEN_11253 = 12'h5 == csrAddrReg ? marchid : _GEN_11230; // @[decode.scala 518:28 573:39]
  wire [63:0] _GEN_11254 = 12'h5 == csrAddrReg ? mimpid : _GEN_11231; // @[decode.scala 519:28 573:39]
  wire [63:0] _GEN_11255 = 12'h5 == csrAddrReg ? mhartid : _GEN_11232; // @[decode.scala 520:28 573:39]
  wire [63:0] _GEN_11262 = 12'h0 == csrAddrReg ? _mstatus_T_1 : _GEN_11238; // @[decode.scala 522:11 573:39]
  wire [126:0] _GEN_11263 = 12'h0 == csrAddrReg ? 127'h8000000000101101 : _GEN_11239; // @[decode.scala 573:39 523:8]
  wire [63:0] _GEN_11270 = 12'h0 == csrAddrReg ? mepc : _GEN_11246; // @[decode.scala 511:28 573:39]
  wire [63:0] _GEN_11271 = 12'h0 == csrAddrReg ? mcause : _GEN_11247; // @[decode.scala 512:28 573:39]
  wire [63:0] _ustatus_T = ustatus | csrWriteData; // @[decode.scala 602:49]
  wire [63:0] _utvec_T = utvec | csrWriteData; // @[decode.scala 603:47]
  wire [63:0] _uepc_T = uepc | csrWriteData; // @[decode.scala 604:46]
  wire [63:0] _ucause_T = ucause | csrWriteData; // @[decode.scala 605:48]
  wire [63:0] _scounteren_T = scounteren | csrWriteData; // @[decode.scala 606:52]
  wire [63:0] _satp_T = satp | csrWriteData; // @[decode.scala 607:46]
  wire [63:0] _mstatus_T_2 = mstatus | csrWriteData; // @[decode.scala 608:49]
  wire [63:0] _misa_T_2 = misa | csrWriteData; // @[decode.scala 609:46]
  wire [63:0] _medeleg_T = medeleg | csrWriteData; // @[decode.scala 610:49]
  wire [63:0] _mideleg_T = mideleg | csrWriteData; // @[decode.scala 611:49]
  wire [63:0] _mie_T = mie | csrWriteData; // @[decode.scala 612:46]
  wire [63:0] _mtvec_T = mtvec | csrWriteData; // @[decode.scala 613:47]
  wire [63:0] _mcounteren_T = mcounteren | csrWriteData; // @[decode.scala 614:52]
  wire [63:0] _mscratch_T = mscratch | csrWriteData; // @[decode.scala 615:50]
  wire [63:0] _mepc_T = mepc | csrWriteData; // @[decode.scala 616:46]
  wire [63:0] _mcause_T = mcause | csrWriteData; // @[decode.scala 617:48]
  wire [63:0] _mtval_T = mtval | csrWriteData; // @[decode.scala 618:47]
  wire [63:0] _mip_T = mip | csrWriteData; // @[decode.scala 619:45]
  wire [63:0] _pmpcfg0_T = pmpcfg0 | csrWriteData; // @[decode.scala 620:49]
  wire [63:0] _pmpaddr0_T = pmpaddr0 | csrWriteData; // @[decode.scala 621:50]
  wire [63:0] _mvendorid_T = mvendorid | csrWriteData; // @[decode.scala 622:51]
  wire [63:0] _marchid_T = marchid | csrWriteData; // @[decode.scala 623:49]
  wire [63:0] _mimpid_T = mimpid | csrWriteData; // @[decode.scala 624:48]
  wire [63:0] _mhartid_T = mhartid | csrWriteData; // @[decode.scala 625:49]
  wire [63:0] _GEN_11280 = _T_289 ? _mhartid_T : mhartid; // @[decode.scala 520:28 601:39 625:38]
  wire [63:0] _GEN_11281 = _T_288 ? _mimpid_T : mimpid; // @[decode.scala 519:28 601:39 624:38]
  wire [63:0] _GEN_11282 = _T_288 ? mhartid : _GEN_11280; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11283 = _T_287 ? _marchid_T : marchid; // @[decode.scala 518:28 601:39 623:38]
  wire [63:0] _GEN_11284 = _T_287 ? mimpid : _GEN_11281; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11285 = _T_287 ? mhartid : _GEN_11282; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11286 = _T_286 ? _mvendorid_T : mvendorid; // @[decode.scala 517:28 601:39 622:38]
  wire [63:0] _GEN_11287 = _T_286 ? marchid : _GEN_11283; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11288 = _T_286 ? mimpid : _GEN_11284; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11289 = _T_286 ? mhartid : _GEN_11285; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11290 = _T_285 ? _pmpaddr0_T : pmpaddr0; // @[decode.scala 516:28 601:39 621:38]
  wire [63:0] _GEN_11291 = _T_285 ? mvendorid : _GEN_11286; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11292 = _T_285 ? marchid : _GEN_11287; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11293 = _T_285 ? mimpid : _GEN_11288; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11294 = _T_285 ? mhartid : _GEN_11289; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11295 = _T_284 ? _pmpcfg0_T : pmpcfg0; // @[decode.scala 515:28 601:39 620:38]
  wire [63:0] _GEN_11296 = _T_284 ? pmpaddr0 : _GEN_11290; // @[decode.scala 516:28 601:39]
  wire [63:0] _GEN_11297 = _T_284 ? mvendorid : _GEN_11291; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11298 = _T_284 ? marchid : _GEN_11292; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11299 = _T_284 ? mimpid : _GEN_11293; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11300 = _T_284 ? mhartid : _GEN_11294; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11301 = _T_283 ? _mip_T : mip; // @[decode.scala 514:28 601:39 619:38]
  wire [63:0] _GEN_11302 = _T_283 ? pmpcfg0 : _GEN_11295; // @[decode.scala 515:28 601:39]
  wire [63:0] _GEN_11303 = _T_283 ? pmpaddr0 : _GEN_11296; // @[decode.scala 516:28 601:39]
  wire [63:0] _GEN_11304 = _T_283 ? mvendorid : _GEN_11297; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11305 = _T_283 ? marchid : _GEN_11298; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11306 = _T_283 ? mimpid : _GEN_11299; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11307 = _T_283 ? mhartid : _GEN_11300; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11308 = _T_282 ? _mtval_T : mtval; // @[decode.scala 513:28 601:39 618:38]
  wire [63:0] _GEN_11309 = _T_282 ? mip : _GEN_11301; // @[decode.scala 514:28 601:39]
  wire [63:0] _GEN_11310 = _T_282 ? pmpcfg0 : _GEN_11302; // @[decode.scala 515:28 601:39]
  wire [63:0] _GEN_11311 = _T_282 ? pmpaddr0 : _GEN_11303; // @[decode.scala 516:28 601:39]
  wire [63:0] _GEN_11312 = _T_282 ? mvendorid : _GEN_11304; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11313 = _T_282 ? marchid : _GEN_11305; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11314 = _T_282 ? mimpid : _GEN_11306; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11315 = _T_282 ? mhartid : _GEN_11307; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11316 = _T_281 ? _mcause_T : mcause; // @[decode.scala 512:28 601:39 617:38]
  wire [63:0] _GEN_11317 = _T_281 ? mtval : _GEN_11308; // @[decode.scala 513:28 601:39]
  wire [63:0] _GEN_11318 = _T_281 ? mip : _GEN_11309; // @[decode.scala 514:28 601:39]
  wire [63:0] _GEN_11319 = _T_281 ? pmpcfg0 : _GEN_11310; // @[decode.scala 515:28 601:39]
  wire [63:0] _GEN_11320 = _T_281 ? pmpaddr0 : _GEN_11311; // @[decode.scala 516:28 601:39]
  wire [63:0] _GEN_11321 = _T_281 ? mvendorid : _GEN_11312; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11322 = _T_281 ? marchid : _GEN_11313; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11323 = _T_281 ? mimpid : _GEN_11314; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11324 = _T_281 ? mhartid : _GEN_11315; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11325 = _T_280 ? _mepc_T : mepc; // @[decode.scala 511:28 601:39 616:38]
  wire [63:0] _GEN_11326 = _T_280 ? mcause : _GEN_11316; // @[decode.scala 512:28 601:39]
  wire [63:0] _GEN_11327 = _T_280 ? mtval : _GEN_11317; // @[decode.scala 513:28 601:39]
  wire [63:0] _GEN_11328 = _T_280 ? mip : _GEN_11318; // @[decode.scala 514:28 601:39]
  wire [63:0] _GEN_11329 = _T_280 ? pmpcfg0 : _GEN_11319; // @[decode.scala 515:28 601:39]
  wire [63:0] _GEN_11330 = _T_280 ? pmpaddr0 : _GEN_11320; // @[decode.scala 516:28 601:39]
  wire [63:0] _GEN_11331 = _T_280 ? mvendorid : _GEN_11321; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11332 = _T_280 ? marchid : _GEN_11322; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11333 = _T_280 ? mimpid : _GEN_11323; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11334 = _T_280 ? mhartid : _GEN_11324; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11335 = _T_279 ? _mscratch_T : mscratch; // @[decode.scala 510:28 601:39 615:38]
  wire [63:0] _GEN_11336 = _T_279 ? mepc : _GEN_11325; // @[decode.scala 511:28 601:39]
  wire [63:0] _GEN_11337 = _T_279 ? mcause : _GEN_11326; // @[decode.scala 512:28 601:39]
  wire [63:0] _GEN_11338 = _T_279 ? mtval : _GEN_11327; // @[decode.scala 513:28 601:39]
  wire [63:0] _GEN_11339 = _T_279 ? mip : _GEN_11328; // @[decode.scala 514:28 601:39]
  wire [63:0] _GEN_11340 = _T_279 ? pmpcfg0 : _GEN_11329; // @[decode.scala 515:28 601:39]
  wire [63:0] _GEN_11341 = _T_279 ? pmpaddr0 : _GEN_11330; // @[decode.scala 516:28 601:39]
  wire [63:0] _GEN_11342 = _T_279 ? mvendorid : _GEN_11331; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11343 = _T_279 ? marchid : _GEN_11332; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11344 = _T_279 ? mimpid : _GEN_11333; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11345 = _T_279 ? mhartid : _GEN_11334; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11346 = _T_278 ? _mcounteren_T : mcounteren; // @[decode.scala 509:28 601:39 614:38]
  wire [63:0] _GEN_11347 = _T_278 ? mscratch : _GEN_11335; // @[decode.scala 510:28 601:39]
  wire [63:0] _GEN_11348 = _T_278 ? mepc : _GEN_11336; // @[decode.scala 511:28 601:39]
  wire [63:0] _GEN_11349 = _T_278 ? mcause : _GEN_11337; // @[decode.scala 512:28 601:39]
  wire [63:0] _GEN_11350 = _T_278 ? mtval : _GEN_11338; // @[decode.scala 513:28 601:39]
  wire [63:0] _GEN_11351 = _T_278 ? mip : _GEN_11339; // @[decode.scala 514:28 601:39]
  wire [63:0] _GEN_11352 = _T_278 ? pmpcfg0 : _GEN_11340; // @[decode.scala 515:28 601:39]
  wire [63:0] _GEN_11353 = _T_278 ? pmpaddr0 : _GEN_11341; // @[decode.scala 516:28 601:39]
  wire [63:0] _GEN_11354 = _T_278 ? mvendorid : _GEN_11342; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11355 = _T_278 ? marchid : _GEN_11343; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11356 = _T_278 ? mimpid : _GEN_11344; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11357 = _T_278 ? mhartid : _GEN_11345; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11358 = _T_277 ? _mtvec_T : mtvec; // @[decode.scala 508:28 601:39 613:38]
  wire [63:0] _GEN_11359 = _T_277 ? mcounteren : _GEN_11346; // @[decode.scala 509:28 601:39]
  wire [63:0] _GEN_11360 = _T_277 ? mscratch : _GEN_11347; // @[decode.scala 510:28 601:39]
  wire [63:0] _GEN_11361 = _T_277 ? mepc : _GEN_11348; // @[decode.scala 511:28 601:39]
  wire [63:0] _GEN_11362 = _T_277 ? mcause : _GEN_11349; // @[decode.scala 512:28 601:39]
  wire [63:0] _GEN_11363 = _T_277 ? mtval : _GEN_11350; // @[decode.scala 513:28 601:39]
  wire [63:0] _GEN_11364 = _T_277 ? mip : _GEN_11351; // @[decode.scala 514:28 601:39]
  wire [63:0] _GEN_11365 = _T_277 ? pmpcfg0 : _GEN_11352; // @[decode.scala 515:28 601:39]
  wire [63:0] _GEN_11366 = _T_277 ? pmpaddr0 : _GEN_11353; // @[decode.scala 516:28 601:39]
  wire [63:0] _GEN_11367 = _T_277 ? mvendorid : _GEN_11354; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11368 = _T_277 ? marchid : _GEN_11355; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11369 = _T_277 ? mimpid : _GEN_11356; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11370 = _T_277 ? mhartid : _GEN_11357; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11371 = _T_276 ? _mie_T : mie; // @[decode.scala 507:28 601:39 612:38]
  wire [63:0] _GEN_11372 = _T_276 ? mtvec : _GEN_11358; // @[decode.scala 508:28 601:39]
  wire [63:0] _GEN_11373 = _T_276 ? mcounteren : _GEN_11359; // @[decode.scala 509:28 601:39]
  wire [63:0] _GEN_11374 = _T_276 ? mscratch : _GEN_11360; // @[decode.scala 510:28 601:39]
  wire [63:0] _GEN_11375 = _T_276 ? mepc : _GEN_11361; // @[decode.scala 511:28 601:39]
  wire [63:0] _GEN_11376 = _T_276 ? mcause : _GEN_11362; // @[decode.scala 512:28 601:39]
  wire [63:0] _GEN_11377 = _T_276 ? mtval : _GEN_11363; // @[decode.scala 513:28 601:39]
  wire [63:0] _GEN_11378 = _T_276 ? mip : _GEN_11364; // @[decode.scala 514:28 601:39]
  wire [63:0] _GEN_11379 = _T_276 ? pmpcfg0 : _GEN_11365; // @[decode.scala 515:28 601:39]
  wire [63:0] _GEN_11380 = _T_276 ? pmpaddr0 : _GEN_11366; // @[decode.scala 516:28 601:39]
  wire [63:0] _GEN_11381 = _T_276 ? mvendorid : _GEN_11367; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11382 = _T_276 ? marchid : _GEN_11368; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11383 = _T_276 ? mimpid : _GEN_11369; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11384 = _T_276 ? mhartid : _GEN_11370; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11385 = _T_275 ? _mideleg_T : mideleg; // @[decode.scala 506:28 601:39 611:38]
  wire [63:0] _GEN_11386 = _T_275 ? mie : _GEN_11371; // @[decode.scala 507:28 601:39]
  wire [63:0] _GEN_11387 = _T_275 ? mtvec : _GEN_11372; // @[decode.scala 508:28 601:39]
  wire [63:0] _GEN_11388 = _T_275 ? mcounteren : _GEN_11373; // @[decode.scala 509:28 601:39]
  wire [63:0] _GEN_11389 = _T_275 ? mscratch : _GEN_11374; // @[decode.scala 510:28 601:39]
  wire [63:0] _GEN_11390 = _T_275 ? mepc : _GEN_11375; // @[decode.scala 511:28 601:39]
  wire [63:0] _GEN_11391 = _T_275 ? mcause : _GEN_11376; // @[decode.scala 512:28 601:39]
  wire [63:0] _GEN_11392 = _T_275 ? mtval : _GEN_11377; // @[decode.scala 513:28 601:39]
  wire [63:0] _GEN_11393 = _T_275 ? mip : _GEN_11378; // @[decode.scala 514:28 601:39]
  wire [63:0] _GEN_11394 = _T_275 ? pmpcfg0 : _GEN_11379; // @[decode.scala 515:28 601:39]
  wire [63:0] _GEN_11395 = _T_275 ? pmpaddr0 : _GEN_11380; // @[decode.scala 516:28 601:39]
  wire [63:0] _GEN_11396 = _T_275 ? mvendorid : _GEN_11381; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11397 = _T_275 ? marchid : _GEN_11382; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11398 = _T_275 ? mimpid : _GEN_11383; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11399 = _T_275 ? mhartid : _GEN_11384; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11400 = _T_274 ? _medeleg_T : medeleg; // @[decode.scala 505:28 601:39 610:38]
  wire [63:0] _GEN_11401 = _T_274 ? mideleg : _GEN_11385; // @[decode.scala 506:28 601:39]
  wire [63:0] _GEN_11402 = _T_274 ? mie : _GEN_11386; // @[decode.scala 507:28 601:39]
  wire [63:0] _GEN_11403 = _T_274 ? mtvec : _GEN_11387; // @[decode.scala 508:28 601:39]
  wire [63:0] _GEN_11404 = _T_274 ? mcounteren : _GEN_11388; // @[decode.scala 509:28 601:39]
  wire [63:0] _GEN_11405 = _T_274 ? mscratch : _GEN_11389; // @[decode.scala 510:28 601:39]
  wire [63:0] _GEN_11406 = _T_274 ? mepc : _GEN_11390; // @[decode.scala 511:28 601:39]
  wire [63:0] _GEN_11407 = _T_274 ? mcause : _GEN_11391; // @[decode.scala 512:28 601:39]
  wire [63:0] _GEN_11408 = _T_274 ? mtval : _GEN_11392; // @[decode.scala 513:28 601:39]
  wire [63:0] _GEN_11409 = _T_274 ? mip : _GEN_11393; // @[decode.scala 514:28 601:39]
  wire [63:0] _GEN_11410 = _T_274 ? pmpcfg0 : _GEN_11394; // @[decode.scala 515:28 601:39]
  wire [63:0] _GEN_11411 = _T_274 ? pmpaddr0 : _GEN_11395; // @[decode.scala 516:28 601:39]
  wire [63:0] _GEN_11412 = _T_274 ? mvendorid : _GEN_11396; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11413 = _T_274 ? marchid : _GEN_11397; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11414 = _T_274 ? mimpid : _GEN_11398; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11415 = _T_274 ? mhartid : _GEN_11399; // @[decode.scala 520:28 601:39]
  wire [126:0] _GEN_11416 = _T_273 ? {{63'd0}, _misa_T_2} : 127'h8000000000101101; // @[decode.scala 601:39 609:38 523:8]
  wire [63:0] _GEN_11417 = _T_273 ? medeleg : _GEN_11400; // @[decode.scala 505:28 601:39]
  wire [63:0] _GEN_11418 = _T_273 ? mideleg : _GEN_11401; // @[decode.scala 506:28 601:39]
  wire [63:0] _GEN_11419 = _T_273 ? mie : _GEN_11402; // @[decode.scala 507:28 601:39]
  wire [63:0] _GEN_11420 = _T_273 ? mtvec : _GEN_11403; // @[decode.scala 508:28 601:39]
  wire [63:0] _GEN_11421 = _T_273 ? mcounteren : _GEN_11404; // @[decode.scala 509:28 601:39]
  wire [63:0] _GEN_11422 = _T_273 ? mscratch : _GEN_11405; // @[decode.scala 510:28 601:39]
  wire [63:0] _GEN_11423 = _T_273 ? mepc : _GEN_11406; // @[decode.scala 511:28 601:39]
  wire [63:0] _GEN_11424 = _T_273 ? mcause : _GEN_11407; // @[decode.scala 512:28 601:39]
  wire [63:0] _GEN_11425 = _T_273 ? mtval : _GEN_11408; // @[decode.scala 513:28 601:39]
  wire [63:0] _GEN_11426 = _T_273 ? mip : _GEN_11409; // @[decode.scala 514:28 601:39]
  wire [63:0] _GEN_11427 = _T_273 ? pmpcfg0 : _GEN_11410; // @[decode.scala 515:28 601:39]
  wire [63:0] _GEN_11428 = _T_273 ? pmpaddr0 : _GEN_11411; // @[decode.scala 516:28 601:39]
  wire [63:0] _GEN_11429 = _T_273 ? mvendorid : _GEN_11412; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11430 = _T_273 ? marchid : _GEN_11413; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11431 = _T_273 ? mimpid : _GEN_11414; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11432 = _T_273 ? mhartid : _GEN_11415; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11433 = _T_272 ? _mstatus_T_2 : _mstatus_T_1; // @[decode.scala 522:11 601:39 608:38]
  wire [126:0] _GEN_11434 = _T_272 ? 127'h8000000000101101 : _GEN_11416; // @[decode.scala 601:39 523:8]
  wire [63:0] _GEN_11435 = _T_272 ? medeleg : _GEN_11417; // @[decode.scala 505:28 601:39]
  wire [63:0] _GEN_11436 = _T_272 ? mideleg : _GEN_11418; // @[decode.scala 506:28 601:39]
  wire [63:0] _GEN_11437 = _T_272 ? mie : _GEN_11419; // @[decode.scala 507:28 601:39]
  wire [63:0] _GEN_11438 = _T_272 ? mtvec : _GEN_11420; // @[decode.scala 508:28 601:39]
  wire [63:0] _GEN_11439 = _T_272 ? mcounteren : _GEN_11421; // @[decode.scala 509:28 601:39]
  wire [63:0] _GEN_11440 = _T_272 ? mscratch : _GEN_11422; // @[decode.scala 510:28 601:39]
  wire [63:0] _GEN_11441 = _T_272 ? mepc : _GEN_11423; // @[decode.scala 511:28 601:39]
  wire [63:0] _GEN_11442 = _T_272 ? mcause : _GEN_11424; // @[decode.scala 512:28 601:39]
  wire [63:0] _GEN_11443 = _T_272 ? mtval : _GEN_11425; // @[decode.scala 513:28 601:39]
  wire [63:0] _GEN_11444 = _T_272 ? mip : _GEN_11426; // @[decode.scala 514:28 601:39]
  wire [63:0] _GEN_11445 = _T_272 ? pmpcfg0 : _GEN_11427; // @[decode.scala 515:28 601:39]
  wire [63:0] _GEN_11446 = _T_272 ? pmpaddr0 : _GEN_11428; // @[decode.scala 516:28 601:39]
  wire [63:0] _GEN_11447 = _T_272 ? mvendorid : _GEN_11429; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11448 = _T_272 ? marchid : _GEN_11430; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11449 = _T_272 ? mimpid : _GEN_11431; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11450 = _T_272 ? mhartid : _GEN_11432; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11451 = _T_271 ? _satp_T : satp; // @[decode.scala 502:28 601:39 607:38]
  wire [63:0] _GEN_11452 = _T_271 ? _mstatus_T_1 : _GEN_11433; // @[decode.scala 522:11 601:39]
  wire [126:0] _GEN_11453 = _T_271 ? 127'h8000000000101101 : _GEN_11434; // @[decode.scala 601:39 523:8]
  wire [63:0] _GEN_11454 = _T_271 ? medeleg : _GEN_11435; // @[decode.scala 505:28 601:39]
  wire [63:0] _GEN_11455 = _T_271 ? mideleg : _GEN_11436; // @[decode.scala 506:28 601:39]
  wire [63:0] _GEN_11456 = _T_271 ? mie : _GEN_11437; // @[decode.scala 507:28 601:39]
  wire [63:0] _GEN_11457 = _T_271 ? mtvec : _GEN_11438; // @[decode.scala 508:28 601:39]
  wire [63:0] _GEN_11458 = _T_271 ? mcounteren : _GEN_11439; // @[decode.scala 509:28 601:39]
  wire [63:0] _GEN_11459 = _T_271 ? mscratch : _GEN_11440; // @[decode.scala 510:28 601:39]
  wire [63:0] _GEN_11460 = _T_271 ? mepc : _GEN_11441; // @[decode.scala 511:28 601:39]
  wire [63:0] _GEN_11461 = _T_271 ? mcause : _GEN_11442; // @[decode.scala 512:28 601:39]
  wire [63:0] _GEN_11462 = _T_271 ? mtval : _GEN_11443; // @[decode.scala 513:28 601:39]
  wire [63:0] _GEN_11463 = _T_271 ? mip : _GEN_11444; // @[decode.scala 514:28 601:39]
  wire [63:0] _GEN_11464 = _T_271 ? pmpcfg0 : _GEN_11445; // @[decode.scala 515:28 601:39]
  wire [63:0] _GEN_11465 = _T_271 ? pmpaddr0 : _GEN_11446; // @[decode.scala 516:28 601:39]
  wire [63:0] _GEN_11466 = _T_271 ? mvendorid : _GEN_11447; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11467 = _T_271 ? marchid : _GEN_11448; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11468 = _T_271 ? mimpid : _GEN_11449; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11469 = _T_271 ? mhartid : _GEN_11450; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11470 = _T_270 ? _scounteren_T : scounteren; // @[decode.scala 501:28 601:39 606:38]
  wire [63:0] _GEN_11471 = _T_270 ? satp : _GEN_11451; // @[decode.scala 502:28 601:39]
  wire [63:0] _GEN_11472 = _T_270 ? _mstatus_T_1 : _GEN_11452; // @[decode.scala 522:11 601:39]
  wire [126:0] _GEN_11473 = _T_270 ? 127'h8000000000101101 : _GEN_11453; // @[decode.scala 601:39 523:8]
  wire [63:0] _GEN_11474 = _T_270 ? medeleg : _GEN_11454; // @[decode.scala 505:28 601:39]
  wire [63:0] _GEN_11475 = _T_270 ? mideleg : _GEN_11455; // @[decode.scala 506:28 601:39]
  wire [63:0] _GEN_11476 = _T_270 ? mie : _GEN_11456; // @[decode.scala 507:28 601:39]
  wire [63:0] _GEN_11477 = _T_270 ? mtvec : _GEN_11457; // @[decode.scala 508:28 601:39]
  wire [63:0] _GEN_11478 = _T_270 ? mcounteren : _GEN_11458; // @[decode.scala 509:28 601:39]
  wire [63:0] _GEN_11479 = _T_270 ? mscratch : _GEN_11459; // @[decode.scala 510:28 601:39]
  wire [63:0] _GEN_11480 = _T_270 ? mepc : _GEN_11460; // @[decode.scala 511:28 601:39]
  wire [63:0] _GEN_11481 = _T_270 ? mcause : _GEN_11461; // @[decode.scala 512:28 601:39]
  wire [63:0] _GEN_11482 = _T_270 ? mtval : _GEN_11462; // @[decode.scala 513:28 601:39]
  wire [63:0] _GEN_11483 = _T_270 ? mip : _GEN_11463; // @[decode.scala 514:28 601:39]
  wire [63:0] _GEN_11484 = _T_270 ? pmpcfg0 : _GEN_11464; // @[decode.scala 515:28 601:39]
  wire [63:0] _GEN_11485 = _T_270 ? pmpaddr0 : _GEN_11465; // @[decode.scala 516:28 601:39]
  wire [63:0] _GEN_11486 = _T_270 ? mvendorid : _GEN_11466; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11487 = _T_270 ? marchid : _GEN_11467; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11488 = _T_270 ? mimpid : _GEN_11468; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11489 = _T_270 ? mhartid : _GEN_11469; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11490 = _T_269 ? _ucause_T : ucause; // @[decode.scala 500:28 601:39 605:38]
  wire [63:0] _GEN_11491 = _T_269 ? scounteren : _GEN_11470; // @[decode.scala 501:28 601:39]
  wire [63:0] _GEN_11492 = _T_269 ? satp : _GEN_11471; // @[decode.scala 502:28 601:39]
  wire [63:0] _GEN_11493 = _T_269 ? _mstatus_T_1 : _GEN_11472; // @[decode.scala 522:11 601:39]
  wire [126:0] _GEN_11494 = _T_269 ? 127'h8000000000101101 : _GEN_11473; // @[decode.scala 601:39 523:8]
  wire [63:0] _GEN_11495 = _T_269 ? medeleg : _GEN_11474; // @[decode.scala 505:28 601:39]
  wire [63:0] _GEN_11496 = _T_269 ? mideleg : _GEN_11475; // @[decode.scala 506:28 601:39]
  wire [63:0] _GEN_11497 = _T_269 ? mie : _GEN_11476; // @[decode.scala 507:28 601:39]
  wire [63:0] _GEN_11498 = _T_269 ? mtvec : _GEN_11477; // @[decode.scala 508:28 601:39]
  wire [63:0] _GEN_11499 = _T_269 ? mcounteren : _GEN_11478; // @[decode.scala 509:28 601:39]
  wire [63:0] _GEN_11500 = _T_269 ? mscratch : _GEN_11479; // @[decode.scala 510:28 601:39]
  wire [63:0] _GEN_11501 = _T_269 ? mepc : _GEN_11480; // @[decode.scala 511:28 601:39]
  wire [63:0] _GEN_11502 = _T_269 ? mcause : _GEN_11481; // @[decode.scala 512:28 601:39]
  wire [63:0] _GEN_11503 = _T_269 ? mtval : _GEN_11482; // @[decode.scala 513:28 601:39]
  wire [63:0] _GEN_11504 = _T_269 ? mip : _GEN_11483; // @[decode.scala 514:28 601:39]
  wire [63:0] _GEN_11505 = _T_269 ? pmpcfg0 : _GEN_11484; // @[decode.scala 515:28 601:39]
  wire [63:0] _GEN_11506 = _T_269 ? pmpaddr0 : _GEN_11485; // @[decode.scala 516:28 601:39]
  wire [63:0] _GEN_11507 = _T_269 ? mvendorid : _GEN_11486; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11508 = _T_269 ? marchid : _GEN_11487; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11509 = _T_269 ? mimpid : _GEN_11488; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11510 = _T_269 ? mhartid : _GEN_11489; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11511 = _T_268 ? _uepc_T : uepc; // @[decode.scala 499:28 601:39 604:38]
  wire [63:0] _GEN_11512 = _T_268 ? ucause : _GEN_11490; // @[decode.scala 500:28 601:39]
  wire [63:0] _GEN_11513 = _T_268 ? scounteren : _GEN_11491; // @[decode.scala 501:28 601:39]
  wire [63:0] _GEN_11514 = _T_268 ? satp : _GEN_11492; // @[decode.scala 502:28 601:39]
  wire [63:0] _GEN_11515 = _T_268 ? _mstatus_T_1 : _GEN_11493; // @[decode.scala 522:11 601:39]
  wire [126:0] _GEN_11516 = _T_268 ? 127'h8000000000101101 : _GEN_11494; // @[decode.scala 601:39 523:8]
  wire [63:0] _GEN_11517 = _T_268 ? medeleg : _GEN_11495; // @[decode.scala 505:28 601:39]
  wire [63:0] _GEN_11518 = _T_268 ? mideleg : _GEN_11496; // @[decode.scala 506:28 601:39]
  wire [63:0] _GEN_11519 = _T_268 ? mie : _GEN_11497; // @[decode.scala 507:28 601:39]
  wire [63:0] _GEN_11520 = _T_268 ? mtvec : _GEN_11498; // @[decode.scala 508:28 601:39]
  wire [63:0] _GEN_11521 = _T_268 ? mcounteren : _GEN_11499; // @[decode.scala 509:28 601:39]
  wire [63:0] _GEN_11522 = _T_268 ? mscratch : _GEN_11500; // @[decode.scala 510:28 601:39]
  wire [63:0] _GEN_11523 = _T_268 ? mepc : _GEN_11501; // @[decode.scala 511:28 601:39]
  wire [63:0] _GEN_11524 = _T_268 ? mcause : _GEN_11502; // @[decode.scala 512:28 601:39]
  wire [63:0] _GEN_11525 = _T_268 ? mtval : _GEN_11503; // @[decode.scala 513:28 601:39]
  wire [63:0] _GEN_11526 = _T_268 ? mip : _GEN_11504; // @[decode.scala 514:28 601:39]
  wire [63:0] _GEN_11527 = _T_268 ? pmpcfg0 : _GEN_11505; // @[decode.scala 515:28 601:39]
  wire [63:0] _GEN_11528 = _T_268 ? pmpaddr0 : _GEN_11506; // @[decode.scala 516:28 601:39]
  wire [63:0] _GEN_11529 = _T_268 ? mvendorid : _GEN_11507; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11530 = _T_268 ? marchid : _GEN_11508; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11531 = _T_268 ? mimpid : _GEN_11509; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11532 = _T_268 ? mhartid : _GEN_11510; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11533 = _T_267 ? _utvec_T : utvec; // @[decode.scala 498:28 601:39 603:38]
  wire [63:0] _GEN_11534 = _T_267 ? uepc : _GEN_11511; // @[decode.scala 499:28 601:39]
  wire [63:0] _GEN_11535 = _T_267 ? ucause : _GEN_11512; // @[decode.scala 500:28 601:39]
  wire [63:0] _GEN_11536 = _T_267 ? scounteren : _GEN_11513; // @[decode.scala 501:28 601:39]
  wire [63:0] _GEN_11537 = _T_267 ? satp : _GEN_11514; // @[decode.scala 502:28 601:39]
  wire [63:0] _GEN_11538 = _T_267 ? _mstatus_T_1 : _GEN_11515; // @[decode.scala 522:11 601:39]
  wire [126:0] _GEN_11539 = _T_267 ? 127'h8000000000101101 : _GEN_11516; // @[decode.scala 601:39 523:8]
  wire [63:0] _GEN_11540 = _T_267 ? medeleg : _GEN_11517; // @[decode.scala 505:28 601:39]
  wire [63:0] _GEN_11541 = _T_267 ? mideleg : _GEN_11518; // @[decode.scala 506:28 601:39]
  wire [63:0] _GEN_11542 = _T_267 ? mie : _GEN_11519; // @[decode.scala 507:28 601:39]
  wire [63:0] _GEN_11543 = _T_267 ? mtvec : _GEN_11520; // @[decode.scala 508:28 601:39]
  wire [63:0] _GEN_11544 = _T_267 ? mcounteren : _GEN_11521; // @[decode.scala 509:28 601:39]
  wire [63:0] _GEN_11545 = _T_267 ? mscratch : _GEN_11522; // @[decode.scala 510:28 601:39]
  wire [63:0] _GEN_11546 = _T_267 ? mepc : _GEN_11523; // @[decode.scala 511:28 601:39]
  wire [63:0] _GEN_11547 = _T_267 ? mcause : _GEN_11524; // @[decode.scala 512:28 601:39]
  wire [63:0] _GEN_11548 = _T_267 ? mtval : _GEN_11525; // @[decode.scala 513:28 601:39]
  wire [63:0] _GEN_11549 = _T_267 ? mip : _GEN_11526; // @[decode.scala 514:28 601:39]
  wire [63:0] _GEN_11550 = _T_267 ? pmpcfg0 : _GEN_11527; // @[decode.scala 515:28 601:39]
  wire [63:0] _GEN_11551 = _T_267 ? pmpaddr0 : _GEN_11528; // @[decode.scala 516:28 601:39]
  wire [63:0] _GEN_11552 = _T_267 ? mvendorid : _GEN_11529; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11553 = _T_267 ? marchid : _GEN_11530; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11554 = _T_267 ? mimpid : _GEN_11531; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11555 = _T_267 ? mhartid : _GEN_11532; // @[decode.scala 520:28 601:39]
  wire [63:0] _GEN_11556 = _T_266 ? _ustatus_T : ustatus; // @[decode.scala 497:28 601:39 602:38]
  wire [63:0] _GEN_11557 = _T_266 ? utvec : _GEN_11533; // @[decode.scala 498:28 601:39]
  wire [63:0] _GEN_11558 = _T_266 ? uepc : _GEN_11534; // @[decode.scala 499:28 601:39]
  wire [63:0] _GEN_11559 = _T_266 ? ucause : _GEN_11535; // @[decode.scala 500:28 601:39]
  wire [63:0] _GEN_11560 = _T_266 ? scounteren : _GEN_11536; // @[decode.scala 501:28 601:39]
  wire [63:0] _GEN_11561 = _T_266 ? satp : _GEN_11537; // @[decode.scala 502:28 601:39]
  wire [63:0] _GEN_11562 = _T_266 ? _mstatus_T_1 : _GEN_11538; // @[decode.scala 522:11 601:39]
  wire [126:0] _GEN_11563 = _T_266 ? 127'h8000000000101101 : _GEN_11539; // @[decode.scala 601:39 523:8]
  wire [63:0] _GEN_11564 = _T_266 ? medeleg : _GEN_11540; // @[decode.scala 505:28 601:39]
  wire [63:0] _GEN_11565 = _T_266 ? mideleg : _GEN_11541; // @[decode.scala 506:28 601:39]
  wire [63:0] _GEN_11566 = _T_266 ? mie : _GEN_11542; // @[decode.scala 507:28 601:39]
  wire [63:0] _GEN_11567 = _T_266 ? mtvec : _GEN_11543; // @[decode.scala 508:28 601:39]
  wire [63:0] _GEN_11568 = _T_266 ? mcounteren : _GEN_11544; // @[decode.scala 509:28 601:39]
  wire [63:0] _GEN_11569 = _T_266 ? mscratch : _GEN_11545; // @[decode.scala 510:28 601:39]
  wire [63:0] _GEN_11570 = _T_266 ? mepc : _GEN_11546; // @[decode.scala 511:28 601:39]
  wire [63:0] _GEN_11571 = _T_266 ? mcause : _GEN_11547; // @[decode.scala 512:28 601:39]
  wire [63:0] _GEN_11572 = _T_266 ? mtval : _GEN_11548; // @[decode.scala 513:28 601:39]
  wire [63:0] _GEN_11573 = _T_266 ? mip : _GEN_11549; // @[decode.scala 514:28 601:39]
  wire [63:0] _GEN_11574 = _T_266 ? pmpcfg0 : _GEN_11550; // @[decode.scala 515:28 601:39]
  wire [63:0] _GEN_11575 = _T_266 ? pmpaddr0 : _GEN_11551; // @[decode.scala 516:28 601:39]
  wire [63:0] _GEN_11576 = _T_266 ? mvendorid : _GEN_11552; // @[decode.scala 517:28 601:39]
  wire [63:0] _GEN_11577 = _T_266 ? marchid : _GEN_11553; // @[decode.scala 518:28 601:39]
  wire [63:0] _GEN_11578 = _T_266 ? mimpid : _GEN_11554; // @[decode.scala 519:28 601:39]
  wire [63:0] _GEN_11579 = _T_266 ? mhartid : _GEN_11555; // @[decode.scala 520:28 601:39]
  wire [63:0] _ustatus_T_1 = ~csrWriteData; // @[decode.scala 630:51]
  wire [63:0] _ustatus_T_2 = ustatus & _ustatus_T_1; // @[decode.scala 630:49]
  wire [63:0] _utvec_T_2 = mtvec & _ustatus_T_1; // @[decode.scala 631:47]
  wire [63:0] _uepc_T_2 = uepc & _ustatus_T_1; // @[decode.scala 632:46]
  wire [63:0] _ucause_T_2 = ucause & _ustatus_T_1; // @[decode.scala 633:48]
  wire [63:0] _scounteren_T_2 = scounteren & _ustatus_T_1; // @[decode.scala 634:52]
  wire [63:0] _satp_T_2 = satp & _ustatus_T_1; // @[decode.scala 635:46]
  wire [63:0] _mstatus_T_4 = mstatus & _ustatus_T_1; // @[decode.scala 636:49]
  wire [63:0] _misa_T_4 = misa & _ustatus_T_1; // @[decode.scala 637:46]
  wire [63:0] _medeleg_T_2 = medeleg & _ustatus_T_1; // @[decode.scala 638:49]
  wire [63:0] _mideleg_T_2 = mideleg & _ustatus_T_1; // @[decode.scala 639:49]
  wire [63:0] _mie_T_2 = mie & _ustatus_T_1; // @[decode.scala 640:45]
  wire [63:0] _mcounteren_T_2 = mcounteren & _ustatus_T_1; // @[decode.scala 642:52]
  wire [63:0] _mscratch_T_2 = mscratch & _ustatus_T_1; // @[decode.scala 643:50]
  wire [63:0] _mepc_T_2 = mepc & _ustatus_T_1; // @[decode.scala 644:46]
  wire [63:0] _mcause_T_2 = mcause & _ustatus_T_1; // @[decode.scala 645:48]
  wire [63:0] _mtval_T_2 = mtval & _ustatus_T_1; // @[decode.scala 646:47]
  wire [63:0] _mip_T_2 = mip & _ustatus_T_1; // @[decode.scala 647:45]
  wire [63:0] _pmpcfg0_T_2 = pmpcfg0 & _ustatus_T_1; // @[decode.scala 648:49]
  wire [63:0] _pmpaddr0_T_2 = pmpaddr0 & _ustatus_T_1; // @[decode.scala 649:50]
  wire [63:0] _mvendorid_T_2 = mvendorid & _ustatus_T_1; // @[decode.scala 650:51]
  wire [63:0] _marchid_T_2 = marchid & _ustatus_T_1; // @[decode.scala 651:49]
  wire [63:0] _mimpid_T_2 = mimpid & _ustatus_T_1; // @[decode.scala 652:48]
  wire [63:0] _mhartid_T_2 = mhartid & _ustatus_T_1; // @[decode.scala 653:49]
  wire [63:0] _GEN_11580 = _T_289 ? _mhartid_T_2 : mhartid; // @[decode.scala 520:28 629:39 653:38]
  wire [63:0] _GEN_11581 = _T_288 ? _mimpid_T_2 : mimpid; // @[decode.scala 519:28 629:39 652:38]
  wire [63:0] _GEN_11582 = _T_288 ? mhartid : _GEN_11580; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11583 = _T_287 ? _marchid_T_2 : marchid; // @[decode.scala 518:28 629:39 651:38]
  wire [63:0] _GEN_11584 = _T_287 ? mimpid : _GEN_11581; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11585 = _T_287 ? mhartid : _GEN_11582; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11586 = _T_286 ? _mvendorid_T_2 : mvendorid; // @[decode.scala 517:28 629:39 650:38]
  wire [63:0] _GEN_11587 = _T_286 ? marchid : _GEN_11583; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11588 = _T_286 ? mimpid : _GEN_11584; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11589 = _T_286 ? mhartid : _GEN_11585; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11590 = _T_285 ? _pmpaddr0_T_2 : pmpaddr0; // @[decode.scala 516:28 629:39 649:38]
  wire [63:0] _GEN_11591 = _T_285 ? mvendorid : _GEN_11586; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11592 = _T_285 ? marchid : _GEN_11587; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11593 = _T_285 ? mimpid : _GEN_11588; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11594 = _T_285 ? mhartid : _GEN_11589; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11595 = _T_284 ? _pmpcfg0_T_2 : pmpcfg0; // @[decode.scala 515:28 629:39 648:38]
  wire [63:0] _GEN_11596 = _T_284 ? pmpaddr0 : _GEN_11590; // @[decode.scala 516:28 629:39]
  wire [63:0] _GEN_11597 = _T_284 ? mvendorid : _GEN_11591; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11598 = _T_284 ? marchid : _GEN_11592; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11599 = _T_284 ? mimpid : _GEN_11593; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11600 = _T_284 ? mhartid : _GEN_11594; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11601 = _T_283 ? _mip_T_2 : mip; // @[decode.scala 514:28 629:39 647:38]
  wire [63:0] _GEN_11602 = _T_283 ? pmpcfg0 : _GEN_11595; // @[decode.scala 515:28 629:39]
  wire [63:0] _GEN_11603 = _T_283 ? pmpaddr0 : _GEN_11596; // @[decode.scala 516:28 629:39]
  wire [63:0] _GEN_11604 = _T_283 ? mvendorid : _GEN_11597; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11605 = _T_283 ? marchid : _GEN_11598; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11606 = _T_283 ? mimpid : _GEN_11599; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11607 = _T_283 ? mhartid : _GEN_11600; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11608 = _T_282 ? _mtval_T_2 : mtval; // @[decode.scala 513:28 629:39 646:38]
  wire [63:0] _GEN_11609 = _T_282 ? mip : _GEN_11601; // @[decode.scala 514:28 629:39]
  wire [63:0] _GEN_11610 = _T_282 ? pmpcfg0 : _GEN_11602; // @[decode.scala 515:28 629:39]
  wire [63:0] _GEN_11611 = _T_282 ? pmpaddr0 : _GEN_11603; // @[decode.scala 516:28 629:39]
  wire [63:0] _GEN_11612 = _T_282 ? mvendorid : _GEN_11604; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11613 = _T_282 ? marchid : _GEN_11605; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11614 = _T_282 ? mimpid : _GEN_11606; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11615 = _T_282 ? mhartid : _GEN_11607; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11616 = _T_281 ? _mcause_T_2 : mcause; // @[decode.scala 512:28 629:39 645:38]
  wire [63:0] _GEN_11617 = _T_281 ? mtval : _GEN_11608; // @[decode.scala 513:28 629:39]
  wire [63:0] _GEN_11618 = _T_281 ? mip : _GEN_11609; // @[decode.scala 514:28 629:39]
  wire [63:0] _GEN_11619 = _T_281 ? pmpcfg0 : _GEN_11610; // @[decode.scala 515:28 629:39]
  wire [63:0] _GEN_11620 = _T_281 ? pmpaddr0 : _GEN_11611; // @[decode.scala 516:28 629:39]
  wire [63:0] _GEN_11621 = _T_281 ? mvendorid : _GEN_11612; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11622 = _T_281 ? marchid : _GEN_11613; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11623 = _T_281 ? mimpid : _GEN_11614; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11624 = _T_281 ? mhartid : _GEN_11615; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11625 = _T_280 ? _mepc_T_2 : mepc; // @[decode.scala 511:28 629:39 644:38]
  wire [63:0] _GEN_11626 = _T_280 ? mcause : _GEN_11616; // @[decode.scala 512:28 629:39]
  wire [63:0] _GEN_11627 = _T_280 ? mtval : _GEN_11617; // @[decode.scala 513:28 629:39]
  wire [63:0] _GEN_11628 = _T_280 ? mip : _GEN_11618; // @[decode.scala 514:28 629:39]
  wire [63:0] _GEN_11629 = _T_280 ? pmpcfg0 : _GEN_11619; // @[decode.scala 515:28 629:39]
  wire [63:0] _GEN_11630 = _T_280 ? pmpaddr0 : _GEN_11620; // @[decode.scala 516:28 629:39]
  wire [63:0] _GEN_11631 = _T_280 ? mvendorid : _GEN_11621; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11632 = _T_280 ? marchid : _GEN_11622; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11633 = _T_280 ? mimpid : _GEN_11623; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11634 = _T_280 ? mhartid : _GEN_11624; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11635 = _T_279 ? _mscratch_T_2 : mscratch; // @[decode.scala 510:28 629:39 643:38]
  wire [63:0] _GEN_11636 = _T_279 ? mepc : _GEN_11625; // @[decode.scala 511:28 629:39]
  wire [63:0] _GEN_11637 = _T_279 ? mcause : _GEN_11626; // @[decode.scala 512:28 629:39]
  wire [63:0] _GEN_11638 = _T_279 ? mtval : _GEN_11627; // @[decode.scala 513:28 629:39]
  wire [63:0] _GEN_11639 = _T_279 ? mip : _GEN_11628; // @[decode.scala 514:28 629:39]
  wire [63:0] _GEN_11640 = _T_279 ? pmpcfg0 : _GEN_11629; // @[decode.scala 515:28 629:39]
  wire [63:0] _GEN_11641 = _T_279 ? pmpaddr0 : _GEN_11630; // @[decode.scala 516:28 629:39]
  wire [63:0] _GEN_11642 = _T_279 ? mvendorid : _GEN_11631; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11643 = _T_279 ? marchid : _GEN_11632; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11644 = _T_279 ? mimpid : _GEN_11633; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11645 = _T_279 ? mhartid : _GEN_11634; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11646 = _T_278 ? _mcounteren_T_2 : mcounteren; // @[decode.scala 509:28 629:39 642:38]
  wire [63:0] _GEN_11647 = _T_278 ? mscratch : _GEN_11635; // @[decode.scala 510:28 629:39]
  wire [63:0] _GEN_11648 = _T_278 ? mepc : _GEN_11636; // @[decode.scala 511:28 629:39]
  wire [63:0] _GEN_11649 = _T_278 ? mcause : _GEN_11637; // @[decode.scala 512:28 629:39]
  wire [63:0] _GEN_11650 = _T_278 ? mtval : _GEN_11638; // @[decode.scala 513:28 629:39]
  wire [63:0] _GEN_11651 = _T_278 ? mip : _GEN_11639; // @[decode.scala 514:28 629:39]
  wire [63:0] _GEN_11652 = _T_278 ? pmpcfg0 : _GEN_11640; // @[decode.scala 515:28 629:39]
  wire [63:0] _GEN_11653 = _T_278 ? pmpaddr0 : _GEN_11641; // @[decode.scala 516:28 629:39]
  wire [63:0] _GEN_11654 = _T_278 ? mvendorid : _GEN_11642; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11655 = _T_278 ? marchid : _GEN_11643; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11656 = _T_278 ? mimpid : _GEN_11644; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11657 = _T_278 ? mhartid : _GEN_11645; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11658 = _T_277 ? _utvec_T_2 : mtvec; // @[decode.scala 508:28 629:39 641:38]
  wire [63:0] _GEN_11659 = _T_277 ? mcounteren : _GEN_11646; // @[decode.scala 509:28 629:39]
  wire [63:0] _GEN_11660 = _T_277 ? mscratch : _GEN_11647; // @[decode.scala 510:28 629:39]
  wire [63:0] _GEN_11661 = _T_277 ? mepc : _GEN_11648; // @[decode.scala 511:28 629:39]
  wire [63:0] _GEN_11662 = _T_277 ? mcause : _GEN_11649; // @[decode.scala 512:28 629:39]
  wire [63:0] _GEN_11663 = _T_277 ? mtval : _GEN_11650; // @[decode.scala 513:28 629:39]
  wire [63:0] _GEN_11664 = _T_277 ? mip : _GEN_11651; // @[decode.scala 514:28 629:39]
  wire [63:0] _GEN_11665 = _T_277 ? pmpcfg0 : _GEN_11652; // @[decode.scala 515:28 629:39]
  wire [63:0] _GEN_11666 = _T_277 ? pmpaddr0 : _GEN_11653; // @[decode.scala 516:28 629:39]
  wire [63:0] _GEN_11667 = _T_277 ? mvendorid : _GEN_11654; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11668 = _T_277 ? marchid : _GEN_11655; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11669 = _T_277 ? mimpid : _GEN_11656; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11670 = _T_277 ? mhartid : _GEN_11657; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11671 = _T_276 ? _mie_T_2 : mie; // @[decode.scala 507:28 629:39 640:38]
  wire [63:0] _GEN_11672 = _T_276 ? mtvec : _GEN_11658; // @[decode.scala 508:28 629:39]
  wire [63:0] _GEN_11673 = _T_276 ? mcounteren : _GEN_11659; // @[decode.scala 509:28 629:39]
  wire [63:0] _GEN_11674 = _T_276 ? mscratch : _GEN_11660; // @[decode.scala 510:28 629:39]
  wire [63:0] _GEN_11675 = _T_276 ? mepc : _GEN_11661; // @[decode.scala 511:28 629:39]
  wire [63:0] _GEN_11676 = _T_276 ? mcause : _GEN_11662; // @[decode.scala 512:28 629:39]
  wire [63:0] _GEN_11677 = _T_276 ? mtval : _GEN_11663; // @[decode.scala 513:28 629:39]
  wire [63:0] _GEN_11678 = _T_276 ? mip : _GEN_11664; // @[decode.scala 514:28 629:39]
  wire [63:0] _GEN_11679 = _T_276 ? pmpcfg0 : _GEN_11665; // @[decode.scala 515:28 629:39]
  wire [63:0] _GEN_11680 = _T_276 ? pmpaddr0 : _GEN_11666; // @[decode.scala 516:28 629:39]
  wire [63:0] _GEN_11681 = _T_276 ? mvendorid : _GEN_11667; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11682 = _T_276 ? marchid : _GEN_11668; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11683 = _T_276 ? mimpid : _GEN_11669; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11684 = _T_276 ? mhartid : _GEN_11670; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11685 = _T_275 ? _mideleg_T_2 : mideleg; // @[decode.scala 506:28 629:39 639:38]
  wire [63:0] _GEN_11686 = _T_275 ? mie : _GEN_11671; // @[decode.scala 507:28 629:39]
  wire [63:0] _GEN_11687 = _T_275 ? mtvec : _GEN_11672; // @[decode.scala 508:28 629:39]
  wire [63:0] _GEN_11688 = _T_275 ? mcounteren : _GEN_11673; // @[decode.scala 509:28 629:39]
  wire [63:0] _GEN_11689 = _T_275 ? mscratch : _GEN_11674; // @[decode.scala 510:28 629:39]
  wire [63:0] _GEN_11690 = _T_275 ? mepc : _GEN_11675; // @[decode.scala 511:28 629:39]
  wire [63:0] _GEN_11691 = _T_275 ? mcause : _GEN_11676; // @[decode.scala 512:28 629:39]
  wire [63:0] _GEN_11692 = _T_275 ? mtval : _GEN_11677; // @[decode.scala 513:28 629:39]
  wire [63:0] _GEN_11693 = _T_275 ? mip : _GEN_11678; // @[decode.scala 514:28 629:39]
  wire [63:0] _GEN_11694 = _T_275 ? pmpcfg0 : _GEN_11679; // @[decode.scala 515:28 629:39]
  wire [63:0] _GEN_11695 = _T_275 ? pmpaddr0 : _GEN_11680; // @[decode.scala 516:28 629:39]
  wire [63:0] _GEN_11696 = _T_275 ? mvendorid : _GEN_11681; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11697 = _T_275 ? marchid : _GEN_11682; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11698 = _T_275 ? mimpid : _GEN_11683; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11699 = _T_275 ? mhartid : _GEN_11684; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11700 = _T_274 ? _medeleg_T_2 : medeleg; // @[decode.scala 505:28 629:39 638:38]
  wire [63:0] _GEN_11701 = _T_274 ? mideleg : _GEN_11685; // @[decode.scala 506:28 629:39]
  wire [63:0] _GEN_11702 = _T_274 ? mie : _GEN_11686; // @[decode.scala 507:28 629:39]
  wire [63:0] _GEN_11703 = _T_274 ? mtvec : _GEN_11687; // @[decode.scala 508:28 629:39]
  wire [63:0] _GEN_11704 = _T_274 ? mcounteren : _GEN_11688; // @[decode.scala 509:28 629:39]
  wire [63:0] _GEN_11705 = _T_274 ? mscratch : _GEN_11689; // @[decode.scala 510:28 629:39]
  wire [63:0] _GEN_11706 = _T_274 ? mepc : _GEN_11690; // @[decode.scala 511:28 629:39]
  wire [63:0] _GEN_11707 = _T_274 ? mcause : _GEN_11691; // @[decode.scala 512:28 629:39]
  wire [63:0] _GEN_11708 = _T_274 ? mtval : _GEN_11692; // @[decode.scala 513:28 629:39]
  wire [63:0] _GEN_11709 = _T_274 ? mip : _GEN_11693; // @[decode.scala 514:28 629:39]
  wire [63:0] _GEN_11710 = _T_274 ? pmpcfg0 : _GEN_11694; // @[decode.scala 515:28 629:39]
  wire [63:0] _GEN_11711 = _T_274 ? pmpaddr0 : _GEN_11695; // @[decode.scala 516:28 629:39]
  wire [63:0] _GEN_11712 = _T_274 ? mvendorid : _GEN_11696; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11713 = _T_274 ? marchid : _GEN_11697; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11714 = _T_274 ? mimpid : _GEN_11698; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11715 = _T_274 ? mhartid : _GEN_11699; // @[decode.scala 520:28 629:39]
  wire [126:0] _GEN_11716 = _T_273 ? {{63'd0}, _misa_T_4} : 127'h8000000000101101; // @[decode.scala 629:39 637:38 523:8]
  wire [63:0] _GEN_11717 = _T_273 ? medeleg : _GEN_11700; // @[decode.scala 505:28 629:39]
  wire [63:0] _GEN_11718 = _T_273 ? mideleg : _GEN_11701; // @[decode.scala 506:28 629:39]
  wire [63:0] _GEN_11719 = _T_273 ? mie : _GEN_11702; // @[decode.scala 507:28 629:39]
  wire [63:0] _GEN_11720 = _T_273 ? mtvec : _GEN_11703; // @[decode.scala 508:28 629:39]
  wire [63:0] _GEN_11721 = _T_273 ? mcounteren : _GEN_11704; // @[decode.scala 509:28 629:39]
  wire [63:0] _GEN_11722 = _T_273 ? mscratch : _GEN_11705; // @[decode.scala 510:28 629:39]
  wire [63:0] _GEN_11723 = _T_273 ? mepc : _GEN_11706; // @[decode.scala 511:28 629:39]
  wire [63:0] _GEN_11724 = _T_273 ? mcause : _GEN_11707; // @[decode.scala 512:28 629:39]
  wire [63:0] _GEN_11725 = _T_273 ? mtval : _GEN_11708; // @[decode.scala 513:28 629:39]
  wire [63:0] _GEN_11726 = _T_273 ? mip : _GEN_11709; // @[decode.scala 514:28 629:39]
  wire [63:0] _GEN_11727 = _T_273 ? pmpcfg0 : _GEN_11710; // @[decode.scala 515:28 629:39]
  wire [63:0] _GEN_11728 = _T_273 ? pmpaddr0 : _GEN_11711; // @[decode.scala 516:28 629:39]
  wire [63:0] _GEN_11729 = _T_273 ? mvendorid : _GEN_11712; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11730 = _T_273 ? marchid : _GEN_11713; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11731 = _T_273 ? mimpid : _GEN_11714; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11732 = _T_273 ? mhartid : _GEN_11715; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11733 = _T_272 ? _mstatus_T_4 : _mstatus_T_1; // @[decode.scala 522:11 629:39 636:38]
  wire [126:0] _GEN_11734 = _T_272 ? 127'h8000000000101101 : _GEN_11716; // @[decode.scala 629:39 523:8]
  wire [63:0] _GEN_11735 = _T_272 ? medeleg : _GEN_11717; // @[decode.scala 505:28 629:39]
  wire [63:0] _GEN_11736 = _T_272 ? mideleg : _GEN_11718; // @[decode.scala 506:28 629:39]
  wire [63:0] _GEN_11737 = _T_272 ? mie : _GEN_11719; // @[decode.scala 507:28 629:39]
  wire [63:0] _GEN_11738 = _T_272 ? mtvec : _GEN_11720; // @[decode.scala 508:28 629:39]
  wire [63:0] _GEN_11739 = _T_272 ? mcounteren : _GEN_11721; // @[decode.scala 509:28 629:39]
  wire [63:0] _GEN_11740 = _T_272 ? mscratch : _GEN_11722; // @[decode.scala 510:28 629:39]
  wire [63:0] _GEN_11741 = _T_272 ? mepc : _GEN_11723; // @[decode.scala 511:28 629:39]
  wire [63:0] _GEN_11742 = _T_272 ? mcause : _GEN_11724; // @[decode.scala 512:28 629:39]
  wire [63:0] _GEN_11743 = _T_272 ? mtval : _GEN_11725; // @[decode.scala 513:28 629:39]
  wire [63:0] _GEN_11744 = _T_272 ? mip : _GEN_11726; // @[decode.scala 514:28 629:39]
  wire [63:0] _GEN_11745 = _T_272 ? pmpcfg0 : _GEN_11727; // @[decode.scala 515:28 629:39]
  wire [63:0] _GEN_11746 = _T_272 ? pmpaddr0 : _GEN_11728; // @[decode.scala 516:28 629:39]
  wire [63:0] _GEN_11747 = _T_272 ? mvendorid : _GEN_11729; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11748 = _T_272 ? marchid : _GEN_11730; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11749 = _T_272 ? mimpid : _GEN_11731; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11750 = _T_272 ? mhartid : _GEN_11732; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11751 = _T_271 ? _satp_T_2 : satp; // @[decode.scala 502:28 629:39 635:38]
  wire [63:0] _GEN_11752 = _T_271 ? _mstatus_T_1 : _GEN_11733; // @[decode.scala 522:11 629:39]
  wire [126:0] _GEN_11753 = _T_271 ? 127'h8000000000101101 : _GEN_11734; // @[decode.scala 629:39 523:8]
  wire [63:0] _GEN_11754 = _T_271 ? medeleg : _GEN_11735; // @[decode.scala 505:28 629:39]
  wire [63:0] _GEN_11755 = _T_271 ? mideleg : _GEN_11736; // @[decode.scala 506:28 629:39]
  wire [63:0] _GEN_11756 = _T_271 ? mie : _GEN_11737; // @[decode.scala 507:28 629:39]
  wire [63:0] _GEN_11757 = _T_271 ? mtvec : _GEN_11738; // @[decode.scala 508:28 629:39]
  wire [63:0] _GEN_11758 = _T_271 ? mcounteren : _GEN_11739; // @[decode.scala 509:28 629:39]
  wire [63:0] _GEN_11759 = _T_271 ? mscratch : _GEN_11740; // @[decode.scala 510:28 629:39]
  wire [63:0] _GEN_11760 = _T_271 ? mepc : _GEN_11741; // @[decode.scala 511:28 629:39]
  wire [63:0] _GEN_11761 = _T_271 ? mcause : _GEN_11742; // @[decode.scala 512:28 629:39]
  wire [63:0] _GEN_11762 = _T_271 ? mtval : _GEN_11743; // @[decode.scala 513:28 629:39]
  wire [63:0] _GEN_11763 = _T_271 ? mip : _GEN_11744; // @[decode.scala 514:28 629:39]
  wire [63:0] _GEN_11764 = _T_271 ? pmpcfg0 : _GEN_11745; // @[decode.scala 515:28 629:39]
  wire [63:0] _GEN_11765 = _T_271 ? pmpaddr0 : _GEN_11746; // @[decode.scala 516:28 629:39]
  wire [63:0] _GEN_11766 = _T_271 ? mvendorid : _GEN_11747; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11767 = _T_271 ? marchid : _GEN_11748; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11768 = _T_271 ? mimpid : _GEN_11749; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11769 = _T_271 ? mhartid : _GEN_11750; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11770 = _T_270 ? _scounteren_T_2 : scounteren; // @[decode.scala 501:28 629:39 634:38]
  wire [63:0] _GEN_11771 = _T_270 ? satp : _GEN_11751; // @[decode.scala 502:28 629:39]
  wire [63:0] _GEN_11772 = _T_270 ? _mstatus_T_1 : _GEN_11752; // @[decode.scala 522:11 629:39]
  wire [126:0] _GEN_11773 = _T_270 ? 127'h8000000000101101 : _GEN_11753; // @[decode.scala 629:39 523:8]
  wire [63:0] _GEN_11774 = _T_270 ? medeleg : _GEN_11754; // @[decode.scala 505:28 629:39]
  wire [63:0] _GEN_11775 = _T_270 ? mideleg : _GEN_11755; // @[decode.scala 506:28 629:39]
  wire [63:0] _GEN_11776 = _T_270 ? mie : _GEN_11756; // @[decode.scala 507:28 629:39]
  wire [63:0] _GEN_11777 = _T_270 ? mtvec : _GEN_11757; // @[decode.scala 508:28 629:39]
  wire [63:0] _GEN_11778 = _T_270 ? mcounteren : _GEN_11758; // @[decode.scala 509:28 629:39]
  wire [63:0] _GEN_11779 = _T_270 ? mscratch : _GEN_11759; // @[decode.scala 510:28 629:39]
  wire [63:0] _GEN_11780 = _T_270 ? mepc : _GEN_11760; // @[decode.scala 511:28 629:39]
  wire [63:0] _GEN_11781 = _T_270 ? mcause : _GEN_11761; // @[decode.scala 512:28 629:39]
  wire [63:0] _GEN_11782 = _T_270 ? mtval : _GEN_11762; // @[decode.scala 513:28 629:39]
  wire [63:0] _GEN_11783 = _T_270 ? mip : _GEN_11763; // @[decode.scala 514:28 629:39]
  wire [63:0] _GEN_11784 = _T_270 ? pmpcfg0 : _GEN_11764; // @[decode.scala 515:28 629:39]
  wire [63:0] _GEN_11785 = _T_270 ? pmpaddr0 : _GEN_11765; // @[decode.scala 516:28 629:39]
  wire [63:0] _GEN_11786 = _T_270 ? mvendorid : _GEN_11766; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11787 = _T_270 ? marchid : _GEN_11767; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11788 = _T_270 ? mimpid : _GEN_11768; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11789 = _T_270 ? mhartid : _GEN_11769; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11790 = _T_269 ? _ucause_T_2 : ucause; // @[decode.scala 500:28 629:39 633:38]
  wire [63:0] _GEN_11791 = _T_269 ? scounteren : _GEN_11770; // @[decode.scala 501:28 629:39]
  wire [63:0] _GEN_11792 = _T_269 ? satp : _GEN_11771; // @[decode.scala 502:28 629:39]
  wire [63:0] _GEN_11793 = _T_269 ? _mstatus_T_1 : _GEN_11772; // @[decode.scala 522:11 629:39]
  wire [126:0] _GEN_11794 = _T_269 ? 127'h8000000000101101 : _GEN_11773; // @[decode.scala 629:39 523:8]
  wire [63:0] _GEN_11795 = _T_269 ? medeleg : _GEN_11774; // @[decode.scala 505:28 629:39]
  wire [63:0] _GEN_11796 = _T_269 ? mideleg : _GEN_11775; // @[decode.scala 506:28 629:39]
  wire [63:0] _GEN_11797 = _T_269 ? mie : _GEN_11776; // @[decode.scala 507:28 629:39]
  wire [63:0] _GEN_11798 = _T_269 ? mtvec : _GEN_11777; // @[decode.scala 508:28 629:39]
  wire [63:0] _GEN_11799 = _T_269 ? mcounteren : _GEN_11778; // @[decode.scala 509:28 629:39]
  wire [63:0] _GEN_11800 = _T_269 ? mscratch : _GEN_11779; // @[decode.scala 510:28 629:39]
  wire [63:0] _GEN_11801 = _T_269 ? mepc : _GEN_11780; // @[decode.scala 511:28 629:39]
  wire [63:0] _GEN_11802 = _T_269 ? mcause : _GEN_11781; // @[decode.scala 512:28 629:39]
  wire [63:0] _GEN_11803 = _T_269 ? mtval : _GEN_11782; // @[decode.scala 513:28 629:39]
  wire [63:0] _GEN_11804 = _T_269 ? mip : _GEN_11783; // @[decode.scala 514:28 629:39]
  wire [63:0] _GEN_11805 = _T_269 ? pmpcfg0 : _GEN_11784; // @[decode.scala 515:28 629:39]
  wire [63:0] _GEN_11806 = _T_269 ? pmpaddr0 : _GEN_11785; // @[decode.scala 516:28 629:39]
  wire [63:0] _GEN_11807 = _T_269 ? mvendorid : _GEN_11786; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11808 = _T_269 ? marchid : _GEN_11787; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11809 = _T_269 ? mimpid : _GEN_11788; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11810 = _T_269 ? mhartid : _GEN_11789; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11811 = _T_268 ? _uepc_T_2 : uepc; // @[decode.scala 499:28 629:39 632:38]
  wire [63:0] _GEN_11812 = _T_268 ? ucause : _GEN_11790; // @[decode.scala 500:28 629:39]
  wire [63:0] _GEN_11813 = _T_268 ? scounteren : _GEN_11791; // @[decode.scala 501:28 629:39]
  wire [63:0] _GEN_11814 = _T_268 ? satp : _GEN_11792; // @[decode.scala 502:28 629:39]
  wire [63:0] _GEN_11815 = _T_268 ? _mstatus_T_1 : _GEN_11793; // @[decode.scala 522:11 629:39]
  wire [126:0] _GEN_11816 = _T_268 ? 127'h8000000000101101 : _GEN_11794; // @[decode.scala 629:39 523:8]
  wire [63:0] _GEN_11817 = _T_268 ? medeleg : _GEN_11795; // @[decode.scala 505:28 629:39]
  wire [63:0] _GEN_11818 = _T_268 ? mideleg : _GEN_11796; // @[decode.scala 506:28 629:39]
  wire [63:0] _GEN_11819 = _T_268 ? mie : _GEN_11797; // @[decode.scala 507:28 629:39]
  wire [63:0] _GEN_11820 = _T_268 ? mtvec : _GEN_11798; // @[decode.scala 508:28 629:39]
  wire [63:0] _GEN_11821 = _T_268 ? mcounteren : _GEN_11799; // @[decode.scala 509:28 629:39]
  wire [63:0] _GEN_11822 = _T_268 ? mscratch : _GEN_11800; // @[decode.scala 510:28 629:39]
  wire [63:0] _GEN_11823 = _T_268 ? mepc : _GEN_11801; // @[decode.scala 511:28 629:39]
  wire [63:0] _GEN_11824 = _T_268 ? mcause : _GEN_11802; // @[decode.scala 512:28 629:39]
  wire [63:0] _GEN_11825 = _T_268 ? mtval : _GEN_11803; // @[decode.scala 513:28 629:39]
  wire [63:0] _GEN_11826 = _T_268 ? mip : _GEN_11804; // @[decode.scala 514:28 629:39]
  wire [63:0] _GEN_11827 = _T_268 ? pmpcfg0 : _GEN_11805; // @[decode.scala 515:28 629:39]
  wire [63:0] _GEN_11828 = _T_268 ? pmpaddr0 : _GEN_11806; // @[decode.scala 516:28 629:39]
  wire [63:0] _GEN_11829 = _T_268 ? mvendorid : _GEN_11807; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11830 = _T_268 ? marchid : _GEN_11808; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11831 = _T_268 ? mimpid : _GEN_11809; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11832 = _T_268 ? mhartid : _GEN_11810; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11833 = _T_267 ? _utvec_T_2 : utvec; // @[decode.scala 498:28 629:39 631:38]
  wire [63:0] _GEN_11834 = _T_267 ? uepc : _GEN_11811; // @[decode.scala 499:28 629:39]
  wire [63:0] _GEN_11835 = _T_267 ? ucause : _GEN_11812; // @[decode.scala 500:28 629:39]
  wire [63:0] _GEN_11836 = _T_267 ? scounteren : _GEN_11813; // @[decode.scala 501:28 629:39]
  wire [63:0] _GEN_11837 = _T_267 ? satp : _GEN_11814; // @[decode.scala 502:28 629:39]
  wire [63:0] _GEN_11838 = _T_267 ? _mstatus_T_1 : _GEN_11815; // @[decode.scala 522:11 629:39]
  wire [126:0] _GEN_11839 = _T_267 ? 127'h8000000000101101 : _GEN_11816; // @[decode.scala 629:39 523:8]
  wire [63:0] _GEN_11840 = _T_267 ? medeleg : _GEN_11817; // @[decode.scala 505:28 629:39]
  wire [63:0] _GEN_11841 = _T_267 ? mideleg : _GEN_11818; // @[decode.scala 506:28 629:39]
  wire [63:0] _GEN_11842 = _T_267 ? mie : _GEN_11819; // @[decode.scala 507:28 629:39]
  wire [63:0] _GEN_11843 = _T_267 ? mtvec : _GEN_11820; // @[decode.scala 508:28 629:39]
  wire [63:0] _GEN_11844 = _T_267 ? mcounteren : _GEN_11821; // @[decode.scala 509:28 629:39]
  wire [63:0] _GEN_11845 = _T_267 ? mscratch : _GEN_11822; // @[decode.scala 510:28 629:39]
  wire [63:0] _GEN_11846 = _T_267 ? mepc : _GEN_11823; // @[decode.scala 511:28 629:39]
  wire [63:0] _GEN_11847 = _T_267 ? mcause : _GEN_11824; // @[decode.scala 512:28 629:39]
  wire [63:0] _GEN_11848 = _T_267 ? mtval : _GEN_11825; // @[decode.scala 513:28 629:39]
  wire [63:0] _GEN_11849 = _T_267 ? mip : _GEN_11826; // @[decode.scala 514:28 629:39]
  wire [63:0] _GEN_11850 = _T_267 ? pmpcfg0 : _GEN_11827; // @[decode.scala 515:28 629:39]
  wire [63:0] _GEN_11851 = _T_267 ? pmpaddr0 : _GEN_11828; // @[decode.scala 516:28 629:39]
  wire [63:0] _GEN_11852 = _T_267 ? mvendorid : _GEN_11829; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11853 = _T_267 ? marchid : _GEN_11830; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11854 = _T_267 ? mimpid : _GEN_11831; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11855 = _T_267 ? mhartid : _GEN_11832; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11856 = _T_266 ? _ustatus_T_2 : ustatus; // @[decode.scala 497:28 629:39 630:38]
  wire [63:0] _GEN_11857 = _T_266 ? utvec : _GEN_11833; // @[decode.scala 498:28 629:39]
  wire [63:0] _GEN_11858 = _T_266 ? uepc : _GEN_11834; // @[decode.scala 499:28 629:39]
  wire [63:0] _GEN_11859 = _T_266 ? ucause : _GEN_11835; // @[decode.scala 500:28 629:39]
  wire [63:0] _GEN_11860 = _T_266 ? scounteren : _GEN_11836; // @[decode.scala 501:28 629:39]
  wire [63:0] _GEN_11861 = _T_266 ? satp : _GEN_11837; // @[decode.scala 502:28 629:39]
  wire [63:0] _GEN_11862 = _T_266 ? _mstatus_T_1 : _GEN_11838; // @[decode.scala 522:11 629:39]
  wire [126:0] _GEN_11863 = _T_266 ? 127'h8000000000101101 : _GEN_11839; // @[decode.scala 629:39 523:8]
  wire [63:0] _GEN_11864 = _T_266 ? medeleg : _GEN_11840; // @[decode.scala 505:28 629:39]
  wire [63:0] _GEN_11865 = _T_266 ? mideleg : _GEN_11841; // @[decode.scala 506:28 629:39]
  wire [63:0] _GEN_11866 = _T_266 ? mie : _GEN_11842; // @[decode.scala 507:28 629:39]
  wire [63:0] _GEN_11867 = _T_266 ? mtvec : _GEN_11843; // @[decode.scala 508:28 629:39]
  wire [63:0] _GEN_11868 = _T_266 ? mcounteren : _GEN_11844; // @[decode.scala 509:28 629:39]
  wire [63:0] _GEN_11869 = _T_266 ? mscratch : _GEN_11845; // @[decode.scala 510:28 629:39]
  wire [63:0] _GEN_11870 = _T_266 ? mepc : _GEN_11846; // @[decode.scala 511:28 629:39]
  wire [63:0] _GEN_11871 = _T_266 ? mcause : _GEN_11847; // @[decode.scala 512:28 629:39]
  wire [63:0] _GEN_11872 = _T_266 ? mtval : _GEN_11848; // @[decode.scala 513:28 629:39]
  wire [63:0] _GEN_11873 = _T_266 ? mip : _GEN_11849; // @[decode.scala 514:28 629:39]
  wire [63:0] _GEN_11874 = _T_266 ? pmpcfg0 : _GEN_11850; // @[decode.scala 515:28 629:39]
  wire [63:0] _GEN_11875 = _T_266 ? pmpaddr0 : _GEN_11851; // @[decode.scala 516:28 629:39]
  wire [63:0] _GEN_11876 = _T_266 ? mvendorid : _GEN_11852; // @[decode.scala 517:28 629:39]
  wire [63:0] _GEN_11877 = _T_266 ? marchid : _GEN_11853; // @[decode.scala 518:28 629:39]
  wire [63:0] _GEN_11878 = _T_266 ? mimpid : _GEN_11854; // @[decode.scala 519:28 629:39]
  wire [63:0] _GEN_11879 = _T_266 ? mhartid : _GEN_11855; // @[decode.scala 520:28 629:39]
  wire [63:0] _GEN_11880 = _T_289 ? csrImmReg : mhartid; // @[decode.scala 520:28 657:39 681:38]
  wire [63:0] _GEN_11881 = _T_288 ? csrImmReg : mimpid; // @[decode.scala 519:28 657:39 680:38]
  wire [63:0] _GEN_11882 = _T_288 ? mhartid : _GEN_11880; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_11883 = _T_287 ? csrImmReg : marchid; // @[decode.scala 518:28 657:39 679:38]
  wire [63:0] _GEN_11884 = _T_287 ? mimpid : _GEN_11881; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_11885 = _T_287 ? mhartid : _GEN_11882; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_11886 = _T_286 ? csrImmReg : mvendorid; // @[decode.scala 517:28 657:39 678:38]
  wire [63:0] _GEN_11887 = _T_286 ? marchid : _GEN_11883; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_11888 = _T_286 ? mimpid : _GEN_11884; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_11889 = _T_286 ? mhartid : _GEN_11885; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_11890 = _T_285 ? csrImmReg : pmpaddr0; // @[decode.scala 516:28 657:39 677:38]
  wire [63:0] _GEN_11891 = _T_285 ? mvendorid : _GEN_11886; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_11892 = _T_285 ? marchid : _GEN_11887; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_11893 = _T_285 ? mimpid : _GEN_11888; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_11894 = _T_285 ? mhartid : _GEN_11889; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_11895 = _T_284 ? csrImmReg : pmpcfg0; // @[decode.scala 515:28 657:39 676:38]
  wire [63:0] _GEN_11896 = _T_284 ? pmpaddr0 : _GEN_11890; // @[decode.scala 516:28 657:39]
  wire [63:0] _GEN_11897 = _T_284 ? mvendorid : _GEN_11891; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_11898 = _T_284 ? marchid : _GEN_11892; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_11899 = _T_284 ? mimpid : _GEN_11893; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_11900 = _T_284 ? mhartid : _GEN_11894; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_11901 = _T_283 ? csrImmReg : mip; // @[decode.scala 514:28 657:39 675:38]
  wire [63:0] _GEN_11902 = _T_283 ? pmpcfg0 : _GEN_11895; // @[decode.scala 515:28 657:39]
  wire [63:0] _GEN_11903 = _T_283 ? pmpaddr0 : _GEN_11896; // @[decode.scala 516:28 657:39]
  wire [63:0] _GEN_11904 = _T_283 ? mvendorid : _GEN_11897; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_11905 = _T_283 ? marchid : _GEN_11898; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_11906 = _T_283 ? mimpid : _GEN_11899; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_11907 = _T_283 ? mhartid : _GEN_11900; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_11908 = _T_282 ? csrImmReg : mtval; // @[decode.scala 513:28 657:39 674:38]
  wire [63:0] _GEN_11909 = _T_282 ? mip : _GEN_11901; // @[decode.scala 514:28 657:39]
  wire [63:0] _GEN_11910 = _T_282 ? pmpcfg0 : _GEN_11902; // @[decode.scala 515:28 657:39]
  wire [63:0] _GEN_11911 = _T_282 ? pmpaddr0 : _GEN_11903; // @[decode.scala 516:28 657:39]
  wire [63:0] _GEN_11912 = _T_282 ? mvendorid : _GEN_11904; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_11913 = _T_282 ? marchid : _GEN_11905; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_11914 = _T_282 ? mimpid : _GEN_11906; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_11915 = _T_282 ? mhartid : _GEN_11907; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_11916 = _T_281 ? csrImmReg : mcause; // @[decode.scala 512:28 657:39 673:38]
  wire [63:0] _GEN_11917 = _T_281 ? mtval : _GEN_11908; // @[decode.scala 513:28 657:39]
  wire [63:0] _GEN_11918 = _T_281 ? mip : _GEN_11909; // @[decode.scala 514:28 657:39]
  wire [63:0] _GEN_11919 = _T_281 ? pmpcfg0 : _GEN_11910; // @[decode.scala 515:28 657:39]
  wire [63:0] _GEN_11920 = _T_281 ? pmpaddr0 : _GEN_11911; // @[decode.scala 516:28 657:39]
  wire [63:0] _GEN_11921 = _T_281 ? mvendorid : _GEN_11912; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_11922 = _T_281 ? marchid : _GEN_11913; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_11923 = _T_281 ? mimpid : _GEN_11914; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_11924 = _T_281 ? mhartid : _GEN_11915; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_11925 = _T_280 ? csrImmReg : mepc; // @[decode.scala 511:28 657:39 672:38]
  wire [63:0] _GEN_11926 = _T_280 ? mcause : _GEN_11916; // @[decode.scala 512:28 657:39]
  wire [63:0] _GEN_11927 = _T_280 ? mtval : _GEN_11917; // @[decode.scala 513:28 657:39]
  wire [63:0] _GEN_11928 = _T_280 ? mip : _GEN_11918; // @[decode.scala 514:28 657:39]
  wire [63:0] _GEN_11929 = _T_280 ? pmpcfg0 : _GEN_11919; // @[decode.scala 515:28 657:39]
  wire [63:0] _GEN_11930 = _T_280 ? pmpaddr0 : _GEN_11920; // @[decode.scala 516:28 657:39]
  wire [63:0] _GEN_11931 = _T_280 ? mvendorid : _GEN_11921; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_11932 = _T_280 ? marchid : _GEN_11922; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_11933 = _T_280 ? mimpid : _GEN_11923; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_11934 = _T_280 ? mhartid : _GEN_11924; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_11935 = _T_279 ? csrImmReg : mscratch; // @[decode.scala 510:28 657:39 671:38]
  wire [63:0] _GEN_11936 = _T_279 ? mepc : _GEN_11925; // @[decode.scala 511:28 657:39]
  wire [63:0] _GEN_11937 = _T_279 ? mcause : _GEN_11926; // @[decode.scala 512:28 657:39]
  wire [63:0] _GEN_11938 = _T_279 ? mtval : _GEN_11927; // @[decode.scala 513:28 657:39]
  wire [63:0] _GEN_11939 = _T_279 ? mip : _GEN_11928; // @[decode.scala 514:28 657:39]
  wire [63:0] _GEN_11940 = _T_279 ? pmpcfg0 : _GEN_11929; // @[decode.scala 515:28 657:39]
  wire [63:0] _GEN_11941 = _T_279 ? pmpaddr0 : _GEN_11930; // @[decode.scala 516:28 657:39]
  wire [63:0] _GEN_11942 = _T_279 ? mvendorid : _GEN_11931; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_11943 = _T_279 ? marchid : _GEN_11932; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_11944 = _T_279 ? mimpid : _GEN_11933; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_11945 = _T_279 ? mhartid : _GEN_11934; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_11946 = _T_278 ? csrImmReg : mcounteren; // @[decode.scala 509:28 657:39 670:38]
  wire [63:0] _GEN_11947 = _T_278 ? mscratch : _GEN_11935; // @[decode.scala 510:28 657:39]
  wire [63:0] _GEN_11948 = _T_278 ? mepc : _GEN_11936; // @[decode.scala 511:28 657:39]
  wire [63:0] _GEN_11949 = _T_278 ? mcause : _GEN_11937; // @[decode.scala 512:28 657:39]
  wire [63:0] _GEN_11950 = _T_278 ? mtval : _GEN_11938; // @[decode.scala 513:28 657:39]
  wire [63:0] _GEN_11951 = _T_278 ? mip : _GEN_11939; // @[decode.scala 514:28 657:39]
  wire [63:0] _GEN_11952 = _T_278 ? pmpcfg0 : _GEN_11940; // @[decode.scala 515:28 657:39]
  wire [63:0] _GEN_11953 = _T_278 ? pmpaddr0 : _GEN_11941; // @[decode.scala 516:28 657:39]
  wire [63:0] _GEN_11954 = _T_278 ? mvendorid : _GEN_11942; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_11955 = _T_278 ? marchid : _GEN_11943; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_11956 = _T_278 ? mimpid : _GEN_11944; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_11957 = _T_278 ? mhartid : _GEN_11945; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_11958 = _T_277 ? csrImmReg : mtvec; // @[decode.scala 508:28 657:39 669:38]
  wire [63:0] _GEN_11959 = _T_277 ? mcounteren : _GEN_11946; // @[decode.scala 509:28 657:39]
  wire [63:0] _GEN_11960 = _T_277 ? mscratch : _GEN_11947; // @[decode.scala 510:28 657:39]
  wire [63:0] _GEN_11961 = _T_277 ? mepc : _GEN_11948; // @[decode.scala 511:28 657:39]
  wire [63:0] _GEN_11962 = _T_277 ? mcause : _GEN_11949; // @[decode.scala 512:28 657:39]
  wire [63:0] _GEN_11963 = _T_277 ? mtval : _GEN_11950; // @[decode.scala 513:28 657:39]
  wire [63:0] _GEN_11964 = _T_277 ? mip : _GEN_11951; // @[decode.scala 514:28 657:39]
  wire [63:0] _GEN_11965 = _T_277 ? pmpcfg0 : _GEN_11952; // @[decode.scala 515:28 657:39]
  wire [63:0] _GEN_11966 = _T_277 ? pmpaddr0 : _GEN_11953; // @[decode.scala 516:28 657:39]
  wire [63:0] _GEN_11967 = _T_277 ? mvendorid : _GEN_11954; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_11968 = _T_277 ? marchid : _GEN_11955; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_11969 = _T_277 ? mimpid : _GEN_11956; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_11970 = _T_277 ? mhartid : _GEN_11957; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_11971 = _T_276 ? csrImmReg : mie; // @[decode.scala 507:28 657:39 668:38]
  wire [63:0] _GEN_11972 = _T_276 ? mtvec : _GEN_11958; // @[decode.scala 508:28 657:39]
  wire [63:0] _GEN_11973 = _T_276 ? mcounteren : _GEN_11959; // @[decode.scala 509:28 657:39]
  wire [63:0] _GEN_11974 = _T_276 ? mscratch : _GEN_11960; // @[decode.scala 510:28 657:39]
  wire [63:0] _GEN_11975 = _T_276 ? mepc : _GEN_11961; // @[decode.scala 511:28 657:39]
  wire [63:0] _GEN_11976 = _T_276 ? mcause : _GEN_11962; // @[decode.scala 512:28 657:39]
  wire [63:0] _GEN_11977 = _T_276 ? mtval : _GEN_11963; // @[decode.scala 513:28 657:39]
  wire [63:0] _GEN_11978 = _T_276 ? mip : _GEN_11964; // @[decode.scala 514:28 657:39]
  wire [63:0] _GEN_11979 = _T_276 ? pmpcfg0 : _GEN_11965; // @[decode.scala 515:28 657:39]
  wire [63:0] _GEN_11980 = _T_276 ? pmpaddr0 : _GEN_11966; // @[decode.scala 516:28 657:39]
  wire [63:0] _GEN_11981 = _T_276 ? mvendorid : _GEN_11967; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_11982 = _T_276 ? marchid : _GEN_11968; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_11983 = _T_276 ? mimpid : _GEN_11969; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_11984 = _T_276 ? mhartid : _GEN_11970; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_11985 = _T_275 ? csrImmReg : mideleg; // @[decode.scala 506:28 657:39 667:38]
  wire [63:0] _GEN_11986 = _T_275 ? mie : _GEN_11971; // @[decode.scala 507:28 657:39]
  wire [63:0] _GEN_11987 = _T_275 ? mtvec : _GEN_11972; // @[decode.scala 508:28 657:39]
  wire [63:0] _GEN_11988 = _T_275 ? mcounteren : _GEN_11973; // @[decode.scala 509:28 657:39]
  wire [63:0] _GEN_11989 = _T_275 ? mscratch : _GEN_11974; // @[decode.scala 510:28 657:39]
  wire [63:0] _GEN_11990 = _T_275 ? mepc : _GEN_11975; // @[decode.scala 511:28 657:39]
  wire [63:0] _GEN_11991 = _T_275 ? mcause : _GEN_11976; // @[decode.scala 512:28 657:39]
  wire [63:0] _GEN_11992 = _T_275 ? mtval : _GEN_11977; // @[decode.scala 513:28 657:39]
  wire [63:0] _GEN_11993 = _T_275 ? mip : _GEN_11978; // @[decode.scala 514:28 657:39]
  wire [63:0] _GEN_11994 = _T_275 ? pmpcfg0 : _GEN_11979; // @[decode.scala 515:28 657:39]
  wire [63:0] _GEN_11995 = _T_275 ? pmpaddr0 : _GEN_11980; // @[decode.scala 516:28 657:39]
  wire [63:0] _GEN_11996 = _T_275 ? mvendorid : _GEN_11981; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_11997 = _T_275 ? marchid : _GEN_11982; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_11998 = _T_275 ? mimpid : _GEN_11983; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_11999 = _T_275 ? mhartid : _GEN_11984; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_12000 = _T_274 ? csrImmReg : medeleg; // @[decode.scala 505:28 657:39 666:38]
  wire [63:0] _GEN_12001 = _T_274 ? mideleg : _GEN_11985; // @[decode.scala 506:28 657:39]
  wire [63:0] _GEN_12002 = _T_274 ? mie : _GEN_11986; // @[decode.scala 507:28 657:39]
  wire [63:0] _GEN_12003 = _T_274 ? mtvec : _GEN_11987; // @[decode.scala 508:28 657:39]
  wire [63:0] _GEN_12004 = _T_274 ? mcounteren : _GEN_11988; // @[decode.scala 509:28 657:39]
  wire [63:0] _GEN_12005 = _T_274 ? mscratch : _GEN_11989; // @[decode.scala 510:28 657:39]
  wire [63:0] _GEN_12006 = _T_274 ? mepc : _GEN_11990; // @[decode.scala 511:28 657:39]
  wire [63:0] _GEN_12007 = _T_274 ? mcause : _GEN_11991; // @[decode.scala 512:28 657:39]
  wire [63:0] _GEN_12008 = _T_274 ? mtval : _GEN_11992; // @[decode.scala 513:28 657:39]
  wire [63:0] _GEN_12009 = _T_274 ? mip : _GEN_11993; // @[decode.scala 514:28 657:39]
  wire [63:0] _GEN_12010 = _T_274 ? pmpcfg0 : _GEN_11994; // @[decode.scala 515:28 657:39]
  wire [63:0] _GEN_12011 = _T_274 ? pmpaddr0 : _GEN_11995; // @[decode.scala 516:28 657:39]
  wire [63:0] _GEN_12012 = _T_274 ? mvendorid : _GEN_11996; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_12013 = _T_274 ? marchid : _GEN_11997; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_12014 = _T_274 ? mimpid : _GEN_11998; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_12015 = _T_274 ? mhartid : _GEN_11999; // @[decode.scala 520:28 657:39]
  wire [126:0] _GEN_12016 = _T_273 ? {{63'd0}, csrImmReg} : 127'h8000000000101101; // @[decode.scala 657:39 665:38 523:8]
  wire [63:0] _GEN_12017 = _T_273 ? medeleg : _GEN_12000; // @[decode.scala 505:28 657:39]
  wire [63:0] _GEN_12018 = _T_273 ? mideleg : _GEN_12001; // @[decode.scala 506:28 657:39]
  wire [63:0] _GEN_12019 = _T_273 ? mie : _GEN_12002; // @[decode.scala 507:28 657:39]
  wire [63:0] _GEN_12020 = _T_273 ? mtvec : _GEN_12003; // @[decode.scala 508:28 657:39]
  wire [63:0] _GEN_12021 = _T_273 ? mcounteren : _GEN_12004; // @[decode.scala 509:28 657:39]
  wire [63:0] _GEN_12022 = _T_273 ? mscratch : _GEN_12005; // @[decode.scala 510:28 657:39]
  wire [63:0] _GEN_12023 = _T_273 ? mepc : _GEN_12006; // @[decode.scala 511:28 657:39]
  wire [63:0] _GEN_12024 = _T_273 ? mcause : _GEN_12007; // @[decode.scala 512:28 657:39]
  wire [63:0] _GEN_12025 = _T_273 ? mtval : _GEN_12008; // @[decode.scala 513:28 657:39]
  wire [63:0] _GEN_12026 = _T_273 ? mip : _GEN_12009; // @[decode.scala 514:28 657:39]
  wire [63:0] _GEN_12027 = _T_273 ? pmpcfg0 : _GEN_12010; // @[decode.scala 515:28 657:39]
  wire [63:0] _GEN_12028 = _T_273 ? pmpaddr0 : _GEN_12011; // @[decode.scala 516:28 657:39]
  wire [63:0] _GEN_12029 = _T_273 ? mvendorid : _GEN_12012; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_12030 = _T_273 ? marchid : _GEN_12013; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_12031 = _T_273 ? mimpid : _GEN_12014; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_12032 = _T_273 ? mhartid : _GEN_12015; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_12033 = _T_272 ? csrImmReg : _mstatus_T_1; // @[decode.scala 522:11 657:39 664:38]
  wire [126:0] _GEN_12034 = _T_272 ? 127'h8000000000101101 : _GEN_12016; // @[decode.scala 657:39 523:8]
  wire [63:0] _GEN_12035 = _T_272 ? medeleg : _GEN_12017; // @[decode.scala 505:28 657:39]
  wire [63:0] _GEN_12036 = _T_272 ? mideleg : _GEN_12018; // @[decode.scala 506:28 657:39]
  wire [63:0] _GEN_12037 = _T_272 ? mie : _GEN_12019; // @[decode.scala 507:28 657:39]
  wire [63:0] _GEN_12038 = _T_272 ? mtvec : _GEN_12020; // @[decode.scala 508:28 657:39]
  wire [63:0] _GEN_12039 = _T_272 ? mcounteren : _GEN_12021; // @[decode.scala 509:28 657:39]
  wire [63:0] _GEN_12040 = _T_272 ? mscratch : _GEN_12022; // @[decode.scala 510:28 657:39]
  wire [63:0] _GEN_12041 = _T_272 ? mepc : _GEN_12023; // @[decode.scala 511:28 657:39]
  wire [63:0] _GEN_12042 = _T_272 ? mcause : _GEN_12024; // @[decode.scala 512:28 657:39]
  wire [63:0] _GEN_12043 = _T_272 ? mtval : _GEN_12025; // @[decode.scala 513:28 657:39]
  wire [63:0] _GEN_12044 = _T_272 ? mip : _GEN_12026; // @[decode.scala 514:28 657:39]
  wire [63:0] _GEN_12045 = _T_272 ? pmpcfg0 : _GEN_12027; // @[decode.scala 515:28 657:39]
  wire [63:0] _GEN_12046 = _T_272 ? pmpaddr0 : _GEN_12028; // @[decode.scala 516:28 657:39]
  wire [63:0] _GEN_12047 = _T_272 ? mvendorid : _GEN_12029; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_12048 = _T_272 ? marchid : _GEN_12030; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_12049 = _T_272 ? mimpid : _GEN_12031; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_12050 = _T_272 ? mhartid : _GEN_12032; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_12051 = _T_271 ? csrImmReg : satp; // @[decode.scala 502:28 657:39 663:38]
  wire [63:0] _GEN_12052 = _T_271 ? _mstatus_T_1 : _GEN_12033; // @[decode.scala 522:11 657:39]
  wire [126:0] _GEN_12053 = _T_271 ? 127'h8000000000101101 : _GEN_12034; // @[decode.scala 657:39 523:8]
  wire [63:0] _GEN_12054 = _T_271 ? medeleg : _GEN_12035; // @[decode.scala 505:28 657:39]
  wire [63:0] _GEN_12055 = _T_271 ? mideleg : _GEN_12036; // @[decode.scala 506:28 657:39]
  wire [63:0] _GEN_12056 = _T_271 ? mie : _GEN_12037; // @[decode.scala 507:28 657:39]
  wire [63:0] _GEN_12057 = _T_271 ? mtvec : _GEN_12038; // @[decode.scala 508:28 657:39]
  wire [63:0] _GEN_12058 = _T_271 ? mcounteren : _GEN_12039; // @[decode.scala 509:28 657:39]
  wire [63:0] _GEN_12059 = _T_271 ? mscratch : _GEN_12040; // @[decode.scala 510:28 657:39]
  wire [63:0] _GEN_12060 = _T_271 ? mepc : _GEN_12041; // @[decode.scala 511:28 657:39]
  wire [63:0] _GEN_12061 = _T_271 ? mcause : _GEN_12042; // @[decode.scala 512:28 657:39]
  wire [63:0] _GEN_12062 = _T_271 ? mtval : _GEN_12043; // @[decode.scala 513:28 657:39]
  wire [63:0] _GEN_12063 = _T_271 ? mip : _GEN_12044; // @[decode.scala 514:28 657:39]
  wire [63:0] _GEN_12064 = _T_271 ? pmpcfg0 : _GEN_12045; // @[decode.scala 515:28 657:39]
  wire [63:0] _GEN_12065 = _T_271 ? pmpaddr0 : _GEN_12046; // @[decode.scala 516:28 657:39]
  wire [63:0] _GEN_12066 = _T_271 ? mvendorid : _GEN_12047; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_12067 = _T_271 ? marchid : _GEN_12048; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_12068 = _T_271 ? mimpid : _GEN_12049; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_12069 = _T_271 ? mhartid : _GEN_12050; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_12070 = _T_270 ? csrImmReg : scounteren; // @[decode.scala 501:28 657:39 662:38]
  wire [63:0] _GEN_12071 = _T_270 ? satp : _GEN_12051; // @[decode.scala 502:28 657:39]
  wire [63:0] _GEN_12072 = _T_270 ? _mstatus_T_1 : _GEN_12052; // @[decode.scala 522:11 657:39]
  wire [126:0] _GEN_12073 = _T_270 ? 127'h8000000000101101 : _GEN_12053; // @[decode.scala 657:39 523:8]
  wire [63:0] _GEN_12074 = _T_270 ? medeleg : _GEN_12054; // @[decode.scala 505:28 657:39]
  wire [63:0] _GEN_12075 = _T_270 ? mideleg : _GEN_12055; // @[decode.scala 506:28 657:39]
  wire [63:0] _GEN_12076 = _T_270 ? mie : _GEN_12056; // @[decode.scala 507:28 657:39]
  wire [63:0] _GEN_12077 = _T_270 ? mtvec : _GEN_12057; // @[decode.scala 508:28 657:39]
  wire [63:0] _GEN_12078 = _T_270 ? mcounteren : _GEN_12058; // @[decode.scala 509:28 657:39]
  wire [63:0] _GEN_12079 = _T_270 ? mscratch : _GEN_12059; // @[decode.scala 510:28 657:39]
  wire [63:0] _GEN_12080 = _T_270 ? mepc : _GEN_12060; // @[decode.scala 511:28 657:39]
  wire [63:0] _GEN_12081 = _T_270 ? mcause : _GEN_12061; // @[decode.scala 512:28 657:39]
  wire [63:0] _GEN_12082 = _T_270 ? mtval : _GEN_12062; // @[decode.scala 513:28 657:39]
  wire [63:0] _GEN_12083 = _T_270 ? mip : _GEN_12063; // @[decode.scala 514:28 657:39]
  wire [63:0] _GEN_12084 = _T_270 ? pmpcfg0 : _GEN_12064; // @[decode.scala 515:28 657:39]
  wire [63:0] _GEN_12085 = _T_270 ? pmpaddr0 : _GEN_12065; // @[decode.scala 516:28 657:39]
  wire [63:0] _GEN_12086 = _T_270 ? mvendorid : _GEN_12066; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_12087 = _T_270 ? marchid : _GEN_12067; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_12088 = _T_270 ? mimpid : _GEN_12068; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_12089 = _T_270 ? mhartid : _GEN_12069; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_12090 = _T_269 ? csrImmReg : ucause; // @[decode.scala 500:28 657:39 661:38]
  wire [63:0] _GEN_12091 = _T_269 ? scounteren : _GEN_12070; // @[decode.scala 501:28 657:39]
  wire [63:0] _GEN_12092 = _T_269 ? satp : _GEN_12071; // @[decode.scala 502:28 657:39]
  wire [63:0] _GEN_12093 = _T_269 ? _mstatus_T_1 : _GEN_12072; // @[decode.scala 522:11 657:39]
  wire [126:0] _GEN_12094 = _T_269 ? 127'h8000000000101101 : _GEN_12073; // @[decode.scala 657:39 523:8]
  wire [63:0] _GEN_12095 = _T_269 ? medeleg : _GEN_12074; // @[decode.scala 505:28 657:39]
  wire [63:0] _GEN_12096 = _T_269 ? mideleg : _GEN_12075; // @[decode.scala 506:28 657:39]
  wire [63:0] _GEN_12097 = _T_269 ? mie : _GEN_12076; // @[decode.scala 507:28 657:39]
  wire [63:0] _GEN_12098 = _T_269 ? mtvec : _GEN_12077; // @[decode.scala 508:28 657:39]
  wire [63:0] _GEN_12099 = _T_269 ? mcounteren : _GEN_12078; // @[decode.scala 509:28 657:39]
  wire [63:0] _GEN_12100 = _T_269 ? mscratch : _GEN_12079; // @[decode.scala 510:28 657:39]
  wire [63:0] _GEN_12101 = _T_269 ? mepc : _GEN_12080; // @[decode.scala 511:28 657:39]
  wire [63:0] _GEN_12102 = _T_269 ? mcause : _GEN_12081; // @[decode.scala 512:28 657:39]
  wire [63:0] _GEN_12103 = _T_269 ? mtval : _GEN_12082; // @[decode.scala 513:28 657:39]
  wire [63:0] _GEN_12104 = _T_269 ? mip : _GEN_12083; // @[decode.scala 514:28 657:39]
  wire [63:0] _GEN_12105 = _T_269 ? pmpcfg0 : _GEN_12084; // @[decode.scala 515:28 657:39]
  wire [63:0] _GEN_12106 = _T_269 ? pmpaddr0 : _GEN_12085; // @[decode.scala 516:28 657:39]
  wire [63:0] _GEN_12107 = _T_269 ? mvendorid : _GEN_12086; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_12108 = _T_269 ? marchid : _GEN_12087; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_12109 = _T_269 ? mimpid : _GEN_12088; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_12110 = _T_269 ? mhartid : _GEN_12089; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_12111 = _T_268 ? csrImmReg : uepc; // @[decode.scala 499:28 657:39 660:38]
  wire [63:0] _GEN_12112 = _T_268 ? ucause : _GEN_12090; // @[decode.scala 500:28 657:39]
  wire [63:0] _GEN_12113 = _T_268 ? scounteren : _GEN_12091; // @[decode.scala 501:28 657:39]
  wire [63:0] _GEN_12114 = _T_268 ? satp : _GEN_12092; // @[decode.scala 502:28 657:39]
  wire [63:0] _GEN_12115 = _T_268 ? _mstatus_T_1 : _GEN_12093; // @[decode.scala 522:11 657:39]
  wire [126:0] _GEN_12116 = _T_268 ? 127'h8000000000101101 : _GEN_12094; // @[decode.scala 657:39 523:8]
  wire [63:0] _GEN_12117 = _T_268 ? medeleg : _GEN_12095; // @[decode.scala 505:28 657:39]
  wire [63:0] _GEN_12118 = _T_268 ? mideleg : _GEN_12096; // @[decode.scala 506:28 657:39]
  wire [63:0] _GEN_12119 = _T_268 ? mie : _GEN_12097; // @[decode.scala 507:28 657:39]
  wire [63:0] _GEN_12120 = _T_268 ? mtvec : _GEN_12098; // @[decode.scala 508:28 657:39]
  wire [63:0] _GEN_12121 = _T_268 ? mcounteren : _GEN_12099; // @[decode.scala 509:28 657:39]
  wire [63:0] _GEN_12122 = _T_268 ? mscratch : _GEN_12100; // @[decode.scala 510:28 657:39]
  wire [63:0] _GEN_12123 = _T_268 ? mepc : _GEN_12101; // @[decode.scala 511:28 657:39]
  wire [63:0] _GEN_12124 = _T_268 ? mcause : _GEN_12102; // @[decode.scala 512:28 657:39]
  wire [63:0] _GEN_12125 = _T_268 ? mtval : _GEN_12103; // @[decode.scala 513:28 657:39]
  wire [63:0] _GEN_12126 = _T_268 ? mip : _GEN_12104; // @[decode.scala 514:28 657:39]
  wire [63:0] _GEN_12127 = _T_268 ? pmpcfg0 : _GEN_12105; // @[decode.scala 515:28 657:39]
  wire [63:0] _GEN_12128 = _T_268 ? pmpaddr0 : _GEN_12106; // @[decode.scala 516:28 657:39]
  wire [63:0] _GEN_12129 = _T_268 ? mvendorid : _GEN_12107; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_12130 = _T_268 ? marchid : _GEN_12108; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_12131 = _T_268 ? mimpid : _GEN_12109; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_12132 = _T_268 ? mhartid : _GEN_12110; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_12133 = _T_267 ? csrImmReg : utvec; // @[decode.scala 498:28 657:39 659:38]
  wire [63:0] _GEN_12134 = _T_267 ? uepc : _GEN_12111; // @[decode.scala 499:28 657:39]
  wire [63:0] _GEN_12135 = _T_267 ? ucause : _GEN_12112; // @[decode.scala 500:28 657:39]
  wire [63:0] _GEN_12136 = _T_267 ? scounteren : _GEN_12113; // @[decode.scala 501:28 657:39]
  wire [63:0] _GEN_12137 = _T_267 ? satp : _GEN_12114; // @[decode.scala 502:28 657:39]
  wire [63:0] _GEN_12138 = _T_267 ? _mstatus_T_1 : _GEN_12115; // @[decode.scala 522:11 657:39]
  wire [126:0] _GEN_12139 = _T_267 ? 127'h8000000000101101 : _GEN_12116; // @[decode.scala 657:39 523:8]
  wire [63:0] _GEN_12140 = _T_267 ? medeleg : _GEN_12117; // @[decode.scala 505:28 657:39]
  wire [63:0] _GEN_12141 = _T_267 ? mideleg : _GEN_12118; // @[decode.scala 506:28 657:39]
  wire [63:0] _GEN_12142 = _T_267 ? mie : _GEN_12119; // @[decode.scala 507:28 657:39]
  wire [63:0] _GEN_12143 = _T_267 ? mtvec : _GEN_12120; // @[decode.scala 508:28 657:39]
  wire [63:0] _GEN_12144 = _T_267 ? mcounteren : _GEN_12121; // @[decode.scala 509:28 657:39]
  wire [63:0] _GEN_12145 = _T_267 ? mscratch : _GEN_12122; // @[decode.scala 510:28 657:39]
  wire [63:0] _GEN_12146 = _T_267 ? mepc : _GEN_12123; // @[decode.scala 511:28 657:39]
  wire [63:0] _GEN_12147 = _T_267 ? mcause : _GEN_12124; // @[decode.scala 512:28 657:39]
  wire [63:0] _GEN_12148 = _T_267 ? mtval : _GEN_12125; // @[decode.scala 513:28 657:39]
  wire [63:0] _GEN_12149 = _T_267 ? mip : _GEN_12126; // @[decode.scala 514:28 657:39]
  wire [63:0] _GEN_12150 = _T_267 ? pmpcfg0 : _GEN_12127; // @[decode.scala 515:28 657:39]
  wire [63:0] _GEN_12151 = _T_267 ? pmpaddr0 : _GEN_12128; // @[decode.scala 516:28 657:39]
  wire [63:0] _GEN_12152 = _T_267 ? mvendorid : _GEN_12129; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_12153 = _T_267 ? marchid : _GEN_12130; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_12154 = _T_267 ? mimpid : _GEN_12131; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_12155 = _T_267 ? mhartid : _GEN_12132; // @[decode.scala 520:28 657:39]
  wire [63:0] _GEN_12156 = _T_266 ? csrImmReg : ustatus; // @[decode.scala 497:28 657:39 658:38]
  wire [63:0] _GEN_12157 = _T_266 ? utvec : _GEN_12133; // @[decode.scala 498:28 657:39]
  wire [63:0] _GEN_12158 = _T_266 ? uepc : _GEN_12134; // @[decode.scala 499:28 657:39]
  wire [63:0] _GEN_12159 = _T_266 ? ucause : _GEN_12135; // @[decode.scala 500:28 657:39]
  wire [63:0] _GEN_12160 = _T_266 ? scounteren : _GEN_12136; // @[decode.scala 501:28 657:39]
  wire [63:0] _GEN_12161 = _T_266 ? satp : _GEN_12137; // @[decode.scala 502:28 657:39]
  wire [63:0] _GEN_12162 = _T_266 ? _mstatus_T_1 : _GEN_12138; // @[decode.scala 522:11 657:39]
  wire [126:0] _GEN_12163 = _T_266 ? 127'h8000000000101101 : _GEN_12139; // @[decode.scala 657:39 523:8]
  wire [63:0] _GEN_12164 = _T_266 ? medeleg : _GEN_12140; // @[decode.scala 505:28 657:39]
  wire [63:0] _GEN_12165 = _T_266 ? mideleg : _GEN_12141; // @[decode.scala 506:28 657:39]
  wire [63:0] _GEN_12166 = _T_266 ? mie : _GEN_12142; // @[decode.scala 507:28 657:39]
  wire [63:0] _GEN_12167 = _T_266 ? mtvec : _GEN_12143; // @[decode.scala 508:28 657:39]
  wire [63:0] _GEN_12168 = _T_266 ? mcounteren : _GEN_12144; // @[decode.scala 509:28 657:39]
  wire [63:0] _GEN_12169 = _T_266 ? mscratch : _GEN_12145; // @[decode.scala 510:28 657:39]
  wire [63:0] _GEN_12170 = _T_266 ? mepc : _GEN_12146; // @[decode.scala 511:28 657:39]
  wire [63:0] _GEN_12171 = _T_266 ? mcause : _GEN_12147; // @[decode.scala 512:28 657:39]
  wire [63:0] _GEN_12172 = _T_266 ? mtval : _GEN_12148; // @[decode.scala 513:28 657:39]
  wire [63:0] _GEN_12173 = _T_266 ? mip : _GEN_12149; // @[decode.scala 514:28 657:39]
  wire [63:0] _GEN_12174 = _T_266 ? pmpcfg0 : _GEN_12150; // @[decode.scala 515:28 657:39]
  wire [63:0] _GEN_12175 = _T_266 ? pmpaddr0 : _GEN_12151; // @[decode.scala 516:28 657:39]
  wire [63:0] _GEN_12176 = _T_266 ? mvendorid : _GEN_12152; // @[decode.scala 517:28 657:39]
  wire [63:0] _GEN_12177 = _T_266 ? marchid : _GEN_12153; // @[decode.scala 518:28 657:39]
  wire [63:0] _GEN_12178 = _T_266 ? mimpid : _GEN_12154; // @[decode.scala 519:28 657:39]
  wire [63:0] _GEN_12179 = _T_266 ? mhartid : _GEN_12155; // @[decode.scala 520:28 657:39]
  wire [63:0] _ustatus_T_3 = ustatus | csrImmReg; // @[decode.scala 686:49]
  wire [63:0] _utvec_T_3 = utvec | csrImmReg; // @[decode.scala 687:47]
  wire [63:0] _uepc_T_3 = uepc | csrImmReg; // @[decode.scala 688:46]
  wire [63:0] _ucause_T_3 = ucause | csrImmReg; // @[decode.scala 689:48]
  wire [63:0] _scounteren_T_3 = scounteren | csrImmReg; // @[decode.scala 690:52]
  wire [63:0] _satp_T_3 = satp | csrImmReg; // @[decode.scala 691:46]
  wire [63:0] _mstatus_T_5 = mstatus | csrImmReg; // @[decode.scala 692:49]
  wire [63:0] _misa_T_5 = misa | csrImmReg; // @[decode.scala 693:46]
  wire [63:0] _medeleg_T_3 = medeleg | csrImmReg; // @[decode.scala 694:49]
  wire [63:0] _mideleg_T_3 = mideleg | csrImmReg; // @[decode.scala 695:49]
  wire [63:0] _mie_T_3 = mie | csrImmReg; // @[decode.scala 696:45]
  wire [63:0] _mtvec_T_3 = mtvec | csrImmReg; // @[decode.scala 697:47]
  wire [63:0] _mcounteren_T_3 = mcounteren | csrImmReg; // @[decode.scala 698:52]
  wire [63:0] _mscratch_T_3 = mscratch | csrImmReg; // @[decode.scala 699:50]
  wire [63:0] _mepc_T_3 = mepc | csrImmReg; // @[decode.scala 700:46]
  wire [63:0] _mcause_T_3 = mcause | csrImmReg; // @[decode.scala 701:48]
  wire [63:0] _mtval_T_3 = mtval | csrImmReg; // @[decode.scala 702:47]
  wire [63:0] _mip_T_3 = mip | csrImmReg; // @[decode.scala 703:45]
  wire [63:0] _pmpcfg0_T_3 = pmpcfg0 | csrImmReg; // @[decode.scala 704:49]
  wire [63:0] _pmpaddr0_T_3 = pmpaddr0 | csrImmReg; // @[decode.scala 705:50]
  wire [63:0] _mvendorid_T_3 = mvendorid | csrImmReg; // @[decode.scala 706:51]
  wire [63:0] _marchid_T_3 = marchid | csrImmReg; // @[decode.scala 707:49]
  wire [63:0] _mimpid_T_3 = mimpid | csrImmReg; // @[decode.scala 708:48]
  wire [63:0] _mhartid_T_3 = mhartid | csrImmReg; // @[decode.scala 709:49]
  wire [63:0] _GEN_12180 = _T_289 ? _mhartid_T_3 : mhartid; // @[decode.scala 520:28 685:39 709:38]
  wire [63:0] _GEN_12181 = _T_288 ? _mimpid_T_3 : mimpid; // @[decode.scala 519:28 685:39 708:38]
  wire [63:0] _GEN_12182 = _T_288 ? mhartid : _GEN_12180; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12183 = _T_287 ? _marchid_T_3 : marchid; // @[decode.scala 518:28 685:39 707:38]
  wire [63:0] _GEN_12184 = _T_287 ? mimpid : _GEN_12181; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12185 = _T_287 ? mhartid : _GEN_12182; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12186 = _T_286 ? _mvendorid_T_3 : mvendorid; // @[decode.scala 517:28 685:39 706:38]
  wire [63:0] _GEN_12187 = _T_286 ? marchid : _GEN_12183; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12188 = _T_286 ? mimpid : _GEN_12184; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12189 = _T_286 ? mhartid : _GEN_12185; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12190 = _T_285 ? _pmpaddr0_T_3 : pmpaddr0; // @[decode.scala 516:28 685:39 705:38]
  wire [63:0] _GEN_12191 = _T_285 ? mvendorid : _GEN_12186; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12192 = _T_285 ? marchid : _GEN_12187; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12193 = _T_285 ? mimpid : _GEN_12188; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12194 = _T_285 ? mhartid : _GEN_12189; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12195 = _T_284 ? _pmpcfg0_T_3 : pmpcfg0; // @[decode.scala 515:28 685:39 704:38]
  wire [63:0] _GEN_12196 = _T_284 ? pmpaddr0 : _GEN_12190; // @[decode.scala 516:28 685:39]
  wire [63:0] _GEN_12197 = _T_284 ? mvendorid : _GEN_12191; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12198 = _T_284 ? marchid : _GEN_12192; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12199 = _T_284 ? mimpid : _GEN_12193; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12200 = _T_284 ? mhartid : _GEN_12194; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12201 = _T_283 ? _mip_T_3 : mip; // @[decode.scala 514:28 685:39 703:38]
  wire [63:0] _GEN_12202 = _T_283 ? pmpcfg0 : _GEN_12195; // @[decode.scala 515:28 685:39]
  wire [63:0] _GEN_12203 = _T_283 ? pmpaddr0 : _GEN_12196; // @[decode.scala 516:28 685:39]
  wire [63:0] _GEN_12204 = _T_283 ? mvendorid : _GEN_12197; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12205 = _T_283 ? marchid : _GEN_12198; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12206 = _T_283 ? mimpid : _GEN_12199; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12207 = _T_283 ? mhartid : _GEN_12200; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12208 = _T_282 ? _mtval_T_3 : mtval; // @[decode.scala 513:28 685:39 702:38]
  wire [63:0] _GEN_12209 = _T_282 ? mip : _GEN_12201; // @[decode.scala 514:28 685:39]
  wire [63:0] _GEN_12210 = _T_282 ? pmpcfg0 : _GEN_12202; // @[decode.scala 515:28 685:39]
  wire [63:0] _GEN_12211 = _T_282 ? pmpaddr0 : _GEN_12203; // @[decode.scala 516:28 685:39]
  wire [63:0] _GEN_12212 = _T_282 ? mvendorid : _GEN_12204; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12213 = _T_282 ? marchid : _GEN_12205; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12214 = _T_282 ? mimpid : _GEN_12206; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12215 = _T_282 ? mhartid : _GEN_12207; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12216 = _T_281 ? _mcause_T_3 : mcause; // @[decode.scala 512:28 685:39 701:38]
  wire [63:0] _GEN_12217 = _T_281 ? mtval : _GEN_12208; // @[decode.scala 513:28 685:39]
  wire [63:0] _GEN_12218 = _T_281 ? mip : _GEN_12209; // @[decode.scala 514:28 685:39]
  wire [63:0] _GEN_12219 = _T_281 ? pmpcfg0 : _GEN_12210; // @[decode.scala 515:28 685:39]
  wire [63:0] _GEN_12220 = _T_281 ? pmpaddr0 : _GEN_12211; // @[decode.scala 516:28 685:39]
  wire [63:0] _GEN_12221 = _T_281 ? mvendorid : _GEN_12212; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12222 = _T_281 ? marchid : _GEN_12213; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12223 = _T_281 ? mimpid : _GEN_12214; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12224 = _T_281 ? mhartid : _GEN_12215; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12225 = _T_280 ? _mepc_T_3 : mepc; // @[decode.scala 511:28 685:39 700:38]
  wire [63:0] _GEN_12226 = _T_280 ? mcause : _GEN_12216; // @[decode.scala 512:28 685:39]
  wire [63:0] _GEN_12227 = _T_280 ? mtval : _GEN_12217; // @[decode.scala 513:28 685:39]
  wire [63:0] _GEN_12228 = _T_280 ? mip : _GEN_12218; // @[decode.scala 514:28 685:39]
  wire [63:0] _GEN_12229 = _T_280 ? pmpcfg0 : _GEN_12219; // @[decode.scala 515:28 685:39]
  wire [63:0] _GEN_12230 = _T_280 ? pmpaddr0 : _GEN_12220; // @[decode.scala 516:28 685:39]
  wire [63:0] _GEN_12231 = _T_280 ? mvendorid : _GEN_12221; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12232 = _T_280 ? marchid : _GEN_12222; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12233 = _T_280 ? mimpid : _GEN_12223; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12234 = _T_280 ? mhartid : _GEN_12224; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12235 = _T_279 ? _mscratch_T_3 : mscratch; // @[decode.scala 510:28 685:39 699:38]
  wire [63:0] _GEN_12236 = _T_279 ? mepc : _GEN_12225; // @[decode.scala 511:28 685:39]
  wire [63:0] _GEN_12237 = _T_279 ? mcause : _GEN_12226; // @[decode.scala 512:28 685:39]
  wire [63:0] _GEN_12238 = _T_279 ? mtval : _GEN_12227; // @[decode.scala 513:28 685:39]
  wire [63:0] _GEN_12239 = _T_279 ? mip : _GEN_12228; // @[decode.scala 514:28 685:39]
  wire [63:0] _GEN_12240 = _T_279 ? pmpcfg0 : _GEN_12229; // @[decode.scala 515:28 685:39]
  wire [63:0] _GEN_12241 = _T_279 ? pmpaddr0 : _GEN_12230; // @[decode.scala 516:28 685:39]
  wire [63:0] _GEN_12242 = _T_279 ? mvendorid : _GEN_12231; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12243 = _T_279 ? marchid : _GEN_12232; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12244 = _T_279 ? mimpid : _GEN_12233; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12245 = _T_279 ? mhartid : _GEN_12234; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12246 = _T_278 ? _mcounteren_T_3 : mcounteren; // @[decode.scala 509:28 685:39 698:38]
  wire [63:0] _GEN_12247 = _T_278 ? mscratch : _GEN_12235; // @[decode.scala 510:28 685:39]
  wire [63:0] _GEN_12248 = _T_278 ? mepc : _GEN_12236; // @[decode.scala 511:28 685:39]
  wire [63:0] _GEN_12249 = _T_278 ? mcause : _GEN_12237; // @[decode.scala 512:28 685:39]
  wire [63:0] _GEN_12250 = _T_278 ? mtval : _GEN_12238; // @[decode.scala 513:28 685:39]
  wire [63:0] _GEN_12251 = _T_278 ? mip : _GEN_12239; // @[decode.scala 514:28 685:39]
  wire [63:0] _GEN_12252 = _T_278 ? pmpcfg0 : _GEN_12240; // @[decode.scala 515:28 685:39]
  wire [63:0] _GEN_12253 = _T_278 ? pmpaddr0 : _GEN_12241; // @[decode.scala 516:28 685:39]
  wire [63:0] _GEN_12254 = _T_278 ? mvendorid : _GEN_12242; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12255 = _T_278 ? marchid : _GEN_12243; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12256 = _T_278 ? mimpid : _GEN_12244; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12257 = _T_278 ? mhartid : _GEN_12245; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12258 = _T_277 ? _mtvec_T_3 : mtvec; // @[decode.scala 508:28 685:39 697:38]
  wire [63:0] _GEN_12259 = _T_277 ? mcounteren : _GEN_12246; // @[decode.scala 509:28 685:39]
  wire [63:0] _GEN_12260 = _T_277 ? mscratch : _GEN_12247; // @[decode.scala 510:28 685:39]
  wire [63:0] _GEN_12261 = _T_277 ? mepc : _GEN_12248; // @[decode.scala 511:28 685:39]
  wire [63:0] _GEN_12262 = _T_277 ? mcause : _GEN_12249; // @[decode.scala 512:28 685:39]
  wire [63:0] _GEN_12263 = _T_277 ? mtval : _GEN_12250; // @[decode.scala 513:28 685:39]
  wire [63:0] _GEN_12264 = _T_277 ? mip : _GEN_12251; // @[decode.scala 514:28 685:39]
  wire [63:0] _GEN_12265 = _T_277 ? pmpcfg0 : _GEN_12252; // @[decode.scala 515:28 685:39]
  wire [63:0] _GEN_12266 = _T_277 ? pmpaddr0 : _GEN_12253; // @[decode.scala 516:28 685:39]
  wire [63:0] _GEN_12267 = _T_277 ? mvendorid : _GEN_12254; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12268 = _T_277 ? marchid : _GEN_12255; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12269 = _T_277 ? mimpid : _GEN_12256; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12270 = _T_277 ? mhartid : _GEN_12257; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12271 = _T_276 ? _mie_T_3 : mie; // @[decode.scala 507:28 685:39 696:38]
  wire [63:0] _GEN_12272 = _T_276 ? mtvec : _GEN_12258; // @[decode.scala 508:28 685:39]
  wire [63:0] _GEN_12273 = _T_276 ? mcounteren : _GEN_12259; // @[decode.scala 509:28 685:39]
  wire [63:0] _GEN_12274 = _T_276 ? mscratch : _GEN_12260; // @[decode.scala 510:28 685:39]
  wire [63:0] _GEN_12275 = _T_276 ? mepc : _GEN_12261; // @[decode.scala 511:28 685:39]
  wire [63:0] _GEN_12276 = _T_276 ? mcause : _GEN_12262; // @[decode.scala 512:28 685:39]
  wire [63:0] _GEN_12277 = _T_276 ? mtval : _GEN_12263; // @[decode.scala 513:28 685:39]
  wire [63:0] _GEN_12278 = _T_276 ? mip : _GEN_12264; // @[decode.scala 514:28 685:39]
  wire [63:0] _GEN_12279 = _T_276 ? pmpcfg0 : _GEN_12265; // @[decode.scala 515:28 685:39]
  wire [63:0] _GEN_12280 = _T_276 ? pmpaddr0 : _GEN_12266; // @[decode.scala 516:28 685:39]
  wire [63:0] _GEN_12281 = _T_276 ? mvendorid : _GEN_12267; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12282 = _T_276 ? marchid : _GEN_12268; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12283 = _T_276 ? mimpid : _GEN_12269; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12284 = _T_276 ? mhartid : _GEN_12270; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12285 = _T_275 ? _mideleg_T_3 : mideleg; // @[decode.scala 506:28 685:39 695:38]
  wire [63:0] _GEN_12286 = _T_275 ? mie : _GEN_12271; // @[decode.scala 507:28 685:39]
  wire [63:0] _GEN_12287 = _T_275 ? mtvec : _GEN_12272; // @[decode.scala 508:28 685:39]
  wire [63:0] _GEN_12288 = _T_275 ? mcounteren : _GEN_12273; // @[decode.scala 509:28 685:39]
  wire [63:0] _GEN_12289 = _T_275 ? mscratch : _GEN_12274; // @[decode.scala 510:28 685:39]
  wire [63:0] _GEN_12290 = _T_275 ? mepc : _GEN_12275; // @[decode.scala 511:28 685:39]
  wire [63:0] _GEN_12291 = _T_275 ? mcause : _GEN_12276; // @[decode.scala 512:28 685:39]
  wire [63:0] _GEN_12292 = _T_275 ? mtval : _GEN_12277; // @[decode.scala 513:28 685:39]
  wire [63:0] _GEN_12293 = _T_275 ? mip : _GEN_12278; // @[decode.scala 514:28 685:39]
  wire [63:0] _GEN_12294 = _T_275 ? pmpcfg0 : _GEN_12279; // @[decode.scala 515:28 685:39]
  wire [63:0] _GEN_12295 = _T_275 ? pmpaddr0 : _GEN_12280; // @[decode.scala 516:28 685:39]
  wire [63:0] _GEN_12296 = _T_275 ? mvendorid : _GEN_12281; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12297 = _T_275 ? marchid : _GEN_12282; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12298 = _T_275 ? mimpid : _GEN_12283; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12299 = _T_275 ? mhartid : _GEN_12284; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12300 = _T_274 ? _medeleg_T_3 : medeleg; // @[decode.scala 505:28 685:39 694:38]
  wire [63:0] _GEN_12301 = _T_274 ? mideleg : _GEN_12285; // @[decode.scala 506:28 685:39]
  wire [63:0] _GEN_12302 = _T_274 ? mie : _GEN_12286; // @[decode.scala 507:28 685:39]
  wire [63:0] _GEN_12303 = _T_274 ? mtvec : _GEN_12287; // @[decode.scala 508:28 685:39]
  wire [63:0] _GEN_12304 = _T_274 ? mcounteren : _GEN_12288; // @[decode.scala 509:28 685:39]
  wire [63:0] _GEN_12305 = _T_274 ? mscratch : _GEN_12289; // @[decode.scala 510:28 685:39]
  wire [63:0] _GEN_12306 = _T_274 ? mepc : _GEN_12290; // @[decode.scala 511:28 685:39]
  wire [63:0] _GEN_12307 = _T_274 ? mcause : _GEN_12291; // @[decode.scala 512:28 685:39]
  wire [63:0] _GEN_12308 = _T_274 ? mtval : _GEN_12292; // @[decode.scala 513:28 685:39]
  wire [63:0] _GEN_12309 = _T_274 ? mip : _GEN_12293; // @[decode.scala 514:28 685:39]
  wire [63:0] _GEN_12310 = _T_274 ? pmpcfg0 : _GEN_12294; // @[decode.scala 515:28 685:39]
  wire [63:0] _GEN_12311 = _T_274 ? pmpaddr0 : _GEN_12295; // @[decode.scala 516:28 685:39]
  wire [63:0] _GEN_12312 = _T_274 ? mvendorid : _GEN_12296; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12313 = _T_274 ? marchid : _GEN_12297; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12314 = _T_274 ? mimpid : _GEN_12298; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12315 = _T_274 ? mhartid : _GEN_12299; // @[decode.scala 520:28 685:39]
  wire [126:0] _GEN_12316 = _T_273 ? {{63'd0}, _misa_T_5} : 127'h8000000000101101; // @[decode.scala 685:39 693:38 523:8]
  wire [63:0] _GEN_12317 = _T_273 ? medeleg : _GEN_12300; // @[decode.scala 505:28 685:39]
  wire [63:0] _GEN_12318 = _T_273 ? mideleg : _GEN_12301; // @[decode.scala 506:28 685:39]
  wire [63:0] _GEN_12319 = _T_273 ? mie : _GEN_12302; // @[decode.scala 507:28 685:39]
  wire [63:0] _GEN_12320 = _T_273 ? mtvec : _GEN_12303; // @[decode.scala 508:28 685:39]
  wire [63:0] _GEN_12321 = _T_273 ? mcounteren : _GEN_12304; // @[decode.scala 509:28 685:39]
  wire [63:0] _GEN_12322 = _T_273 ? mscratch : _GEN_12305; // @[decode.scala 510:28 685:39]
  wire [63:0] _GEN_12323 = _T_273 ? mepc : _GEN_12306; // @[decode.scala 511:28 685:39]
  wire [63:0] _GEN_12324 = _T_273 ? mcause : _GEN_12307; // @[decode.scala 512:28 685:39]
  wire [63:0] _GEN_12325 = _T_273 ? mtval : _GEN_12308; // @[decode.scala 513:28 685:39]
  wire [63:0] _GEN_12326 = _T_273 ? mip : _GEN_12309; // @[decode.scala 514:28 685:39]
  wire [63:0] _GEN_12327 = _T_273 ? pmpcfg0 : _GEN_12310; // @[decode.scala 515:28 685:39]
  wire [63:0] _GEN_12328 = _T_273 ? pmpaddr0 : _GEN_12311; // @[decode.scala 516:28 685:39]
  wire [63:0] _GEN_12329 = _T_273 ? mvendorid : _GEN_12312; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12330 = _T_273 ? marchid : _GEN_12313; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12331 = _T_273 ? mimpid : _GEN_12314; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12332 = _T_273 ? mhartid : _GEN_12315; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12333 = _T_272 ? _mstatus_T_5 : _mstatus_T_1; // @[decode.scala 522:11 685:39 692:38]
  wire [126:0] _GEN_12334 = _T_272 ? 127'h8000000000101101 : _GEN_12316; // @[decode.scala 685:39 523:8]
  wire [63:0] _GEN_12335 = _T_272 ? medeleg : _GEN_12317; // @[decode.scala 505:28 685:39]
  wire [63:0] _GEN_12336 = _T_272 ? mideleg : _GEN_12318; // @[decode.scala 506:28 685:39]
  wire [63:0] _GEN_12337 = _T_272 ? mie : _GEN_12319; // @[decode.scala 507:28 685:39]
  wire [63:0] _GEN_12338 = _T_272 ? mtvec : _GEN_12320; // @[decode.scala 508:28 685:39]
  wire [63:0] _GEN_12339 = _T_272 ? mcounteren : _GEN_12321; // @[decode.scala 509:28 685:39]
  wire [63:0] _GEN_12340 = _T_272 ? mscratch : _GEN_12322; // @[decode.scala 510:28 685:39]
  wire [63:0] _GEN_12341 = _T_272 ? mepc : _GEN_12323; // @[decode.scala 511:28 685:39]
  wire [63:0] _GEN_12342 = _T_272 ? mcause : _GEN_12324; // @[decode.scala 512:28 685:39]
  wire [63:0] _GEN_12343 = _T_272 ? mtval : _GEN_12325; // @[decode.scala 513:28 685:39]
  wire [63:0] _GEN_12344 = _T_272 ? mip : _GEN_12326; // @[decode.scala 514:28 685:39]
  wire [63:0] _GEN_12345 = _T_272 ? pmpcfg0 : _GEN_12327; // @[decode.scala 515:28 685:39]
  wire [63:0] _GEN_12346 = _T_272 ? pmpaddr0 : _GEN_12328; // @[decode.scala 516:28 685:39]
  wire [63:0] _GEN_12347 = _T_272 ? mvendorid : _GEN_12329; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12348 = _T_272 ? marchid : _GEN_12330; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12349 = _T_272 ? mimpid : _GEN_12331; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12350 = _T_272 ? mhartid : _GEN_12332; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12351 = _T_271 ? _satp_T_3 : satp; // @[decode.scala 502:28 685:39 691:38]
  wire [63:0] _GEN_12352 = _T_271 ? _mstatus_T_1 : _GEN_12333; // @[decode.scala 522:11 685:39]
  wire [126:0] _GEN_12353 = _T_271 ? 127'h8000000000101101 : _GEN_12334; // @[decode.scala 685:39 523:8]
  wire [63:0] _GEN_12354 = _T_271 ? medeleg : _GEN_12335; // @[decode.scala 505:28 685:39]
  wire [63:0] _GEN_12355 = _T_271 ? mideleg : _GEN_12336; // @[decode.scala 506:28 685:39]
  wire [63:0] _GEN_12356 = _T_271 ? mie : _GEN_12337; // @[decode.scala 507:28 685:39]
  wire [63:0] _GEN_12357 = _T_271 ? mtvec : _GEN_12338; // @[decode.scala 508:28 685:39]
  wire [63:0] _GEN_12358 = _T_271 ? mcounteren : _GEN_12339; // @[decode.scala 509:28 685:39]
  wire [63:0] _GEN_12359 = _T_271 ? mscratch : _GEN_12340; // @[decode.scala 510:28 685:39]
  wire [63:0] _GEN_12360 = _T_271 ? mepc : _GEN_12341; // @[decode.scala 511:28 685:39]
  wire [63:0] _GEN_12361 = _T_271 ? mcause : _GEN_12342; // @[decode.scala 512:28 685:39]
  wire [63:0] _GEN_12362 = _T_271 ? mtval : _GEN_12343; // @[decode.scala 513:28 685:39]
  wire [63:0] _GEN_12363 = _T_271 ? mip : _GEN_12344; // @[decode.scala 514:28 685:39]
  wire [63:0] _GEN_12364 = _T_271 ? pmpcfg0 : _GEN_12345; // @[decode.scala 515:28 685:39]
  wire [63:0] _GEN_12365 = _T_271 ? pmpaddr0 : _GEN_12346; // @[decode.scala 516:28 685:39]
  wire [63:0] _GEN_12366 = _T_271 ? mvendorid : _GEN_12347; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12367 = _T_271 ? marchid : _GEN_12348; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12368 = _T_271 ? mimpid : _GEN_12349; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12369 = _T_271 ? mhartid : _GEN_12350; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12370 = _T_270 ? _scounteren_T_3 : scounteren; // @[decode.scala 501:28 685:39 690:38]
  wire [63:0] _GEN_12371 = _T_270 ? satp : _GEN_12351; // @[decode.scala 502:28 685:39]
  wire [63:0] _GEN_12372 = _T_270 ? _mstatus_T_1 : _GEN_12352; // @[decode.scala 522:11 685:39]
  wire [126:0] _GEN_12373 = _T_270 ? 127'h8000000000101101 : _GEN_12353; // @[decode.scala 685:39 523:8]
  wire [63:0] _GEN_12374 = _T_270 ? medeleg : _GEN_12354; // @[decode.scala 505:28 685:39]
  wire [63:0] _GEN_12375 = _T_270 ? mideleg : _GEN_12355; // @[decode.scala 506:28 685:39]
  wire [63:0] _GEN_12376 = _T_270 ? mie : _GEN_12356; // @[decode.scala 507:28 685:39]
  wire [63:0] _GEN_12377 = _T_270 ? mtvec : _GEN_12357; // @[decode.scala 508:28 685:39]
  wire [63:0] _GEN_12378 = _T_270 ? mcounteren : _GEN_12358; // @[decode.scala 509:28 685:39]
  wire [63:0] _GEN_12379 = _T_270 ? mscratch : _GEN_12359; // @[decode.scala 510:28 685:39]
  wire [63:0] _GEN_12380 = _T_270 ? mepc : _GEN_12360; // @[decode.scala 511:28 685:39]
  wire [63:0] _GEN_12381 = _T_270 ? mcause : _GEN_12361; // @[decode.scala 512:28 685:39]
  wire [63:0] _GEN_12382 = _T_270 ? mtval : _GEN_12362; // @[decode.scala 513:28 685:39]
  wire [63:0] _GEN_12383 = _T_270 ? mip : _GEN_12363; // @[decode.scala 514:28 685:39]
  wire [63:0] _GEN_12384 = _T_270 ? pmpcfg0 : _GEN_12364; // @[decode.scala 515:28 685:39]
  wire [63:0] _GEN_12385 = _T_270 ? pmpaddr0 : _GEN_12365; // @[decode.scala 516:28 685:39]
  wire [63:0] _GEN_12386 = _T_270 ? mvendorid : _GEN_12366; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12387 = _T_270 ? marchid : _GEN_12367; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12388 = _T_270 ? mimpid : _GEN_12368; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12389 = _T_270 ? mhartid : _GEN_12369; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12390 = _T_269 ? _ucause_T_3 : ucause; // @[decode.scala 500:28 685:39 689:38]
  wire [63:0] _GEN_12391 = _T_269 ? scounteren : _GEN_12370; // @[decode.scala 501:28 685:39]
  wire [63:0] _GEN_12392 = _T_269 ? satp : _GEN_12371; // @[decode.scala 502:28 685:39]
  wire [63:0] _GEN_12393 = _T_269 ? _mstatus_T_1 : _GEN_12372; // @[decode.scala 522:11 685:39]
  wire [126:0] _GEN_12394 = _T_269 ? 127'h8000000000101101 : _GEN_12373; // @[decode.scala 685:39 523:8]
  wire [63:0] _GEN_12395 = _T_269 ? medeleg : _GEN_12374; // @[decode.scala 505:28 685:39]
  wire [63:0] _GEN_12396 = _T_269 ? mideleg : _GEN_12375; // @[decode.scala 506:28 685:39]
  wire [63:0] _GEN_12397 = _T_269 ? mie : _GEN_12376; // @[decode.scala 507:28 685:39]
  wire [63:0] _GEN_12398 = _T_269 ? mtvec : _GEN_12377; // @[decode.scala 508:28 685:39]
  wire [63:0] _GEN_12399 = _T_269 ? mcounteren : _GEN_12378; // @[decode.scala 509:28 685:39]
  wire [63:0] _GEN_12400 = _T_269 ? mscratch : _GEN_12379; // @[decode.scala 510:28 685:39]
  wire [63:0] _GEN_12401 = _T_269 ? mepc : _GEN_12380; // @[decode.scala 511:28 685:39]
  wire [63:0] _GEN_12402 = _T_269 ? mcause : _GEN_12381; // @[decode.scala 512:28 685:39]
  wire [63:0] _GEN_12403 = _T_269 ? mtval : _GEN_12382; // @[decode.scala 513:28 685:39]
  wire [63:0] _GEN_12404 = _T_269 ? mip : _GEN_12383; // @[decode.scala 514:28 685:39]
  wire [63:0] _GEN_12405 = _T_269 ? pmpcfg0 : _GEN_12384; // @[decode.scala 515:28 685:39]
  wire [63:0] _GEN_12406 = _T_269 ? pmpaddr0 : _GEN_12385; // @[decode.scala 516:28 685:39]
  wire [63:0] _GEN_12407 = _T_269 ? mvendorid : _GEN_12386; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12408 = _T_269 ? marchid : _GEN_12387; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12409 = _T_269 ? mimpid : _GEN_12388; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12410 = _T_269 ? mhartid : _GEN_12389; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12411 = _T_268 ? _uepc_T_3 : uepc; // @[decode.scala 499:28 685:39 688:38]
  wire [63:0] _GEN_12412 = _T_268 ? ucause : _GEN_12390; // @[decode.scala 500:28 685:39]
  wire [63:0] _GEN_12413 = _T_268 ? scounteren : _GEN_12391; // @[decode.scala 501:28 685:39]
  wire [63:0] _GEN_12414 = _T_268 ? satp : _GEN_12392; // @[decode.scala 502:28 685:39]
  wire [63:0] _GEN_12415 = _T_268 ? _mstatus_T_1 : _GEN_12393; // @[decode.scala 522:11 685:39]
  wire [126:0] _GEN_12416 = _T_268 ? 127'h8000000000101101 : _GEN_12394; // @[decode.scala 685:39 523:8]
  wire [63:0] _GEN_12417 = _T_268 ? medeleg : _GEN_12395; // @[decode.scala 505:28 685:39]
  wire [63:0] _GEN_12418 = _T_268 ? mideleg : _GEN_12396; // @[decode.scala 506:28 685:39]
  wire [63:0] _GEN_12419 = _T_268 ? mie : _GEN_12397; // @[decode.scala 507:28 685:39]
  wire [63:0] _GEN_12420 = _T_268 ? mtvec : _GEN_12398; // @[decode.scala 508:28 685:39]
  wire [63:0] _GEN_12421 = _T_268 ? mcounteren : _GEN_12399; // @[decode.scala 509:28 685:39]
  wire [63:0] _GEN_12422 = _T_268 ? mscratch : _GEN_12400; // @[decode.scala 510:28 685:39]
  wire [63:0] _GEN_12423 = _T_268 ? mepc : _GEN_12401; // @[decode.scala 511:28 685:39]
  wire [63:0] _GEN_12424 = _T_268 ? mcause : _GEN_12402; // @[decode.scala 512:28 685:39]
  wire [63:0] _GEN_12425 = _T_268 ? mtval : _GEN_12403; // @[decode.scala 513:28 685:39]
  wire [63:0] _GEN_12426 = _T_268 ? mip : _GEN_12404; // @[decode.scala 514:28 685:39]
  wire [63:0] _GEN_12427 = _T_268 ? pmpcfg0 : _GEN_12405; // @[decode.scala 515:28 685:39]
  wire [63:0] _GEN_12428 = _T_268 ? pmpaddr0 : _GEN_12406; // @[decode.scala 516:28 685:39]
  wire [63:0] _GEN_12429 = _T_268 ? mvendorid : _GEN_12407; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12430 = _T_268 ? marchid : _GEN_12408; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12431 = _T_268 ? mimpid : _GEN_12409; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12432 = _T_268 ? mhartid : _GEN_12410; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12433 = _T_267 ? _utvec_T_3 : utvec; // @[decode.scala 498:28 685:39 687:38]
  wire [63:0] _GEN_12434 = _T_267 ? uepc : _GEN_12411; // @[decode.scala 499:28 685:39]
  wire [63:0] _GEN_12435 = _T_267 ? ucause : _GEN_12412; // @[decode.scala 500:28 685:39]
  wire [63:0] _GEN_12436 = _T_267 ? scounteren : _GEN_12413; // @[decode.scala 501:28 685:39]
  wire [63:0] _GEN_12437 = _T_267 ? satp : _GEN_12414; // @[decode.scala 502:28 685:39]
  wire [63:0] _GEN_12438 = _T_267 ? _mstatus_T_1 : _GEN_12415; // @[decode.scala 522:11 685:39]
  wire [126:0] _GEN_12439 = _T_267 ? 127'h8000000000101101 : _GEN_12416; // @[decode.scala 685:39 523:8]
  wire [63:0] _GEN_12440 = _T_267 ? medeleg : _GEN_12417; // @[decode.scala 505:28 685:39]
  wire [63:0] _GEN_12441 = _T_267 ? mideleg : _GEN_12418; // @[decode.scala 506:28 685:39]
  wire [63:0] _GEN_12442 = _T_267 ? mie : _GEN_12419; // @[decode.scala 507:28 685:39]
  wire [63:0] _GEN_12443 = _T_267 ? mtvec : _GEN_12420; // @[decode.scala 508:28 685:39]
  wire [63:0] _GEN_12444 = _T_267 ? mcounteren : _GEN_12421; // @[decode.scala 509:28 685:39]
  wire [63:0] _GEN_12445 = _T_267 ? mscratch : _GEN_12422; // @[decode.scala 510:28 685:39]
  wire [63:0] _GEN_12446 = _T_267 ? mepc : _GEN_12423; // @[decode.scala 511:28 685:39]
  wire [63:0] _GEN_12447 = _T_267 ? mcause : _GEN_12424; // @[decode.scala 512:28 685:39]
  wire [63:0] _GEN_12448 = _T_267 ? mtval : _GEN_12425; // @[decode.scala 513:28 685:39]
  wire [63:0] _GEN_12449 = _T_267 ? mip : _GEN_12426; // @[decode.scala 514:28 685:39]
  wire [63:0] _GEN_12450 = _T_267 ? pmpcfg0 : _GEN_12427; // @[decode.scala 515:28 685:39]
  wire [63:0] _GEN_12451 = _T_267 ? pmpaddr0 : _GEN_12428; // @[decode.scala 516:28 685:39]
  wire [63:0] _GEN_12452 = _T_267 ? mvendorid : _GEN_12429; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12453 = _T_267 ? marchid : _GEN_12430; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12454 = _T_267 ? mimpid : _GEN_12431; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12455 = _T_267 ? mhartid : _GEN_12432; // @[decode.scala 520:28 685:39]
  wire [63:0] _GEN_12456 = _T_266 ? _ustatus_T_3 : ustatus; // @[decode.scala 497:28 685:39 686:38]
  wire [63:0] _GEN_12457 = _T_266 ? utvec : _GEN_12433; // @[decode.scala 498:28 685:39]
  wire [63:0] _GEN_12458 = _T_266 ? uepc : _GEN_12434; // @[decode.scala 499:28 685:39]
  wire [63:0] _GEN_12459 = _T_266 ? ucause : _GEN_12435; // @[decode.scala 500:28 685:39]
  wire [63:0] _GEN_12460 = _T_266 ? scounteren : _GEN_12436; // @[decode.scala 501:28 685:39]
  wire [63:0] _GEN_12461 = _T_266 ? satp : _GEN_12437; // @[decode.scala 502:28 685:39]
  wire [63:0] _GEN_12462 = _T_266 ? _mstatus_T_1 : _GEN_12438; // @[decode.scala 522:11 685:39]
  wire [126:0] _GEN_12463 = _T_266 ? 127'h8000000000101101 : _GEN_12439; // @[decode.scala 685:39 523:8]
  wire [63:0] _GEN_12464 = _T_266 ? medeleg : _GEN_12440; // @[decode.scala 505:28 685:39]
  wire [63:0] _GEN_12465 = _T_266 ? mideleg : _GEN_12441; // @[decode.scala 506:28 685:39]
  wire [63:0] _GEN_12466 = _T_266 ? mie : _GEN_12442; // @[decode.scala 507:28 685:39]
  wire [63:0] _GEN_12467 = _T_266 ? mtvec : _GEN_12443; // @[decode.scala 508:28 685:39]
  wire [63:0] _GEN_12468 = _T_266 ? mcounteren : _GEN_12444; // @[decode.scala 509:28 685:39]
  wire [63:0] _GEN_12469 = _T_266 ? mscratch : _GEN_12445; // @[decode.scala 510:28 685:39]
  wire [63:0] _GEN_12470 = _T_266 ? mepc : _GEN_12446; // @[decode.scala 511:28 685:39]
  wire [63:0] _GEN_12471 = _T_266 ? mcause : _GEN_12447; // @[decode.scala 512:28 685:39]
  wire [63:0] _GEN_12472 = _T_266 ? mtval : _GEN_12448; // @[decode.scala 513:28 685:39]
  wire [63:0] _GEN_12473 = _T_266 ? mip : _GEN_12449; // @[decode.scala 514:28 685:39]
  wire [63:0] _GEN_12474 = _T_266 ? pmpcfg0 : _GEN_12450; // @[decode.scala 515:28 685:39]
  wire [63:0] _GEN_12475 = _T_266 ? pmpaddr0 : _GEN_12451; // @[decode.scala 516:28 685:39]
  wire [63:0] _GEN_12476 = _T_266 ? mvendorid : _GEN_12452; // @[decode.scala 517:28 685:39]
  wire [63:0] _GEN_12477 = _T_266 ? marchid : _GEN_12453; // @[decode.scala 518:28 685:39]
  wire [63:0] _GEN_12478 = _T_266 ? mimpid : _GEN_12454; // @[decode.scala 519:28 685:39]
  wire [63:0] _GEN_12479 = _T_266 ? mhartid : _GEN_12455; // @[decode.scala 520:28 685:39]
  wire [63:0] _ustatus_T_4 = ~csrImmReg; // @[decode.scala 714:51]
  wire [63:0] _ustatus_T_5 = ustatus & _ustatus_T_4; // @[decode.scala 714:49]
  wire [63:0] _utvec_T_5 = utvec & _ustatus_T_4; // @[decode.scala 715:47]
  wire [63:0] _uepc_T_5 = uepc & _ustatus_T_4; // @[decode.scala 716:46]
  wire [63:0] _ucause_T_5 = ucause & _ustatus_T_4; // @[decode.scala 717:48]
  wire [63:0] _scounteren_T_5 = scounteren & _ustatus_T_4; // @[decode.scala 718:52]
  wire [63:0] _satp_T_5 = satp & _ustatus_T_4; // @[decode.scala 719:46]
  wire [63:0] _mstatus_T_7 = mstatus & _ustatus_T_4; // @[decode.scala 720:49]
  wire [63:0] _misa_T_7 = misa & _ustatus_T_4; // @[decode.scala 721:46]
  wire [63:0] _medeleg_T_5 = medeleg & _ustatus_T_4; // @[decode.scala 722:49]
  wire [63:0] _mideleg_T_5 = mideleg & _ustatus_T_4; // @[decode.scala 723:49]
  wire [63:0] _mie_T_5 = mie & _ustatus_T_4; // @[decode.scala 724:45]
  wire [63:0] _mtvec_T_5 = mtvec & _ustatus_T_4; // @[decode.scala 725:47]
  wire [63:0] _mcounteren_T_5 = mcounteren & _ustatus_T_4; // @[decode.scala 726:52]
  wire [63:0] _mscratch_T_5 = mscratch & _ustatus_T_4; // @[decode.scala 727:50]
  wire [63:0] _mepc_T_5 = mepc & _ustatus_T_4; // @[decode.scala 728:46]
  wire [63:0] _mcause_T_5 = mcause & _ustatus_T_4; // @[decode.scala 729:48]
  wire [63:0] _mtval_T_5 = mtval & _ustatus_T_4; // @[decode.scala 730:47]
  wire [63:0] _mip_T_5 = mip & _ustatus_T_4; // @[decode.scala 731:45]
  wire [63:0] _pmpcfg0_T_5 = pmpcfg0 & _ustatus_T_4; // @[decode.scala 732:49]
  wire [63:0] _pmpaddr0_T_5 = pmpaddr0 & _ustatus_T_4; // @[decode.scala 733:50]
  wire [63:0] _mvendorid_T_5 = mvendorid & _ustatus_T_4; // @[decode.scala 734:51]
  wire [63:0] _marchid_T_5 = marchid & _ustatus_T_4; // @[decode.scala 735:49]
  wire [63:0] _mimpid_T_5 = mimpid & _ustatus_T_4; // @[decode.scala 736:48]
  wire [63:0] _mhartid_T_5 = mhartid & _ustatus_T_4; // @[decode.scala 737:49]
  wire [63:0] _GEN_12480 = _T_289 ? _mhartid_T_5 : mhartid; // @[decode.scala 520:28 713:39 737:38]
  wire [63:0] _GEN_12481 = _T_288 ? _mimpid_T_5 : mimpid; // @[decode.scala 519:28 713:39 736:38]
  wire [63:0] _GEN_12482 = _T_288 ? mhartid : _GEN_12480; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12483 = _T_287 ? _marchid_T_5 : marchid; // @[decode.scala 518:28 713:39 735:38]
  wire [63:0] _GEN_12484 = _T_287 ? mimpid : _GEN_12481; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12485 = _T_287 ? mhartid : _GEN_12482; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12486 = _T_286 ? _mvendorid_T_5 : mvendorid; // @[decode.scala 517:28 713:39 734:38]
  wire [63:0] _GEN_12487 = _T_286 ? marchid : _GEN_12483; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12488 = _T_286 ? mimpid : _GEN_12484; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12489 = _T_286 ? mhartid : _GEN_12485; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12490 = _T_285 ? _pmpaddr0_T_5 : pmpaddr0; // @[decode.scala 516:28 713:39 733:38]
  wire [63:0] _GEN_12491 = _T_285 ? mvendorid : _GEN_12486; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12492 = _T_285 ? marchid : _GEN_12487; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12493 = _T_285 ? mimpid : _GEN_12488; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12494 = _T_285 ? mhartid : _GEN_12489; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12495 = _T_284 ? _pmpcfg0_T_5 : pmpcfg0; // @[decode.scala 515:28 713:39 732:38]
  wire [63:0] _GEN_12496 = _T_284 ? pmpaddr0 : _GEN_12490; // @[decode.scala 516:28 713:39]
  wire [63:0] _GEN_12497 = _T_284 ? mvendorid : _GEN_12491; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12498 = _T_284 ? marchid : _GEN_12492; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12499 = _T_284 ? mimpid : _GEN_12493; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12500 = _T_284 ? mhartid : _GEN_12494; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12501 = _T_283 ? _mip_T_5 : mip; // @[decode.scala 514:28 713:39 731:38]
  wire [63:0] _GEN_12502 = _T_283 ? pmpcfg0 : _GEN_12495; // @[decode.scala 515:28 713:39]
  wire [63:0] _GEN_12503 = _T_283 ? pmpaddr0 : _GEN_12496; // @[decode.scala 516:28 713:39]
  wire [63:0] _GEN_12504 = _T_283 ? mvendorid : _GEN_12497; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12505 = _T_283 ? marchid : _GEN_12498; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12506 = _T_283 ? mimpid : _GEN_12499; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12507 = _T_283 ? mhartid : _GEN_12500; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12508 = _T_282 ? _mtval_T_5 : mtval; // @[decode.scala 513:28 713:39 730:38]
  wire [63:0] _GEN_12509 = _T_282 ? mip : _GEN_12501; // @[decode.scala 514:28 713:39]
  wire [63:0] _GEN_12510 = _T_282 ? pmpcfg0 : _GEN_12502; // @[decode.scala 515:28 713:39]
  wire [63:0] _GEN_12511 = _T_282 ? pmpaddr0 : _GEN_12503; // @[decode.scala 516:28 713:39]
  wire [63:0] _GEN_12512 = _T_282 ? mvendorid : _GEN_12504; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12513 = _T_282 ? marchid : _GEN_12505; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12514 = _T_282 ? mimpid : _GEN_12506; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12515 = _T_282 ? mhartid : _GEN_12507; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12516 = _T_281 ? _mcause_T_5 : mcause; // @[decode.scala 512:28 713:39 729:38]
  wire [63:0] _GEN_12517 = _T_281 ? mtval : _GEN_12508; // @[decode.scala 513:28 713:39]
  wire [63:0] _GEN_12518 = _T_281 ? mip : _GEN_12509; // @[decode.scala 514:28 713:39]
  wire [63:0] _GEN_12519 = _T_281 ? pmpcfg0 : _GEN_12510; // @[decode.scala 515:28 713:39]
  wire [63:0] _GEN_12520 = _T_281 ? pmpaddr0 : _GEN_12511; // @[decode.scala 516:28 713:39]
  wire [63:0] _GEN_12521 = _T_281 ? mvendorid : _GEN_12512; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12522 = _T_281 ? marchid : _GEN_12513; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12523 = _T_281 ? mimpid : _GEN_12514; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12524 = _T_281 ? mhartid : _GEN_12515; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12525 = _T_280 ? _mepc_T_5 : mepc; // @[decode.scala 511:28 713:39 728:38]
  wire [63:0] _GEN_12526 = _T_280 ? mcause : _GEN_12516; // @[decode.scala 512:28 713:39]
  wire [63:0] _GEN_12527 = _T_280 ? mtval : _GEN_12517; // @[decode.scala 513:28 713:39]
  wire [63:0] _GEN_12528 = _T_280 ? mip : _GEN_12518; // @[decode.scala 514:28 713:39]
  wire [63:0] _GEN_12529 = _T_280 ? pmpcfg0 : _GEN_12519; // @[decode.scala 515:28 713:39]
  wire [63:0] _GEN_12530 = _T_280 ? pmpaddr0 : _GEN_12520; // @[decode.scala 516:28 713:39]
  wire [63:0] _GEN_12531 = _T_280 ? mvendorid : _GEN_12521; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12532 = _T_280 ? marchid : _GEN_12522; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12533 = _T_280 ? mimpid : _GEN_12523; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12534 = _T_280 ? mhartid : _GEN_12524; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12535 = _T_279 ? _mscratch_T_5 : mscratch; // @[decode.scala 510:28 713:39 727:38]
  wire [63:0] _GEN_12536 = _T_279 ? mepc : _GEN_12525; // @[decode.scala 511:28 713:39]
  wire [63:0] _GEN_12537 = _T_279 ? mcause : _GEN_12526; // @[decode.scala 512:28 713:39]
  wire [63:0] _GEN_12538 = _T_279 ? mtval : _GEN_12527; // @[decode.scala 513:28 713:39]
  wire [63:0] _GEN_12539 = _T_279 ? mip : _GEN_12528; // @[decode.scala 514:28 713:39]
  wire [63:0] _GEN_12540 = _T_279 ? pmpcfg0 : _GEN_12529; // @[decode.scala 515:28 713:39]
  wire [63:0] _GEN_12541 = _T_279 ? pmpaddr0 : _GEN_12530; // @[decode.scala 516:28 713:39]
  wire [63:0] _GEN_12542 = _T_279 ? mvendorid : _GEN_12531; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12543 = _T_279 ? marchid : _GEN_12532; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12544 = _T_279 ? mimpid : _GEN_12533; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12545 = _T_279 ? mhartid : _GEN_12534; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12546 = _T_278 ? _mcounteren_T_5 : mcounteren; // @[decode.scala 509:28 713:39 726:38]
  wire [63:0] _GEN_12547 = _T_278 ? mscratch : _GEN_12535; // @[decode.scala 510:28 713:39]
  wire [63:0] _GEN_12548 = _T_278 ? mepc : _GEN_12536; // @[decode.scala 511:28 713:39]
  wire [63:0] _GEN_12549 = _T_278 ? mcause : _GEN_12537; // @[decode.scala 512:28 713:39]
  wire [63:0] _GEN_12550 = _T_278 ? mtval : _GEN_12538; // @[decode.scala 513:28 713:39]
  wire [63:0] _GEN_12551 = _T_278 ? mip : _GEN_12539; // @[decode.scala 514:28 713:39]
  wire [63:0] _GEN_12552 = _T_278 ? pmpcfg0 : _GEN_12540; // @[decode.scala 515:28 713:39]
  wire [63:0] _GEN_12553 = _T_278 ? pmpaddr0 : _GEN_12541; // @[decode.scala 516:28 713:39]
  wire [63:0] _GEN_12554 = _T_278 ? mvendorid : _GEN_12542; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12555 = _T_278 ? marchid : _GEN_12543; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12556 = _T_278 ? mimpid : _GEN_12544; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12557 = _T_278 ? mhartid : _GEN_12545; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12558 = _T_277 ? _mtvec_T_5 : mtvec; // @[decode.scala 508:28 713:39 725:38]
  wire [63:0] _GEN_12559 = _T_277 ? mcounteren : _GEN_12546; // @[decode.scala 509:28 713:39]
  wire [63:0] _GEN_12560 = _T_277 ? mscratch : _GEN_12547; // @[decode.scala 510:28 713:39]
  wire [63:0] _GEN_12561 = _T_277 ? mepc : _GEN_12548; // @[decode.scala 511:28 713:39]
  wire [63:0] _GEN_12562 = _T_277 ? mcause : _GEN_12549; // @[decode.scala 512:28 713:39]
  wire [63:0] _GEN_12563 = _T_277 ? mtval : _GEN_12550; // @[decode.scala 513:28 713:39]
  wire [63:0] _GEN_12564 = _T_277 ? mip : _GEN_12551; // @[decode.scala 514:28 713:39]
  wire [63:0] _GEN_12565 = _T_277 ? pmpcfg0 : _GEN_12552; // @[decode.scala 515:28 713:39]
  wire [63:0] _GEN_12566 = _T_277 ? pmpaddr0 : _GEN_12553; // @[decode.scala 516:28 713:39]
  wire [63:0] _GEN_12567 = _T_277 ? mvendorid : _GEN_12554; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12568 = _T_277 ? marchid : _GEN_12555; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12569 = _T_277 ? mimpid : _GEN_12556; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12570 = _T_277 ? mhartid : _GEN_12557; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12571 = _T_276 ? _mie_T_5 : mie; // @[decode.scala 507:28 713:39 724:38]
  wire [63:0] _GEN_12572 = _T_276 ? mtvec : _GEN_12558; // @[decode.scala 508:28 713:39]
  wire [63:0] _GEN_12573 = _T_276 ? mcounteren : _GEN_12559; // @[decode.scala 509:28 713:39]
  wire [63:0] _GEN_12574 = _T_276 ? mscratch : _GEN_12560; // @[decode.scala 510:28 713:39]
  wire [63:0] _GEN_12575 = _T_276 ? mepc : _GEN_12561; // @[decode.scala 511:28 713:39]
  wire [63:0] _GEN_12576 = _T_276 ? mcause : _GEN_12562; // @[decode.scala 512:28 713:39]
  wire [63:0] _GEN_12577 = _T_276 ? mtval : _GEN_12563; // @[decode.scala 513:28 713:39]
  wire [63:0] _GEN_12578 = _T_276 ? mip : _GEN_12564; // @[decode.scala 514:28 713:39]
  wire [63:0] _GEN_12579 = _T_276 ? pmpcfg0 : _GEN_12565; // @[decode.scala 515:28 713:39]
  wire [63:0] _GEN_12580 = _T_276 ? pmpaddr0 : _GEN_12566; // @[decode.scala 516:28 713:39]
  wire [63:0] _GEN_12581 = _T_276 ? mvendorid : _GEN_12567; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12582 = _T_276 ? marchid : _GEN_12568; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12583 = _T_276 ? mimpid : _GEN_12569; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12584 = _T_276 ? mhartid : _GEN_12570; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12585 = _T_275 ? _mideleg_T_5 : mideleg; // @[decode.scala 506:28 713:39 723:38]
  wire [63:0] _GEN_12586 = _T_275 ? mie : _GEN_12571; // @[decode.scala 507:28 713:39]
  wire [63:0] _GEN_12587 = _T_275 ? mtvec : _GEN_12572; // @[decode.scala 508:28 713:39]
  wire [63:0] _GEN_12588 = _T_275 ? mcounteren : _GEN_12573; // @[decode.scala 509:28 713:39]
  wire [63:0] _GEN_12589 = _T_275 ? mscratch : _GEN_12574; // @[decode.scala 510:28 713:39]
  wire [63:0] _GEN_12590 = _T_275 ? mepc : _GEN_12575; // @[decode.scala 511:28 713:39]
  wire [63:0] _GEN_12591 = _T_275 ? mcause : _GEN_12576; // @[decode.scala 512:28 713:39]
  wire [63:0] _GEN_12592 = _T_275 ? mtval : _GEN_12577; // @[decode.scala 513:28 713:39]
  wire [63:0] _GEN_12593 = _T_275 ? mip : _GEN_12578; // @[decode.scala 514:28 713:39]
  wire [63:0] _GEN_12594 = _T_275 ? pmpcfg0 : _GEN_12579; // @[decode.scala 515:28 713:39]
  wire [63:0] _GEN_12595 = _T_275 ? pmpaddr0 : _GEN_12580; // @[decode.scala 516:28 713:39]
  wire [63:0] _GEN_12596 = _T_275 ? mvendorid : _GEN_12581; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12597 = _T_275 ? marchid : _GEN_12582; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12598 = _T_275 ? mimpid : _GEN_12583; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12599 = _T_275 ? mhartid : _GEN_12584; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12600 = _T_274 ? _medeleg_T_5 : medeleg; // @[decode.scala 505:28 713:39 722:38]
  wire [63:0] _GEN_12601 = _T_274 ? mideleg : _GEN_12585; // @[decode.scala 506:28 713:39]
  wire [63:0] _GEN_12602 = _T_274 ? mie : _GEN_12586; // @[decode.scala 507:28 713:39]
  wire [63:0] _GEN_12603 = _T_274 ? mtvec : _GEN_12587; // @[decode.scala 508:28 713:39]
  wire [63:0] _GEN_12604 = _T_274 ? mcounteren : _GEN_12588; // @[decode.scala 509:28 713:39]
  wire [63:0] _GEN_12605 = _T_274 ? mscratch : _GEN_12589; // @[decode.scala 510:28 713:39]
  wire [63:0] _GEN_12606 = _T_274 ? mepc : _GEN_12590; // @[decode.scala 511:28 713:39]
  wire [63:0] _GEN_12607 = _T_274 ? mcause : _GEN_12591; // @[decode.scala 512:28 713:39]
  wire [63:0] _GEN_12608 = _T_274 ? mtval : _GEN_12592; // @[decode.scala 513:28 713:39]
  wire [63:0] _GEN_12609 = _T_274 ? mip : _GEN_12593; // @[decode.scala 514:28 713:39]
  wire [63:0] _GEN_12610 = _T_274 ? pmpcfg0 : _GEN_12594; // @[decode.scala 515:28 713:39]
  wire [63:0] _GEN_12611 = _T_274 ? pmpaddr0 : _GEN_12595; // @[decode.scala 516:28 713:39]
  wire [63:0] _GEN_12612 = _T_274 ? mvendorid : _GEN_12596; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12613 = _T_274 ? marchid : _GEN_12597; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12614 = _T_274 ? mimpid : _GEN_12598; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12615 = _T_274 ? mhartid : _GEN_12599; // @[decode.scala 520:28 713:39]
  wire [126:0] _GEN_12616 = _T_273 ? {{63'd0}, _misa_T_7} : 127'h8000000000101101; // @[decode.scala 713:39 721:38 523:8]
  wire [63:0] _GEN_12617 = _T_273 ? medeleg : _GEN_12600; // @[decode.scala 505:28 713:39]
  wire [63:0] _GEN_12618 = _T_273 ? mideleg : _GEN_12601; // @[decode.scala 506:28 713:39]
  wire [63:0] _GEN_12619 = _T_273 ? mie : _GEN_12602; // @[decode.scala 507:28 713:39]
  wire [63:0] _GEN_12620 = _T_273 ? mtvec : _GEN_12603; // @[decode.scala 508:28 713:39]
  wire [63:0] _GEN_12621 = _T_273 ? mcounteren : _GEN_12604; // @[decode.scala 509:28 713:39]
  wire [63:0] _GEN_12622 = _T_273 ? mscratch : _GEN_12605; // @[decode.scala 510:28 713:39]
  wire [63:0] _GEN_12623 = _T_273 ? mepc : _GEN_12606; // @[decode.scala 511:28 713:39]
  wire [63:0] _GEN_12624 = _T_273 ? mcause : _GEN_12607; // @[decode.scala 512:28 713:39]
  wire [63:0] _GEN_12625 = _T_273 ? mtval : _GEN_12608; // @[decode.scala 513:28 713:39]
  wire [63:0] _GEN_12626 = _T_273 ? mip : _GEN_12609; // @[decode.scala 514:28 713:39]
  wire [63:0] _GEN_12627 = _T_273 ? pmpcfg0 : _GEN_12610; // @[decode.scala 515:28 713:39]
  wire [63:0] _GEN_12628 = _T_273 ? pmpaddr0 : _GEN_12611; // @[decode.scala 516:28 713:39]
  wire [63:0] _GEN_12629 = _T_273 ? mvendorid : _GEN_12612; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12630 = _T_273 ? marchid : _GEN_12613; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12631 = _T_273 ? mimpid : _GEN_12614; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12632 = _T_273 ? mhartid : _GEN_12615; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12633 = _T_272 ? _mstatus_T_7 : _mstatus_T_1; // @[decode.scala 522:11 713:39 720:38]
  wire [126:0] _GEN_12634 = _T_272 ? 127'h8000000000101101 : _GEN_12616; // @[decode.scala 713:39 523:8]
  wire [63:0] _GEN_12635 = _T_272 ? medeleg : _GEN_12617; // @[decode.scala 505:28 713:39]
  wire [63:0] _GEN_12636 = _T_272 ? mideleg : _GEN_12618; // @[decode.scala 506:28 713:39]
  wire [63:0] _GEN_12637 = _T_272 ? mie : _GEN_12619; // @[decode.scala 507:28 713:39]
  wire [63:0] _GEN_12638 = _T_272 ? mtvec : _GEN_12620; // @[decode.scala 508:28 713:39]
  wire [63:0] _GEN_12639 = _T_272 ? mcounteren : _GEN_12621; // @[decode.scala 509:28 713:39]
  wire [63:0] _GEN_12640 = _T_272 ? mscratch : _GEN_12622; // @[decode.scala 510:28 713:39]
  wire [63:0] _GEN_12641 = _T_272 ? mepc : _GEN_12623; // @[decode.scala 511:28 713:39]
  wire [63:0] _GEN_12642 = _T_272 ? mcause : _GEN_12624; // @[decode.scala 512:28 713:39]
  wire [63:0] _GEN_12643 = _T_272 ? mtval : _GEN_12625; // @[decode.scala 513:28 713:39]
  wire [63:0] _GEN_12644 = _T_272 ? mip : _GEN_12626; // @[decode.scala 514:28 713:39]
  wire [63:0] _GEN_12645 = _T_272 ? pmpcfg0 : _GEN_12627; // @[decode.scala 515:28 713:39]
  wire [63:0] _GEN_12646 = _T_272 ? pmpaddr0 : _GEN_12628; // @[decode.scala 516:28 713:39]
  wire [63:0] _GEN_12647 = _T_272 ? mvendorid : _GEN_12629; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12648 = _T_272 ? marchid : _GEN_12630; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12649 = _T_272 ? mimpid : _GEN_12631; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12650 = _T_272 ? mhartid : _GEN_12632; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12651 = _T_271 ? _satp_T_5 : satp; // @[decode.scala 502:28 713:39 719:38]
  wire [63:0] _GEN_12652 = _T_271 ? _mstatus_T_1 : _GEN_12633; // @[decode.scala 522:11 713:39]
  wire [126:0] _GEN_12653 = _T_271 ? 127'h8000000000101101 : _GEN_12634; // @[decode.scala 713:39 523:8]
  wire [63:0] _GEN_12654 = _T_271 ? medeleg : _GEN_12635; // @[decode.scala 505:28 713:39]
  wire [63:0] _GEN_12655 = _T_271 ? mideleg : _GEN_12636; // @[decode.scala 506:28 713:39]
  wire [63:0] _GEN_12656 = _T_271 ? mie : _GEN_12637; // @[decode.scala 507:28 713:39]
  wire [63:0] _GEN_12657 = _T_271 ? mtvec : _GEN_12638; // @[decode.scala 508:28 713:39]
  wire [63:0] _GEN_12658 = _T_271 ? mcounteren : _GEN_12639; // @[decode.scala 509:28 713:39]
  wire [63:0] _GEN_12659 = _T_271 ? mscratch : _GEN_12640; // @[decode.scala 510:28 713:39]
  wire [63:0] _GEN_12660 = _T_271 ? mepc : _GEN_12641; // @[decode.scala 511:28 713:39]
  wire [63:0] _GEN_12661 = _T_271 ? mcause : _GEN_12642; // @[decode.scala 512:28 713:39]
  wire [63:0] _GEN_12662 = _T_271 ? mtval : _GEN_12643; // @[decode.scala 513:28 713:39]
  wire [63:0] _GEN_12663 = _T_271 ? mip : _GEN_12644; // @[decode.scala 514:28 713:39]
  wire [63:0] _GEN_12664 = _T_271 ? pmpcfg0 : _GEN_12645; // @[decode.scala 515:28 713:39]
  wire [63:0] _GEN_12665 = _T_271 ? pmpaddr0 : _GEN_12646; // @[decode.scala 516:28 713:39]
  wire [63:0] _GEN_12666 = _T_271 ? mvendorid : _GEN_12647; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12667 = _T_271 ? marchid : _GEN_12648; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12668 = _T_271 ? mimpid : _GEN_12649; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12669 = _T_271 ? mhartid : _GEN_12650; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12670 = _T_270 ? _scounteren_T_5 : scounteren; // @[decode.scala 501:28 713:39 718:38]
  wire [63:0] _GEN_12671 = _T_270 ? satp : _GEN_12651; // @[decode.scala 502:28 713:39]
  wire [63:0] _GEN_12672 = _T_270 ? _mstatus_T_1 : _GEN_12652; // @[decode.scala 522:11 713:39]
  wire [126:0] _GEN_12673 = _T_270 ? 127'h8000000000101101 : _GEN_12653; // @[decode.scala 713:39 523:8]
  wire [63:0] _GEN_12674 = _T_270 ? medeleg : _GEN_12654; // @[decode.scala 505:28 713:39]
  wire [63:0] _GEN_12675 = _T_270 ? mideleg : _GEN_12655; // @[decode.scala 506:28 713:39]
  wire [63:0] _GEN_12676 = _T_270 ? mie : _GEN_12656; // @[decode.scala 507:28 713:39]
  wire [63:0] _GEN_12677 = _T_270 ? mtvec : _GEN_12657; // @[decode.scala 508:28 713:39]
  wire [63:0] _GEN_12678 = _T_270 ? mcounteren : _GEN_12658; // @[decode.scala 509:28 713:39]
  wire [63:0] _GEN_12679 = _T_270 ? mscratch : _GEN_12659; // @[decode.scala 510:28 713:39]
  wire [63:0] _GEN_12680 = _T_270 ? mepc : _GEN_12660; // @[decode.scala 511:28 713:39]
  wire [63:0] _GEN_12681 = _T_270 ? mcause : _GEN_12661; // @[decode.scala 512:28 713:39]
  wire [63:0] _GEN_12682 = _T_270 ? mtval : _GEN_12662; // @[decode.scala 513:28 713:39]
  wire [63:0] _GEN_12683 = _T_270 ? mip : _GEN_12663; // @[decode.scala 514:28 713:39]
  wire [63:0] _GEN_12684 = _T_270 ? pmpcfg0 : _GEN_12664; // @[decode.scala 515:28 713:39]
  wire [63:0] _GEN_12685 = _T_270 ? pmpaddr0 : _GEN_12665; // @[decode.scala 516:28 713:39]
  wire [63:0] _GEN_12686 = _T_270 ? mvendorid : _GEN_12666; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12687 = _T_270 ? marchid : _GEN_12667; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12688 = _T_270 ? mimpid : _GEN_12668; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12689 = _T_270 ? mhartid : _GEN_12669; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12690 = _T_269 ? _ucause_T_5 : ucause; // @[decode.scala 500:28 713:39 717:38]
  wire [63:0] _GEN_12691 = _T_269 ? scounteren : _GEN_12670; // @[decode.scala 501:28 713:39]
  wire [63:0] _GEN_12692 = _T_269 ? satp : _GEN_12671; // @[decode.scala 502:28 713:39]
  wire [63:0] _GEN_12693 = _T_269 ? _mstatus_T_1 : _GEN_12672; // @[decode.scala 522:11 713:39]
  wire [126:0] _GEN_12694 = _T_269 ? 127'h8000000000101101 : _GEN_12673; // @[decode.scala 713:39 523:8]
  wire [63:0] _GEN_12695 = _T_269 ? medeleg : _GEN_12674; // @[decode.scala 505:28 713:39]
  wire [63:0] _GEN_12696 = _T_269 ? mideleg : _GEN_12675; // @[decode.scala 506:28 713:39]
  wire [63:0] _GEN_12697 = _T_269 ? mie : _GEN_12676; // @[decode.scala 507:28 713:39]
  wire [63:0] _GEN_12698 = _T_269 ? mtvec : _GEN_12677; // @[decode.scala 508:28 713:39]
  wire [63:0] _GEN_12699 = _T_269 ? mcounteren : _GEN_12678; // @[decode.scala 509:28 713:39]
  wire [63:0] _GEN_12700 = _T_269 ? mscratch : _GEN_12679; // @[decode.scala 510:28 713:39]
  wire [63:0] _GEN_12701 = _T_269 ? mepc : _GEN_12680; // @[decode.scala 511:28 713:39]
  wire [63:0] _GEN_12702 = _T_269 ? mcause : _GEN_12681; // @[decode.scala 512:28 713:39]
  wire [63:0] _GEN_12703 = _T_269 ? mtval : _GEN_12682; // @[decode.scala 513:28 713:39]
  wire [63:0] _GEN_12704 = _T_269 ? mip : _GEN_12683; // @[decode.scala 514:28 713:39]
  wire [63:0] _GEN_12705 = _T_269 ? pmpcfg0 : _GEN_12684; // @[decode.scala 515:28 713:39]
  wire [63:0] _GEN_12706 = _T_269 ? pmpaddr0 : _GEN_12685; // @[decode.scala 516:28 713:39]
  wire [63:0] _GEN_12707 = _T_269 ? mvendorid : _GEN_12686; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12708 = _T_269 ? marchid : _GEN_12687; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12709 = _T_269 ? mimpid : _GEN_12688; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12710 = _T_269 ? mhartid : _GEN_12689; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12711 = _T_268 ? _uepc_T_5 : uepc; // @[decode.scala 499:28 713:39 716:38]
  wire [63:0] _GEN_12712 = _T_268 ? ucause : _GEN_12690; // @[decode.scala 500:28 713:39]
  wire [63:0] _GEN_12713 = _T_268 ? scounteren : _GEN_12691; // @[decode.scala 501:28 713:39]
  wire [63:0] _GEN_12714 = _T_268 ? satp : _GEN_12692; // @[decode.scala 502:28 713:39]
  wire [63:0] _GEN_12715 = _T_268 ? _mstatus_T_1 : _GEN_12693; // @[decode.scala 522:11 713:39]
  wire [126:0] _GEN_12716 = _T_268 ? 127'h8000000000101101 : _GEN_12694; // @[decode.scala 713:39 523:8]
  wire [63:0] _GEN_12717 = _T_268 ? medeleg : _GEN_12695; // @[decode.scala 505:28 713:39]
  wire [63:0] _GEN_12718 = _T_268 ? mideleg : _GEN_12696; // @[decode.scala 506:28 713:39]
  wire [63:0] _GEN_12719 = _T_268 ? mie : _GEN_12697; // @[decode.scala 507:28 713:39]
  wire [63:0] _GEN_12720 = _T_268 ? mtvec : _GEN_12698; // @[decode.scala 508:28 713:39]
  wire [63:0] _GEN_12721 = _T_268 ? mcounteren : _GEN_12699; // @[decode.scala 509:28 713:39]
  wire [63:0] _GEN_12722 = _T_268 ? mscratch : _GEN_12700; // @[decode.scala 510:28 713:39]
  wire [63:0] _GEN_12723 = _T_268 ? mepc : _GEN_12701; // @[decode.scala 511:28 713:39]
  wire [63:0] _GEN_12724 = _T_268 ? mcause : _GEN_12702; // @[decode.scala 512:28 713:39]
  wire [63:0] _GEN_12725 = _T_268 ? mtval : _GEN_12703; // @[decode.scala 513:28 713:39]
  wire [63:0] _GEN_12726 = _T_268 ? mip : _GEN_12704; // @[decode.scala 514:28 713:39]
  wire [63:0] _GEN_12727 = _T_268 ? pmpcfg0 : _GEN_12705; // @[decode.scala 515:28 713:39]
  wire [63:0] _GEN_12728 = _T_268 ? pmpaddr0 : _GEN_12706; // @[decode.scala 516:28 713:39]
  wire [63:0] _GEN_12729 = _T_268 ? mvendorid : _GEN_12707; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12730 = _T_268 ? marchid : _GEN_12708; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12731 = _T_268 ? mimpid : _GEN_12709; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12732 = _T_268 ? mhartid : _GEN_12710; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12733 = _T_267 ? _utvec_T_5 : utvec; // @[decode.scala 498:28 713:39 715:38]
  wire [63:0] _GEN_12734 = _T_267 ? uepc : _GEN_12711; // @[decode.scala 499:28 713:39]
  wire [63:0] _GEN_12735 = _T_267 ? ucause : _GEN_12712; // @[decode.scala 500:28 713:39]
  wire [63:0] _GEN_12736 = _T_267 ? scounteren : _GEN_12713; // @[decode.scala 501:28 713:39]
  wire [63:0] _GEN_12737 = _T_267 ? satp : _GEN_12714; // @[decode.scala 502:28 713:39]
  wire [63:0] _GEN_12738 = _T_267 ? _mstatus_T_1 : _GEN_12715; // @[decode.scala 522:11 713:39]
  wire [126:0] _GEN_12739 = _T_267 ? 127'h8000000000101101 : _GEN_12716; // @[decode.scala 713:39 523:8]
  wire [63:0] _GEN_12740 = _T_267 ? medeleg : _GEN_12717; // @[decode.scala 505:28 713:39]
  wire [63:0] _GEN_12741 = _T_267 ? mideleg : _GEN_12718; // @[decode.scala 506:28 713:39]
  wire [63:0] _GEN_12742 = _T_267 ? mie : _GEN_12719; // @[decode.scala 507:28 713:39]
  wire [63:0] _GEN_12743 = _T_267 ? mtvec : _GEN_12720; // @[decode.scala 508:28 713:39]
  wire [63:0] _GEN_12744 = _T_267 ? mcounteren : _GEN_12721; // @[decode.scala 509:28 713:39]
  wire [63:0] _GEN_12745 = _T_267 ? mscratch : _GEN_12722; // @[decode.scala 510:28 713:39]
  wire [63:0] _GEN_12746 = _T_267 ? mepc : _GEN_12723; // @[decode.scala 511:28 713:39]
  wire [63:0] _GEN_12747 = _T_267 ? mcause : _GEN_12724; // @[decode.scala 512:28 713:39]
  wire [63:0] _GEN_12748 = _T_267 ? mtval : _GEN_12725; // @[decode.scala 513:28 713:39]
  wire [63:0] _GEN_12749 = _T_267 ? mip : _GEN_12726; // @[decode.scala 514:28 713:39]
  wire [63:0] _GEN_12750 = _T_267 ? pmpcfg0 : _GEN_12727; // @[decode.scala 515:28 713:39]
  wire [63:0] _GEN_12751 = _T_267 ? pmpaddr0 : _GEN_12728; // @[decode.scala 516:28 713:39]
  wire [63:0] _GEN_12752 = _T_267 ? mvendorid : _GEN_12729; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12753 = _T_267 ? marchid : _GEN_12730; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12754 = _T_267 ? mimpid : _GEN_12731; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12755 = _T_267 ? mhartid : _GEN_12732; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12756 = _T_266 ? _ustatus_T_5 : ustatus; // @[decode.scala 497:28 713:39 714:38]
  wire [63:0] _GEN_12757 = _T_266 ? utvec : _GEN_12733; // @[decode.scala 498:28 713:39]
  wire [63:0] _GEN_12758 = _T_266 ? uepc : _GEN_12734; // @[decode.scala 499:28 713:39]
  wire [63:0] _GEN_12759 = _T_266 ? ucause : _GEN_12735; // @[decode.scala 500:28 713:39]
  wire [63:0] _GEN_12760 = _T_266 ? scounteren : _GEN_12736; // @[decode.scala 501:28 713:39]
  wire [63:0] _GEN_12761 = _T_266 ? satp : _GEN_12737; // @[decode.scala 502:28 713:39]
  wire [63:0] _GEN_12762 = _T_266 ? _mstatus_T_1 : _GEN_12738; // @[decode.scala 522:11 713:39]
  wire [126:0] _GEN_12763 = _T_266 ? 127'h8000000000101101 : _GEN_12739; // @[decode.scala 713:39 523:8]
  wire [63:0] _GEN_12764 = _T_266 ? medeleg : _GEN_12740; // @[decode.scala 505:28 713:39]
  wire [63:0] _GEN_12765 = _T_266 ? mideleg : _GEN_12741; // @[decode.scala 506:28 713:39]
  wire [63:0] _GEN_12766 = _T_266 ? mie : _GEN_12742; // @[decode.scala 507:28 713:39]
  wire [63:0] _GEN_12767 = _T_266 ? mtvec : _GEN_12743; // @[decode.scala 508:28 713:39]
  wire [63:0] _GEN_12768 = _T_266 ? mcounteren : _GEN_12744; // @[decode.scala 509:28 713:39]
  wire [63:0] _GEN_12769 = _T_266 ? mscratch : _GEN_12745; // @[decode.scala 510:28 713:39]
  wire [63:0] _GEN_12770 = _T_266 ? mepc : _GEN_12746; // @[decode.scala 511:28 713:39]
  wire [63:0] _GEN_12771 = _T_266 ? mcause : _GEN_12747; // @[decode.scala 512:28 713:39]
  wire [63:0] _GEN_12772 = _T_266 ? mtval : _GEN_12748; // @[decode.scala 513:28 713:39]
  wire [63:0] _GEN_12773 = _T_266 ? mip : _GEN_12749; // @[decode.scala 514:28 713:39]
  wire [63:0] _GEN_12774 = _T_266 ? pmpcfg0 : _GEN_12750; // @[decode.scala 515:28 713:39]
  wire [63:0] _GEN_12775 = _T_266 ? pmpaddr0 : _GEN_12751; // @[decode.scala 516:28 713:39]
  wire [63:0] _GEN_12776 = _T_266 ? mvendorid : _GEN_12752; // @[decode.scala 517:28 713:39]
  wire [63:0] _GEN_12777 = _T_266 ? marchid : _GEN_12753; // @[decode.scala 518:28 713:39]
  wire [63:0] _GEN_12778 = _T_266 ? mimpid : _GEN_12754; // @[decode.scala 519:28 713:39]
  wire [63:0] _GEN_12779 = _T_266 ? mhartid : _GEN_12755; // @[decode.scala 520:28 713:39]
  wire [63:0] _GEN_12780 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12756 : ustatus; // @[decode.scala 497:28 571:48]
  wire [63:0] _GEN_12781 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12757 : utvec; // @[decode.scala 498:28 571:48]
  wire [63:0] _GEN_12782 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12758 : uepc; // @[decode.scala 499:28 571:48]
  wire [63:0] _GEN_12783 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12759 : ucause; // @[decode.scala 500:28 571:48]
  wire [63:0] _GEN_12784 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12760 : scounteren; // @[decode.scala 501:28 571:48]
  wire [63:0] _GEN_12785 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12761 : satp; // @[decode.scala 502:28 571:48]
  wire [63:0] _GEN_12786 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12762 : _mstatus_T_1; // @[decode.scala 522:11 571:48]
  wire [126:0] _GEN_12787 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12763 : 127'h8000000000101101; // @[decode.scala 571:48 523:8]
  wire [63:0] _GEN_12788 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12764 : medeleg; // @[decode.scala 505:28 571:48]
  wire [63:0] _GEN_12789 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12765 : mideleg; // @[decode.scala 506:28 571:48]
  wire [63:0] _GEN_12790 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12766 : mie; // @[decode.scala 507:28 571:48]
  wire [63:0] _GEN_12791 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12767 : mtvec; // @[decode.scala 508:28 571:48]
  wire [63:0] _GEN_12792 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12768 : mcounteren; // @[decode.scala 509:28 571:48]
  wire [63:0] _GEN_12793 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12769 : mscratch; // @[decode.scala 510:28 571:48]
  wire [63:0] _GEN_12794 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12770 : mepc; // @[decode.scala 511:28 571:48]
  wire [63:0] _GEN_12795 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12771 : mcause; // @[decode.scala 512:28 571:48]
  wire [63:0] _GEN_12796 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12772 : mtval; // @[decode.scala 513:28 571:48]
  wire [63:0] _GEN_12797 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12773 : mip; // @[decode.scala 514:28 571:48]
  wire [63:0] _GEN_12798 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12774 : pmpcfg0; // @[decode.scala 515:28 571:48]
  wire [63:0] _GEN_12799 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12775 : pmpaddr0; // @[decode.scala 516:28 571:48]
  wire [63:0] _GEN_12800 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12776 : mvendorid; // @[decode.scala 517:28 571:48]
  wire [63:0] _GEN_12801 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12777 : marchid; // @[decode.scala 518:28 571:48]
  wire [63:0] _GEN_12802 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12778 : mimpid; // @[decode.scala 519:28 571:48]
  wire [63:0] _GEN_12803 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_12779 : mhartid; // @[decode.scala 520:28 571:48]
  wire [63:0] _GEN_12804 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12456 : _GEN_12780; // @[decode.scala 571:48]
  wire [63:0] _GEN_12805 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12457 : _GEN_12781; // @[decode.scala 571:48]
  wire [63:0] _GEN_12806 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12458 : _GEN_12782; // @[decode.scala 571:48]
  wire [63:0] _GEN_12807 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12459 : _GEN_12783; // @[decode.scala 571:48]
  wire [63:0] _GEN_12808 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12460 : _GEN_12784; // @[decode.scala 571:48]
  wire [63:0] _GEN_12809 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12461 : _GEN_12785; // @[decode.scala 571:48]
  wire [63:0] _GEN_12810 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12462 : _GEN_12786; // @[decode.scala 571:48]
  wire [126:0] _GEN_12811 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12463 : _GEN_12787; // @[decode.scala 571:48]
  wire [63:0] _GEN_12812 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12464 : _GEN_12788; // @[decode.scala 571:48]
  wire [63:0] _GEN_12813 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12465 : _GEN_12789; // @[decode.scala 571:48]
  wire [63:0] _GEN_12814 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12466 : _GEN_12790; // @[decode.scala 571:48]
  wire [63:0] _GEN_12815 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12467 : _GEN_12791; // @[decode.scala 571:48]
  wire [63:0] _GEN_12816 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12468 : _GEN_12792; // @[decode.scala 571:48]
  wire [63:0] _GEN_12817 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12469 : _GEN_12793; // @[decode.scala 571:48]
  wire [63:0] _GEN_12818 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12470 : _GEN_12794; // @[decode.scala 571:48]
  wire [63:0] _GEN_12819 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12471 : _GEN_12795; // @[decode.scala 571:48]
  wire [63:0] _GEN_12820 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12472 : _GEN_12796; // @[decode.scala 571:48]
  wire [63:0] _GEN_12821 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12473 : _GEN_12797; // @[decode.scala 571:48]
  wire [63:0] _GEN_12822 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12474 : _GEN_12798; // @[decode.scala 571:48]
  wire [63:0] _GEN_12823 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12475 : _GEN_12799; // @[decode.scala 571:48]
  wire [63:0] _GEN_12824 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12476 : _GEN_12800; // @[decode.scala 571:48]
  wire [63:0] _GEN_12825 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12477 : _GEN_12801; // @[decode.scala 571:48]
  wire [63:0] _GEN_12826 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12478 : _GEN_12802; // @[decode.scala 571:48]
  wire [63:0] _GEN_12827 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_12479 : _GEN_12803; // @[decode.scala 571:48]
  wire [63:0] _GEN_12828 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12156 : _GEN_12804; // @[decode.scala 571:48]
  wire [63:0] _GEN_12829 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12157 : _GEN_12805; // @[decode.scala 571:48]
  wire [63:0] _GEN_12830 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12158 : _GEN_12806; // @[decode.scala 571:48]
  wire [63:0] _GEN_12831 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12159 : _GEN_12807; // @[decode.scala 571:48]
  wire [63:0] _GEN_12832 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12160 : _GEN_12808; // @[decode.scala 571:48]
  wire [63:0] _GEN_12833 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12161 : _GEN_12809; // @[decode.scala 571:48]
  wire [63:0] _GEN_12834 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12162 : _GEN_12810; // @[decode.scala 571:48]
  wire [126:0] _GEN_12835 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12163 : _GEN_12811; // @[decode.scala 571:48]
  wire [63:0] _GEN_12836 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12164 : _GEN_12812; // @[decode.scala 571:48]
  wire [63:0] _GEN_12837 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12165 : _GEN_12813; // @[decode.scala 571:48]
  wire [63:0] _GEN_12838 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12166 : _GEN_12814; // @[decode.scala 571:48]
  wire [63:0] _GEN_12839 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12167 : _GEN_12815; // @[decode.scala 571:48]
  wire [63:0] _GEN_12840 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12168 : _GEN_12816; // @[decode.scala 571:48]
  wire [63:0] _GEN_12841 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12169 : _GEN_12817; // @[decode.scala 571:48]
  wire [63:0] _GEN_12842 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12170 : _GEN_12818; // @[decode.scala 571:48]
  wire [63:0] _GEN_12843 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12171 : _GEN_12819; // @[decode.scala 571:48]
  wire [63:0] _GEN_12844 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12172 : _GEN_12820; // @[decode.scala 571:48]
  wire [63:0] _GEN_12845 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12173 : _GEN_12821; // @[decode.scala 571:48]
  wire [63:0] _GEN_12846 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12174 : _GEN_12822; // @[decode.scala 571:48]
  wire [63:0] _GEN_12847 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12175 : _GEN_12823; // @[decode.scala 571:48]
  wire [63:0] _GEN_12848 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12176 : _GEN_12824; // @[decode.scala 571:48]
  wire [63:0] _GEN_12849 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12177 : _GEN_12825; // @[decode.scala 571:48]
  wire [63:0] _GEN_12850 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12178 : _GEN_12826; // @[decode.scala 571:48]
  wire [63:0] _GEN_12851 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_12179 : _GEN_12827; // @[decode.scala 571:48]
  wire [63:0] _GEN_12852 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11856 : _GEN_12828; // @[decode.scala 571:48]
  wire [63:0] _GEN_12853 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11857 : _GEN_12829; // @[decode.scala 571:48]
  wire [63:0] _GEN_12854 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11858 : _GEN_12830; // @[decode.scala 571:48]
  wire [63:0] _GEN_12855 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11859 : _GEN_12831; // @[decode.scala 571:48]
  wire [63:0] _GEN_12856 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11860 : _GEN_12832; // @[decode.scala 571:48]
  wire [63:0] _GEN_12857 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11861 : _GEN_12833; // @[decode.scala 571:48]
  wire [63:0] _GEN_12858 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11862 : _GEN_12834; // @[decode.scala 571:48]
  wire [126:0] _GEN_12859 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11863 : _GEN_12835; // @[decode.scala 571:48]
  wire [63:0] _GEN_12860 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11864 : _GEN_12836; // @[decode.scala 571:48]
  wire [63:0] _GEN_12861 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11865 : _GEN_12837; // @[decode.scala 571:48]
  wire [63:0] _GEN_12862 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11866 : _GEN_12838; // @[decode.scala 571:48]
  wire [63:0] _GEN_12863 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11867 : _GEN_12839; // @[decode.scala 571:48]
  wire [63:0] _GEN_12864 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11868 : _GEN_12840; // @[decode.scala 571:48]
  wire [63:0] _GEN_12865 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11869 : _GEN_12841; // @[decode.scala 571:48]
  wire [63:0] _GEN_12866 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11870 : _GEN_12842; // @[decode.scala 571:48]
  wire [63:0] _GEN_12867 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11871 : _GEN_12843; // @[decode.scala 571:48]
  wire [63:0] _GEN_12868 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11872 : _GEN_12844; // @[decode.scala 571:48]
  wire [63:0] _GEN_12869 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11873 : _GEN_12845; // @[decode.scala 571:48]
  wire [63:0] _GEN_12870 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11874 : _GEN_12846; // @[decode.scala 571:48]
  wire [63:0] _GEN_12871 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11875 : _GEN_12847; // @[decode.scala 571:48]
  wire [63:0] _GEN_12872 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11876 : _GEN_12848; // @[decode.scala 571:48]
  wire [63:0] _GEN_12873 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11877 : _GEN_12849; // @[decode.scala 571:48]
  wire [63:0] _GEN_12874 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11878 : _GEN_12850; // @[decode.scala 571:48]
  wire [63:0] _GEN_12875 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_11879 : _GEN_12851; // @[decode.scala 571:48]
  wire [63:0] _GEN_12882 = 3'h2 == writeBackResult_instruction[14:12] ? _GEN_11562 : _GEN_12858; // @[decode.scala 571:48]
  wire [126:0] _GEN_12883 = 3'h2 == writeBackResult_instruction[14:12] ? _GEN_11563 : _GEN_12859; // @[decode.scala 571:48]
  wire [63:0] _GEN_12890 = 3'h2 == writeBackResult_instruction[14:12] ? _GEN_11570 : _GEN_12866; // @[decode.scala 571:48]
  wire [63:0] _GEN_12891 = 3'h2 == writeBackResult_instruction[14:12] ? _GEN_11571 : _GEN_12867; // @[decode.scala 571:48]
  wire [63:0] _GEN_12906 = 3'h1 == writeBackResult_instruction[14:12] ? _GEN_11262 : _GEN_12882; // @[decode.scala 571:48]
  wire [126:0] _GEN_12907 = 3'h1 == writeBackResult_instruction[14:12] ? _GEN_11263 : _GEN_12883; // @[decode.scala 571:48]
  wire [63:0] _GEN_12914 = 3'h1 == writeBackResult_instruction[14:12] ? _GEN_11270 : _GEN_12890; // @[decode.scala 571:48]
  wire [63:0] _GEN_12915 = 3'h1 == writeBackResult_instruction[14:12] ? _GEN_11271 : _GEN_12891; // @[decode.scala 571:48]
  wire [63:0] _GEN_12931 = _T_256 & writeBackResult_instruction[14:12] != 3'h0 ? _GEN_12906 : _mstatus_T_1; // @[decode.scala 522:11 568:126]
  wire [126:0] _GEN_12932 = _T_256 & writeBackResult_instruction[14:12] != 3'h0 ? _GEN_12907 : 127'h8000000000101101; // @[decode.scala 568:126 523:8]
  wire [63:0] _GEN_12939 = _T_256 & writeBackResult_instruction[14:12] != 3'h0 ? _GEN_12914 : mepc; // @[decode.scala 568:126 511:28]
  wire [63:0] _GEN_12940 = _T_256 & writeBackResult_instruction[14:12] != 3'h0 ? _GEN_12915 : mcause; // @[decode.scala 568:126 512:28]
  reg [63:0] currentPrivilege; // @[decode.scala 743:33]
  wire [37:0] _GEN_12950 = mstatus[12] ? 38'h2200000000 : 38'h2200001800; // @[decode.scala 747:{24,24}]
  wire [63:0] _mstatus_T_9 = {60'ha0000008,mstatus[7:4]}; // @[Cat.scala 33:92]
  wire  _T_431 = currentPrivilege == 64'h2200000000; // @[decode.scala 753:29]
  wire [3:0] _GEN_12951 = currentPrivilege == 64'h2200000000 ? 4'hb : 4'h8; // @[decode.scala 753:{42,51} 754:27]
  wire [4:0] _mstatus_T_11 = _T_431 ? 5'h18 : 5'h0; // @[decode.scala 757:66]
  wire [63:0] _mstatus_T_13 = {51'h0,_mstatus_T_11,mstatus[3:0],4'h0}; // @[Cat.scala 33:92]
  wire [63:0] _mstatus_T_14 = 64'ha00000000 | _mstatus_T_13; // @[decode.scala 757:46]
  wire [63:0] _GEN_16101 = {{32'd0}, writeBackResult_instruction}; // @[decode.scala 758:44]
  wire [63:0] _mepc_T_6 = stallReg ? ecallPC : interruptedPC; // @[decode.scala 761:18]
  wire [63:0] _GEN_12952 = _GEN_16101 == 64'h80000073 ? _mepc_T_6 : _GEN_12939; // @[decode.scala 758:69 761:12]
  wire [63:0] _GEN_12953 = _GEN_16101 == 64'h80000073 ? 64'h8000000000000007 : _GEN_12940; // @[decode.scala 758:69 762:14]
  wire [63:0] _GEN_12954 = _GEN_16101 == 64'h80000073 ? 64'h2200000000 : currentPrivilege; // @[decode.scala 758:69 763:24 743:33]
  wire [63:0] _GEN_12955 = _GEN_16101 == 64'h80000073 ? mtvec : _GEN_10945; // @[decode.scala 758:69 764:18]
  wire [63:0] _GEN_12956 = _GEN_16101 == 64'h80000073 ? _mstatus_T_14 : _GEN_12931; // @[decode.scala 758:69 765:15]
  wire  _GEN_13036 = writeAddrPRF_exec1Valid ? 6'h0 == writeAddrPRF_exec1Addr | _GEN_6212 : _GEN_6212; // @[decode.scala 784:33]
  wire  _GEN_13037 = writeAddrPRF_exec1Valid ? 6'h1 == writeAddrPRF_exec1Addr | _GEN_6213 : _GEN_6213; // @[decode.scala 784:33]
  wire  _GEN_13038 = writeAddrPRF_exec1Valid ? 6'h2 == writeAddrPRF_exec1Addr | _GEN_6214 : _GEN_6214; // @[decode.scala 784:33]
  wire  _GEN_13039 = writeAddrPRF_exec1Valid ? 6'h3 == writeAddrPRF_exec1Addr | _GEN_6215 : _GEN_6215; // @[decode.scala 784:33]
  wire  _GEN_13040 = writeAddrPRF_exec1Valid ? 6'h4 == writeAddrPRF_exec1Addr | _GEN_6216 : _GEN_6216; // @[decode.scala 784:33]
  wire  _GEN_13041 = writeAddrPRF_exec1Valid ? 6'h5 == writeAddrPRF_exec1Addr | _GEN_6217 : _GEN_6217; // @[decode.scala 784:33]
  wire  _GEN_13042 = writeAddrPRF_exec1Valid ? 6'h6 == writeAddrPRF_exec1Addr | _GEN_6218 : _GEN_6218; // @[decode.scala 784:33]
  wire  _GEN_13043 = writeAddrPRF_exec1Valid ? 6'h7 == writeAddrPRF_exec1Addr | _GEN_6219 : _GEN_6219; // @[decode.scala 784:33]
  wire  _GEN_13044 = writeAddrPRF_exec1Valid ? 6'h8 == writeAddrPRF_exec1Addr | _GEN_6220 : _GEN_6220; // @[decode.scala 784:33]
  wire  _GEN_13045 = writeAddrPRF_exec1Valid ? 6'h9 == writeAddrPRF_exec1Addr | _GEN_6221 : _GEN_6221; // @[decode.scala 784:33]
  wire  _GEN_13046 = writeAddrPRF_exec1Valid ? 6'ha == writeAddrPRF_exec1Addr | _GEN_6222 : _GEN_6222; // @[decode.scala 784:33]
  wire  _GEN_13047 = writeAddrPRF_exec1Valid ? 6'hb == writeAddrPRF_exec1Addr | _GEN_6223 : _GEN_6223; // @[decode.scala 784:33]
  wire  _GEN_13048 = writeAddrPRF_exec1Valid ? 6'hc == writeAddrPRF_exec1Addr | _GEN_6224 : _GEN_6224; // @[decode.scala 784:33]
  wire  _GEN_13049 = writeAddrPRF_exec1Valid ? 6'hd == writeAddrPRF_exec1Addr | _GEN_6225 : _GEN_6225; // @[decode.scala 784:33]
  wire  _GEN_13050 = writeAddrPRF_exec1Valid ? 6'he == writeAddrPRF_exec1Addr | _GEN_6226 : _GEN_6226; // @[decode.scala 784:33]
  wire  _GEN_13051 = writeAddrPRF_exec1Valid ? 6'hf == writeAddrPRF_exec1Addr | _GEN_6227 : _GEN_6227; // @[decode.scala 784:33]
  wire  _GEN_13052 = writeAddrPRF_exec1Valid ? 6'h10 == writeAddrPRF_exec1Addr | _GEN_6228 : _GEN_6228; // @[decode.scala 784:33]
  wire  _GEN_13053 = writeAddrPRF_exec1Valid ? 6'h11 == writeAddrPRF_exec1Addr | _GEN_6229 : _GEN_6229; // @[decode.scala 784:33]
  wire  _GEN_13054 = writeAddrPRF_exec1Valid ? 6'h12 == writeAddrPRF_exec1Addr | _GEN_6230 : _GEN_6230; // @[decode.scala 784:33]
  wire  _GEN_13055 = writeAddrPRF_exec1Valid ? 6'h13 == writeAddrPRF_exec1Addr | _GEN_6231 : _GEN_6231; // @[decode.scala 784:33]
  wire  _GEN_13056 = writeAddrPRF_exec1Valid ? 6'h14 == writeAddrPRF_exec1Addr | _GEN_6232 : _GEN_6232; // @[decode.scala 784:33]
  wire  _GEN_13057 = writeAddrPRF_exec1Valid ? 6'h15 == writeAddrPRF_exec1Addr | _GEN_6233 : _GEN_6233; // @[decode.scala 784:33]
  wire  _GEN_13058 = writeAddrPRF_exec1Valid ? 6'h16 == writeAddrPRF_exec1Addr | _GEN_6234 : _GEN_6234; // @[decode.scala 784:33]
  wire  _GEN_13059 = writeAddrPRF_exec1Valid ? 6'h17 == writeAddrPRF_exec1Addr | _GEN_6235 : _GEN_6235; // @[decode.scala 784:33]
  wire  _GEN_13060 = writeAddrPRF_exec1Valid ? 6'h18 == writeAddrPRF_exec1Addr | _GEN_6236 : _GEN_6236; // @[decode.scala 784:33]
  wire  _GEN_13061 = writeAddrPRF_exec1Valid ? 6'h19 == writeAddrPRF_exec1Addr | _GEN_6237 : _GEN_6237; // @[decode.scala 784:33]
  wire  _GEN_13062 = writeAddrPRF_exec1Valid ? 6'h1a == writeAddrPRF_exec1Addr | _GEN_6238 : _GEN_6238; // @[decode.scala 784:33]
  wire  _GEN_13063 = writeAddrPRF_exec1Valid ? 6'h1b == writeAddrPRF_exec1Addr | _GEN_6239 : _GEN_6239; // @[decode.scala 784:33]
  wire  _GEN_13064 = writeAddrPRF_exec1Valid ? 6'h1c == writeAddrPRF_exec1Addr | _GEN_6240 : _GEN_6240; // @[decode.scala 784:33]
  wire  _GEN_13065 = writeAddrPRF_exec1Valid ? 6'h1d == writeAddrPRF_exec1Addr | _GEN_6241 : _GEN_6241; // @[decode.scala 784:33]
  wire  _GEN_13066 = writeAddrPRF_exec1Valid ? 6'h1e == writeAddrPRF_exec1Addr | _GEN_6242 : _GEN_6242; // @[decode.scala 784:33]
  wire  _GEN_13067 = writeAddrPRF_exec1Valid ? 6'h1f == writeAddrPRF_exec1Addr | _GEN_6243 : _GEN_6243; // @[decode.scala 784:33]
  wire  _GEN_13068 = writeAddrPRF_exec1Valid ? 6'h20 == writeAddrPRF_exec1Addr | _GEN_6244 : _GEN_6244; // @[decode.scala 784:33]
  wire  _GEN_13069 = writeAddrPRF_exec1Valid ? 6'h21 == writeAddrPRF_exec1Addr | _GEN_6245 : _GEN_6245; // @[decode.scala 784:33]
  wire  _GEN_13070 = writeAddrPRF_exec1Valid ? 6'h22 == writeAddrPRF_exec1Addr | _GEN_6246 : _GEN_6246; // @[decode.scala 784:33]
  wire  _GEN_13071 = writeAddrPRF_exec1Valid ? 6'h23 == writeAddrPRF_exec1Addr | _GEN_6247 : _GEN_6247; // @[decode.scala 784:33]
  wire  _GEN_13072 = writeAddrPRF_exec1Valid ? 6'h24 == writeAddrPRF_exec1Addr | _GEN_6248 : _GEN_6248; // @[decode.scala 784:33]
  wire  _GEN_13073 = writeAddrPRF_exec1Valid ? 6'h25 == writeAddrPRF_exec1Addr | _GEN_6249 : _GEN_6249; // @[decode.scala 784:33]
  wire  _GEN_13074 = writeAddrPRF_exec1Valid ? 6'h26 == writeAddrPRF_exec1Addr | _GEN_6250 : _GEN_6250; // @[decode.scala 784:33]
  wire  _GEN_13075 = writeAddrPRF_exec1Valid ? 6'h27 == writeAddrPRF_exec1Addr | _GEN_6251 : _GEN_6251; // @[decode.scala 784:33]
  wire  _GEN_13076 = writeAddrPRF_exec1Valid ? 6'h28 == writeAddrPRF_exec1Addr | _GEN_6252 : _GEN_6252; // @[decode.scala 784:33]
  wire  _GEN_13077 = writeAddrPRF_exec1Valid ? 6'h29 == writeAddrPRF_exec1Addr | _GEN_6253 : _GEN_6253; // @[decode.scala 784:33]
  wire  _GEN_13078 = writeAddrPRF_exec1Valid ? 6'h2a == writeAddrPRF_exec1Addr | _GEN_6254 : _GEN_6254; // @[decode.scala 784:33]
  wire  _GEN_13079 = writeAddrPRF_exec1Valid ? 6'h2b == writeAddrPRF_exec1Addr | _GEN_6255 : _GEN_6255; // @[decode.scala 784:33]
  wire  _GEN_13080 = writeAddrPRF_exec1Valid ? 6'h2c == writeAddrPRF_exec1Addr | _GEN_6256 : _GEN_6256; // @[decode.scala 784:33]
  wire  _GEN_13081 = writeAddrPRF_exec1Valid ? 6'h2d == writeAddrPRF_exec1Addr | _GEN_6257 : _GEN_6257; // @[decode.scala 784:33]
  wire  _GEN_13082 = writeAddrPRF_exec1Valid ? 6'h2e == writeAddrPRF_exec1Addr | _GEN_6258 : _GEN_6258; // @[decode.scala 784:33]
  wire  _GEN_13083 = writeAddrPRF_exec1Valid ? 6'h2f == writeAddrPRF_exec1Addr | _GEN_6259 : _GEN_6259; // @[decode.scala 784:33]
  wire  _GEN_13084 = writeAddrPRF_exec1Valid ? 6'h30 == writeAddrPRF_exec1Addr | _GEN_6260 : _GEN_6260; // @[decode.scala 784:33]
  wire  _GEN_13085 = writeAddrPRF_exec1Valid ? 6'h31 == writeAddrPRF_exec1Addr | _GEN_6261 : _GEN_6261; // @[decode.scala 784:33]
  wire  _GEN_13086 = writeAddrPRF_exec1Valid ? 6'h32 == writeAddrPRF_exec1Addr | _GEN_6262 : _GEN_6262; // @[decode.scala 784:33]
  wire  _GEN_13087 = writeAddrPRF_exec1Valid ? 6'h33 == writeAddrPRF_exec1Addr | _GEN_6263 : _GEN_6263; // @[decode.scala 784:33]
  wire  _GEN_13088 = writeAddrPRF_exec1Valid ? 6'h34 == writeAddrPRF_exec1Addr | _GEN_6264 : _GEN_6264; // @[decode.scala 784:33]
  wire  _GEN_13089 = writeAddrPRF_exec1Valid ? 6'h35 == writeAddrPRF_exec1Addr | _GEN_6265 : _GEN_6265; // @[decode.scala 784:33]
  wire  _GEN_13090 = writeAddrPRF_exec1Valid ? 6'h36 == writeAddrPRF_exec1Addr | _GEN_6266 : _GEN_6266; // @[decode.scala 784:33]
  wire  _GEN_13091 = writeAddrPRF_exec1Valid ? 6'h37 == writeAddrPRF_exec1Addr | _GEN_6267 : _GEN_6267; // @[decode.scala 784:33]
  wire  _GEN_13092 = writeAddrPRF_exec1Valid ? 6'h38 == writeAddrPRF_exec1Addr | _GEN_6268 : _GEN_6268; // @[decode.scala 784:33]
  wire  _GEN_13093 = writeAddrPRF_exec1Valid ? 6'h39 == writeAddrPRF_exec1Addr | _GEN_6269 : _GEN_6269; // @[decode.scala 784:33]
  wire  _GEN_13094 = writeAddrPRF_exec1Valid ? 6'h3a == writeAddrPRF_exec1Addr | _GEN_6270 : _GEN_6270; // @[decode.scala 784:33]
  wire  _GEN_13095 = writeAddrPRF_exec1Valid ? 6'h3b == writeAddrPRF_exec1Addr | _GEN_6271 : _GEN_6271; // @[decode.scala 784:33]
  wire  _GEN_13096 = writeAddrPRF_exec1Valid ? 6'h3c == writeAddrPRF_exec1Addr | _GEN_6272 : _GEN_6272; // @[decode.scala 784:33]
  wire  _GEN_13097 = writeAddrPRF_exec1Valid ? 6'h3d == writeAddrPRF_exec1Addr | _GEN_6273 : _GEN_6273; // @[decode.scala 784:33]
  wire  _GEN_13098 = writeAddrPRF_exec1Valid ? 6'h3e == writeAddrPRF_exec1Addr | _GEN_6274 : _GEN_6274; // @[decode.scala 784:33]
  wire  _GEN_13099 = writeAddrPRF_exec1Valid ? 6'h3f == writeAddrPRF_exec1Addr | _GEN_6275 : _GEN_6275; // @[decode.scala 784:33]
  wire  _GEN_13164 = writeAddrPRF_exec2Valid ? 6'h0 == writeAddrPRF_exec2Addr | _GEN_13036 : _GEN_13036; // @[decode.scala 785:33]
  wire  _GEN_13165 = writeAddrPRF_exec2Valid ? 6'h1 == writeAddrPRF_exec2Addr | _GEN_13037 : _GEN_13037; // @[decode.scala 785:33]
  wire  _GEN_13166 = writeAddrPRF_exec2Valid ? 6'h2 == writeAddrPRF_exec2Addr | _GEN_13038 : _GEN_13038; // @[decode.scala 785:33]
  wire  _GEN_13167 = writeAddrPRF_exec2Valid ? 6'h3 == writeAddrPRF_exec2Addr | _GEN_13039 : _GEN_13039; // @[decode.scala 785:33]
  wire  _GEN_13168 = writeAddrPRF_exec2Valid ? 6'h4 == writeAddrPRF_exec2Addr | _GEN_13040 : _GEN_13040; // @[decode.scala 785:33]
  wire  _GEN_13169 = writeAddrPRF_exec2Valid ? 6'h5 == writeAddrPRF_exec2Addr | _GEN_13041 : _GEN_13041; // @[decode.scala 785:33]
  wire  _GEN_13170 = writeAddrPRF_exec2Valid ? 6'h6 == writeAddrPRF_exec2Addr | _GEN_13042 : _GEN_13042; // @[decode.scala 785:33]
  wire  _GEN_13171 = writeAddrPRF_exec2Valid ? 6'h7 == writeAddrPRF_exec2Addr | _GEN_13043 : _GEN_13043; // @[decode.scala 785:33]
  wire  _GEN_13172 = writeAddrPRF_exec2Valid ? 6'h8 == writeAddrPRF_exec2Addr | _GEN_13044 : _GEN_13044; // @[decode.scala 785:33]
  wire  _GEN_13173 = writeAddrPRF_exec2Valid ? 6'h9 == writeAddrPRF_exec2Addr | _GEN_13045 : _GEN_13045; // @[decode.scala 785:33]
  wire  _GEN_13174 = writeAddrPRF_exec2Valid ? 6'ha == writeAddrPRF_exec2Addr | _GEN_13046 : _GEN_13046; // @[decode.scala 785:33]
  wire  _GEN_13175 = writeAddrPRF_exec2Valid ? 6'hb == writeAddrPRF_exec2Addr | _GEN_13047 : _GEN_13047; // @[decode.scala 785:33]
  wire  _GEN_13176 = writeAddrPRF_exec2Valid ? 6'hc == writeAddrPRF_exec2Addr | _GEN_13048 : _GEN_13048; // @[decode.scala 785:33]
  wire  _GEN_13177 = writeAddrPRF_exec2Valid ? 6'hd == writeAddrPRF_exec2Addr | _GEN_13049 : _GEN_13049; // @[decode.scala 785:33]
  wire  _GEN_13178 = writeAddrPRF_exec2Valid ? 6'he == writeAddrPRF_exec2Addr | _GEN_13050 : _GEN_13050; // @[decode.scala 785:33]
  wire  _GEN_13179 = writeAddrPRF_exec2Valid ? 6'hf == writeAddrPRF_exec2Addr | _GEN_13051 : _GEN_13051; // @[decode.scala 785:33]
  wire  _GEN_13180 = writeAddrPRF_exec2Valid ? 6'h10 == writeAddrPRF_exec2Addr | _GEN_13052 : _GEN_13052; // @[decode.scala 785:33]
  wire  _GEN_13181 = writeAddrPRF_exec2Valid ? 6'h11 == writeAddrPRF_exec2Addr | _GEN_13053 : _GEN_13053; // @[decode.scala 785:33]
  wire  _GEN_13182 = writeAddrPRF_exec2Valid ? 6'h12 == writeAddrPRF_exec2Addr | _GEN_13054 : _GEN_13054; // @[decode.scala 785:33]
  wire  _GEN_13183 = writeAddrPRF_exec2Valid ? 6'h13 == writeAddrPRF_exec2Addr | _GEN_13055 : _GEN_13055; // @[decode.scala 785:33]
  wire  _GEN_13184 = writeAddrPRF_exec2Valid ? 6'h14 == writeAddrPRF_exec2Addr | _GEN_13056 : _GEN_13056; // @[decode.scala 785:33]
  wire  _GEN_13185 = writeAddrPRF_exec2Valid ? 6'h15 == writeAddrPRF_exec2Addr | _GEN_13057 : _GEN_13057; // @[decode.scala 785:33]
  wire  _GEN_13186 = writeAddrPRF_exec2Valid ? 6'h16 == writeAddrPRF_exec2Addr | _GEN_13058 : _GEN_13058; // @[decode.scala 785:33]
  wire  _GEN_13187 = writeAddrPRF_exec2Valid ? 6'h17 == writeAddrPRF_exec2Addr | _GEN_13059 : _GEN_13059; // @[decode.scala 785:33]
  wire  _GEN_13188 = writeAddrPRF_exec2Valid ? 6'h18 == writeAddrPRF_exec2Addr | _GEN_13060 : _GEN_13060; // @[decode.scala 785:33]
  wire  _GEN_13189 = writeAddrPRF_exec2Valid ? 6'h19 == writeAddrPRF_exec2Addr | _GEN_13061 : _GEN_13061; // @[decode.scala 785:33]
  wire  _GEN_13190 = writeAddrPRF_exec2Valid ? 6'h1a == writeAddrPRF_exec2Addr | _GEN_13062 : _GEN_13062; // @[decode.scala 785:33]
  wire  _GEN_13191 = writeAddrPRF_exec2Valid ? 6'h1b == writeAddrPRF_exec2Addr | _GEN_13063 : _GEN_13063; // @[decode.scala 785:33]
  wire  _GEN_13192 = writeAddrPRF_exec2Valid ? 6'h1c == writeAddrPRF_exec2Addr | _GEN_13064 : _GEN_13064; // @[decode.scala 785:33]
  wire  _GEN_13193 = writeAddrPRF_exec2Valid ? 6'h1d == writeAddrPRF_exec2Addr | _GEN_13065 : _GEN_13065; // @[decode.scala 785:33]
  wire  _GEN_13194 = writeAddrPRF_exec2Valid ? 6'h1e == writeAddrPRF_exec2Addr | _GEN_13066 : _GEN_13066; // @[decode.scala 785:33]
  wire  _GEN_13195 = writeAddrPRF_exec2Valid ? 6'h1f == writeAddrPRF_exec2Addr | _GEN_13067 : _GEN_13067; // @[decode.scala 785:33]
  wire  _GEN_13196 = writeAddrPRF_exec2Valid ? 6'h20 == writeAddrPRF_exec2Addr | _GEN_13068 : _GEN_13068; // @[decode.scala 785:33]
  wire  _GEN_13197 = writeAddrPRF_exec2Valid ? 6'h21 == writeAddrPRF_exec2Addr | _GEN_13069 : _GEN_13069; // @[decode.scala 785:33]
  wire  _GEN_13198 = writeAddrPRF_exec2Valid ? 6'h22 == writeAddrPRF_exec2Addr | _GEN_13070 : _GEN_13070; // @[decode.scala 785:33]
  wire  _GEN_13199 = writeAddrPRF_exec2Valid ? 6'h23 == writeAddrPRF_exec2Addr | _GEN_13071 : _GEN_13071; // @[decode.scala 785:33]
  wire  _GEN_13200 = writeAddrPRF_exec2Valid ? 6'h24 == writeAddrPRF_exec2Addr | _GEN_13072 : _GEN_13072; // @[decode.scala 785:33]
  wire  _GEN_13201 = writeAddrPRF_exec2Valid ? 6'h25 == writeAddrPRF_exec2Addr | _GEN_13073 : _GEN_13073; // @[decode.scala 785:33]
  wire  _GEN_13202 = writeAddrPRF_exec2Valid ? 6'h26 == writeAddrPRF_exec2Addr | _GEN_13074 : _GEN_13074; // @[decode.scala 785:33]
  wire  _GEN_13203 = writeAddrPRF_exec2Valid ? 6'h27 == writeAddrPRF_exec2Addr | _GEN_13075 : _GEN_13075; // @[decode.scala 785:33]
  wire  _GEN_13204 = writeAddrPRF_exec2Valid ? 6'h28 == writeAddrPRF_exec2Addr | _GEN_13076 : _GEN_13076; // @[decode.scala 785:33]
  wire  _GEN_13205 = writeAddrPRF_exec2Valid ? 6'h29 == writeAddrPRF_exec2Addr | _GEN_13077 : _GEN_13077; // @[decode.scala 785:33]
  wire  _GEN_13206 = writeAddrPRF_exec2Valid ? 6'h2a == writeAddrPRF_exec2Addr | _GEN_13078 : _GEN_13078; // @[decode.scala 785:33]
  wire  _GEN_13207 = writeAddrPRF_exec2Valid ? 6'h2b == writeAddrPRF_exec2Addr | _GEN_13079 : _GEN_13079; // @[decode.scala 785:33]
  wire  _GEN_13208 = writeAddrPRF_exec2Valid ? 6'h2c == writeAddrPRF_exec2Addr | _GEN_13080 : _GEN_13080; // @[decode.scala 785:33]
  wire  _GEN_13209 = writeAddrPRF_exec2Valid ? 6'h2d == writeAddrPRF_exec2Addr | _GEN_13081 : _GEN_13081; // @[decode.scala 785:33]
  wire  _GEN_13210 = writeAddrPRF_exec2Valid ? 6'h2e == writeAddrPRF_exec2Addr | _GEN_13082 : _GEN_13082; // @[decode.scala 785:33]
  wire  _GEN_13211 = writeAddrPRF_exec2Valid ? 6'h2f == writeAddrPRF_exec2Addr | _GEN_13083 : _GEN_13083; // @[decode.scala 785:33]
  wire  _GEN_13212 = writeAddrPRF_exec2Valid ? 6'h30 == writeAddrPRF_exec2Addr | _GEN_13084 : _GEN_13084; // @[decode.scala 785:33]
  wire  _GEN_13213 = writeAddrPRF_exec2Valid ? 6'h31 == writeAddrPRF_exec2Addr | _GEN_13085 : _GEN_13085; // @[decode.scala 785:33]
  wire  _GEN_13214 = writeAddrPRF_exec2Valid ? 6'h32 == writeAddrPRF_exec2Addr | _GEN_13086 : _GEN_13086; // @[decode.scala 785:33]
  wire  _GEN_13215 = writeAddrPRF_exec2Valid ? 6'h33 == writeAddrPRF_exec2Addr | _GEN_13087 : _GEN_13087; // @[decode.scala 785:33]
  wire  _GEN_13216 = writeAddrPRF_exec2Valid ? 6'h34 == writeAddrPRF_exec2Addr | _GEN_13088 : _GEN_13088; // @[decode.scala 785:33]
  wire  _GEN_13217 = writeAddrPRF_exec2Valid ? 6'h35 == writeAddrPRF_exec2Addr | _GEN_13089 : _GEN_13089; // @[decode.scala 785:33]
  wire  _GEN_13218 = writeAddrPRF_exec2Valid ? 6'h36 == writeAddrPRF_exec2Addr | _GEN_13090 : _GEN_13090; // @[decode.scala 785:33]
  wire  _GEN_13219 = writeAddrPRF_exec2Valid ? 6'h37 == writeAddrPRF_exec2Addr | _GEN_13091 : _GEN_13091; // @[decode.scala 785:33]
  wire  _GEN_13220 = writeAddrPRF_exec2Valid ? 6'h38 == writeAddrPRF_exec2Addr | _GEN_13092 : _GEN_13092; // @[decode.scala 785:33]
  wire  _GEN_13221 = writeAddrPRF_exec2Valid ? 6'h39 == writeAddrPRF_exec2Addr | _GEN_13093 : _GEN_13093; // @[decode.scala 785:33]
  wire  _GEN_13222 = writeAddrPRF_exec2Valid ? 6'h3a == writeAddrPRF_exec2Addr | _GEN_13094 : _GEN_13094; // @[decode.scala 785:33]
  wire  _GEN_13223 = writeAddrPRF_exec2Valid ? 6'h3b == writeAddrPRF_exec2Addr | _GEN_13095 : _GEN_13095; // @[decode.scala 785:33]
  wire  _GEN_13224 = writeAddrPRF_exec2Valid ? 6'h3c == writeAddrPRF_exec2Addr | _GEN_13096 : _GEN_13096; // @[decode.scala 785:33]
  wire  _GEN_13225 = writeAddrPRF_exec2Valid ? 6'h3d == writeAddrPRF_exec2Addr | _GEN_13097 : _GEN_13097; // @[decode.scala 785:33]
  wire  _GEN_13226 = writeAddrPRF_exec2Valid ? 6'h3e == writeAddrPRF_exec2Addr | _GEN_13098 : _GEN_13098; // @[decode.scala 785:33]
  wire  _GEN_13227 = writeAddrPRF_exec2Valid ? 6'h3f == writeAddrPRF_exec2Addr | _GEN_13099 : _GEN_13099; // @[decode.scala 785:33]
  wire  _GEN_13292 = writeAddrPRF_exec3Valid ? 6'h0 == writeAddrPRF_exec3Addr | _GEN_13164 : _GEN_13164; // @[decode.scala 786:33]
  wire  _GEN_13293 = writeAddrPRF_exec3Valid ? 6'h1 == writeAddrPRF_exec3Addr | _GEN_13165 : _GEN_13165; // @[decode.scala 786:33]
  wire  _GEN_13294 = writeAddrPRF_exec3Valid ? 6'h2 == writeAddrPRF_exec3Addr | _GEN_13166 : _GEN_13166; // @[decode.scala 786:33]
  wire  _GEN_13295 = writeAddrPRF_exec3Valid ? 6'h3 == writeAddrPRF_exec3Addr | _GEN_13167 : _GEN_13167; // @[decode.scala 786:33]
  wire  _GEN_13296 = writeAddrPRF_exec3Valid ? 6'h4 == writeAddrPRF_exec3Addr | _GEN_13168 : _GEN_13168; // @[decode.scala 786:33]
  wire  _GEN_13297 = writeAddrPRF_exec3Valid ? 6'h5 == writeAddrPRF_exec3Addr | _GEN_13169 : _GEN_13169; // @[decode.scala 786:33]
  wire  _GEN_13298 = writeAddrPRF_exec3Valid ? 6'h6 == writeAddrPRF_exec3Addr | _GEN_13170 : _GEN_13170; // @[decode.scala 786:33]
  wire  _GEN_13299 = writeAddrPRF_exec3Valid ? 6'h7 == writeAddrPRF_exec3Addr | _GEN_13171 : _GEN_13171; // @[decode.scala 786:33]
  wire  _GEN_13300 = writeAddrPRF_exec3Valid ? 6'h8 == writeAddrPRF_exec3Addr | _GEN_13172 : _GEN_13172; // @[decode.scala 786:33]
  wire  _GEN_13301 = writeAddrPRF_exec3Valid ? 6'h9 == writeAddrPRF_exec3Addr | _GEN_13173 : _GEN_13173; // @[decode.scala 786:33]
  wire  _GEN_13302 = writeAddrPRF_exec3Valid ? 6'ha == writeAddrPRF_exec3Addr | _GEN_13174 : _GEN_13174; // @[decode.scala 786:33]
  wire  _GEN_13303 = writeAddrPRF_exec3Valid ? 6'hb == writeAddrPRF_exec3Addr | _GEN_13175 : _GEN_13175; // @[decode.scala 786:33]
  wire  _GEN_13304 = writeAddrPRF_exec3Valid ? 6'hc == writeAddrPRF_exec3Addr | _GEN_13176 : _GEN_13176; // @[decode.scala 786:33]
  wire  _GEN_13305 = writeAddrPRF_exec3Valid ? 6'hd == writeAddrPRF_exec3Addr | _GEN_13177 : _GEN_13177; // @[decode.scala 786:33]
  wire  _GEN_13306 = writeAddrPRF_exec3Valid ? 6'he == writeAddrPRF_exec3Addr | _GEN_13178 : _GEN_13178; // @[decode.scala 786:33]
  wire  _GEN_13307 = writeAddrPRF_exec3Valid ? 6'hf == writeAddrPRF_exec3Addr | _GEN_13179 : _GEN_13179; // @[decode.scala 786:33]
  wire  _GEN_13308 = writeAddrPRF_exec3Valid ? 6'h10 == writeAddrPRF_exec3Addr | _GEN_13180 : _GEN_13180; // @[decode.scala 786:33]
  wire  _GEN_13309 = writeAddrPRF_exec3Valid ? 6'h11 == writeAddrPRF_exec3Addr | _GEN_13181 : _GEN_13181; // @[decode.scala 786:33]
  wire  _GEN_13310 = writeAddrPRF_exec3Valid ? 6'h12 == writeAddrPRF_exec3Addr | _GEN_13182 : _GEN_13182; // @[decode.scala 786:33]
  wire  _GEN_13311 = writeAddrPRF_exec3Valid ? 6'h13 == writeAddrPRF_exec3Addr | _GEN_13183 : _GEN_13183; // @[decode.scala 786:33]
  wire  _GEN_13312 = writeAddrPRF_exec3Valid ? 6'h14 == writeAddrPRF_exec3Addr | _GEN_13184 : _GEN_13184; // @[decode.scala 786:33]
  wire  _GEN_13313 = writeAddrPRF_exec3Valid ? 6'h15 == writeAddrPRF_exec3Addr | _GEN_13185 : _GEN_13185; // @[decode.scala 786:33]
  wire  _GEN_13314 = writeAddrPRF_exec3Valid ? 6'h16 == writeAddrPRF_exec3Addr | _GEN_13186 : _GEN_13186; // @[decode.scala 786:33]
  wire  _GEN_13315 = writeAddrPRF_exec3Valid ? 6'h17 == writeAddrPRF_exec3Addr | _GEN_13187 : _GEN_13187; // @[decode.scala 786:33]
  wire  _GEN_13316 = writeAddrPRF_exec3Valid ? 6'h18 == writeAddrPRF_exec3Addr | _GEN_13188 : _GEN_13188; // @[decode.scala 786:33]
  wire  _GEN_13317 = writeAddrPRF_exec3Valid ? 6'h19 == writeAddrPRF_exec3Addr | _GEN_13189 : _GEN_13189; // @[decode.scala 786:33]
  wire  _GEN_13318 = writeAddrPRF_exec3Valid ? 6'h1a == writeAddrPRF_exec3Addr | _GEN_13190 : _GEN_13190; // @[decode.scala 786:33]
  wire  _GEN_13319 = writeAddrPRF_exec3Valid ? 6'h1b == writeAddrPRF_exec3Addr | _GEN_13191 : _GEN_13191; // @[decode.scala 786:33]
  wire  _GEN_13320 = writeAddrPRF_exec3Valid ? 6'h1c == writeAddrPRF_exec3Addr | _GEN_13192 : _GEN_13192; // @[decode.scala 786:33]
  wire  _GEN_13321 = writeAddrPRF_exec3Valid ? 6'h1d == writeAddrPRF_exec3Addr | _GEN_13193 : _GEN_13193; // @[decode.scala 786:33]
  wire  _GEN_13322 = writeAddrPRF_exec3Valid ? 6'h1e == writeAddrPRF_exec3Addr | _GEN_13194 : _GEN_13194; // @[decode.scala 786:33]
  wire  _GEN_13323 = writeAddrPRF_exec3Valid ? 6'h1f == writeAddrPRF_exec3Addr | _GEN_13195 : _GEN_13195; // @[decode.scala 786:33]
  wire  _GEN_13356 = _T_222 | stateRegInputBuf; // @[decode.scala 804:58 805:32 193:34]
  wire  _GEN_13357 = fromFetch_expected_valid ? _GEN_13356 : 1'h1; // @[decode.scala 803:42 808:30]
  wire  _GEN_13362 = branchEvalIn_fired & ~branchEvalIn_passFail ? 1'h0 : _GEN_10979; // @[decode.scala 794:58 798:18]
  wire  _GEN_13364 = ~fromFetch_fired | _T_224 & fun3 == 3'h0 & immediate_immediate == 64'h302 ? 1'h0 : stateRegInputBuf
    ; // @[decode.scala 827:100 828:32 193:34]
  wire  _GEN_13366 = readyOutputBuf ? _GEN_13364 : stateRegInputBuf; // @[decode.scala 825:32 193:34]
  wire  _GEN_13369 = ~stall & ~(branchEvalIn_fired & (opcode == 7'h63 | opcode == 7'h6f | opcode == 7'h67)) ? _GEN_13366
     : stateRegInputBuf; // @[decode.scala 823:114 193:34]
  wire  _GEN_13383 = validInputBuf | stateRegOutputBuf; // @[decode.scala 855:29 856:29 194:34]
  wire  _GEN_13387 = ~validInputBuf ? 1'h0 : stateRegOutputBuf; // @[decode.scala 869:32 870:31 194:34]
  wire  _GEN_13389 = toExec_fired ? _GEN_13387 : stateRegOutputBuf; // @[decode.scala 867:28 194:34]
  wire  _T_466 = writeBackResult_instruction[6:0] != 7'h63; // @[decode.scala 885:38]
  wire  _T_467 = writeBackResult_fired & writeBackResult_rdAddr != 5'h0 & _T_466; // @[decode.scala 884:61]
  wire  _T_469 = writeBackResult_instruction[6:0] != 7'h23; // @[decode.scala 886:38]
  wire  _T_470 = _T_467 & _T_469; // @[decode.scala 885:50]
  wire [5:0] _GEN_13400 = 5'h1 == writeBackResult_rdAddr ? architecturalRegMap_1 : architecturalRegMap_0; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13401 = 5'h2 == writeBackResult_rdAddr ? architecturalRegMap_2 : _GEN_13400; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13402 = 5'h3 == writeBackResult_rdAddr ? architecturalRegMap_3 : _GEN_13401; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13403 = 5'h4 == writeBackResult_rdAddr ? architecturalRegMap_4 : _GEN_13402; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13404 = 5'h5 == writeBackResult_rdAddr ? architecturalRegMap_5 : _GEN_13403; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13405 = 5'h6 == writeBackResult_rdAddr ? architecturalRegMap_6 : _GEN_13404; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13406 = 5'h7 == writeBackResult_rdAddr ? architecturalRegMap_7 : _GEN_13405; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13407 = 5'h8 == writeBackResult_rdAddr ? architecturalRegMap_8 : _GEN_13406; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13408 = 5'h9 == writeBackResult_rdAddr ? architecturalRegMap_9 : _GEN_13407; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13409 = 5'ha == writeBackResult_rdAddr ? architecturalRegMap_10 : _GEN_13408; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13410 = 5'hb == writeBackResult_rdAddr ? architecturalRegMap_11 : _GEN_13409; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13411 = 5'hc == writeBackResult_rdAddr ? architecturalRegMap_12 : _GEN_13410; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13412 = 5'hd == writeBackResult_rdAddr ? architecturalRegMap_13 : _GEN_13411; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13413 = 5'he == writeBackResult_rdAddr ? architecturalRegMap_14 : _GEN_13412; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13414 = 5'hf == writeBackResult_rdAddr ? architecturalRegMap_15 : _GEN_13413; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13415 = 5'h10 == writeBackResult_rdAddr ? architecturalRegMap_16 : _GEN_13414; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13416 = 5'h11 == writeBackResult_rdAddr ? architecturalRegMap_17 : _GEN_13415; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13417 = 5'h12 == writeBackResult_rdAddr ? architecturalRegMap_18 : _GEN_13416; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13418 = 5'h13 == writeBackResult_rdAddr ? architecturalRegMap_19 : _GEN_13417; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13419 = 5'h14 == writeBackResult_rdAddr ? architecturalRegMap_20 : _GEN_13418; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13420 = 5'h15 == writeBackResult_rdAddr ? architecturalRegMap_21 : _GEN_13419; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13421 = 5'h16 == writeBackResult_rdAddr ? architecturalRegMap_22 : _GEN_13420; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13422 = 5'h17 == writeBackResult_rdAddr ? architecturalRegMap_23 : _GEN_13421; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13423 = 5'h18 == writeBackResult_rdAddr ? architecturalRegMap_24 : _GEN_13422; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13424 = 5'h19 == writeBackResult_rdAddr ? architecturalRegMap_25 : _GEN_13423; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13425 = 5'h1a == writeBackResult_rdAddr ? architecturalRegMap_26 : _GEN_13424; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13426 = 5'h1b == writeBackResult_rdAddr ? architecturalRegMap_27 : _GEN_13425; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13427 = 5'h1c == writeBackResult_rdAddr ? architecturalRegMap_28 : _GEN_13426; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13428 = 5'h1d == writeBackResult_rdAddr ? architecturalRegMap_29 : _GEN_13427; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13429 = 5'h1e == writeBackResult_rdAddr ? architecturalRegMap_30 : _GEN_13428; // @[decode.scala 887:{49,49}]
  wire [5:0] _GEN_13430 = 5'h1f == writeBackResult_rdAddr ? architecturalRegMap_31 : _GEN_13429; // @[decode.scala 887:{49,49}]
  wire  _T_471 = _GEN_13430 != writeBackResult_PRFDest; // @[decode.scala 887:49]
  wire  _T_472 = _T_470 & _T_471; // @[decode.scala 886:50]
  wire  _T_473 = writeBackResult_instruction != 32'h80000073; // @[decode.scala 888:33]
  wire  _T_474 = _T_472 & _T_473; // @[decode.scala 887:77]
  wire  _GEN_16294 = 6'h0 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13463 = 6'h0 == _GEN_13430 | _GEN_6148; // @[decode.scala 891:{62,62}]
  wire  _GEN_16295 = 6'h1 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13464 = 6'h1 == _GEN_13430 | _GEN_6149; // @[decode.scala 891:{62,62}]
  wire  _GEN_16296 = 6'h2 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13465 = 6'h2 == _GEN_13430 | _GEN_6150; // @[decode.scala 891:{62,62}]
  wire  _GEN_16297 = 6'h3 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13466 = 6'h3 == _GEN_13430 | _GEN_6151; // @[decode.scala 891:{62,62}]
  wire  _GEN_16298 = 6'h4 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13467 = 6'h4 == _GEN_13430 | _GEN_6152; // @[decode.scala 891:{62,62}]
  wire  _GEN_16299 = 6'h5 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13468 = 6'h5 == _GEN_13430 | _GEN_6153; // @[decode.scala 891:{62,62}]
  wire  _GEN_16300 = 6'h6 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13469 = 6'h6 == _GEN_13430 | _GEN_6154; // @[decode.scala 891:{62,62}]
  wire  _GEN_16301 = 6'h7 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13470 = 6'h7 == _GEN_13430 | _GEN_6155; // @[decode.scala 891:{62,62}]
  wire  _GEN_16302 = 6'h8 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13471 = 6'h8 == _GEN_13430 | _GEN_6156; // @[decode.scala 891:{62,62}]
  wire  _GEN_16303 = 6'h9 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13472 = 6'h9 == _GEN_13430 | _GEN_6157; // @[decode.scala 891:{62,62}]
  wire  _GEN_16304 = 6'ha == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13473 = 6'ha == _GEN_13430 | _GEN_6158; // @[decode.scala 891:{62,62}]
  wire  _GEN_16305 = 6'hb == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13474 = 6'hb == _GEN_13430 | _GEN_6159; // @[decode.scala 891:{62,62}]
  wire  _GEN_16306 = 6'hc == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13475 = 6'hc == _GEN_13430 | _GEN_6160; // @[decode.scala 891:{62,62}]
  wire  _GEN_16307 = 6'hd == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13476 = 6'hd == _GEN_13430 | _GEN_6161; // @[decode.scala 891:{62,62}]
  wire  _GEN_16308 = 6'he == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13477 = 6'he == _GEN_13430 | _GEN_6162; // @[decode.scala 891:{62,62}]
  wire  _GEN_16309 = 6'hf == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13478 = 6'hf == _GEN_13430 | _GEN_6163; // @[decode.scala 891:{62,62}]
  wire  _GEN_16310 = 6'h10 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13479 = 6'h10 == _GEN_13430 | _GEN_6164; // @[decode.scala 891:{62,62}]
  wire  _GEN_16311 = 6'h11 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13480 = 6'h11 == _GEN_13430 | _GEN_6165; // @[decode.scala 891:{62,62}]
  wire  _GEN_16312 = 6'h12 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13481 = 6'h12 == _GEN_13430 | _GEN_6166; // @[decode.scala 891:{62,62}]
  wire  _GEN_16313 = 6'h13 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13482 = 6'h13 == _GEN_13430 | _GEN_6167; // @[decode.scala 891:{62,62}]
  wire  _GEN_16314 = 6'h14 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13483 = 6'h14 == _GEN_13430 | _GEN_6168; // @[decode.scala 891:{62,62}]
  wire  _GEN_16315 = 6'h15 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13484 = 6'h15 == _GEN_13430 | _GEN_6169; // @[decode.scala 891:{62,62}]
  wire  _GEN_16316 = 6'h16 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13485 = 6'h16 == _GEN_13430 | _GEN_6170; // @[decode.scala 891:{62,62}]
  wire  _GEN_16317 = 6'h17 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13486 = 6'h17 == _GEN_13430 | _GEN_6171; // @[decode.scala 891:{62,62}]
  wire  _GEN_16318 = 6'h18 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13487 = 6'h18 == _GEN_13430 | _GEN_6172; // @[decode.scala 891:{62,62}]
  wire  _GEN_16319 = 6'h19 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13488 = 6'h19 == _GEN_13430 | _GEN_6173; // @[decode.scala 891:{62,62}]
  wire  _GEN_16320 = 6'h1a == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13489 = 6'h1a == _GEN_13430 | _GEN_6174; // @[decode.scala 891:{62,62}]
  wire  _GEN_16321 = 6'h1b == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13490 = 6'h1b == _GEN_13430 | _GEN_6175; // @[decode.scala 891:{62,62}]
  wire  _GEN_16322 = 6'h1c == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13491 = 6'h1c == _GEN_13430 | _GEN_6176; // @[decode.scala 891:{62,62}]
  wire  _GEN_16323 = 6'h1d == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13492 = 6'h1d == _GEN_13430 | _GEN_6177; // @[decode.scala 891:{62,62}]
  wire  _GEN_16324 = 6'h1e == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13493 = 6'h1e == _GEN_13430 | _GEN_6178; // @[decode.scala 891:{62,62}]
  wire  _GEN_16325 = 6'h1f == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13494 = 6'h1f == _GEN_13430 | _GEN_6179; // @[decode.scala 891:{62,62}]
  wire  _GEN_16326 = 6'h20 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13495 = 6'h20 == _GEN_13430 | _GEN_6180; // @[decode.scala 891:{62,62}]
  wire  _GEN_16327 = 6'h21 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13496 = 6'h21 == _GEN_13430 | _GEN_6181; // @[decode.scala 891:{62,62}]
  wire  _GEN_16328 = 6'h22 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13497 = 6'h22 == _GEN_13430 | _GEN_6182; // @[decode.scala 891:{62,62}]
  wire  _GEN_16329 = 6'h23 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13498 = 6'h23 == _GEN_13430 | _GEN_6183; // @[decode.scala 891:{62,62}]
  wire  _GEN_16330 = 6'h24 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13499 = 6'h24 == _GEN_13430 | _GEN_6184; // @[decode.scala 891:{62,62}]
  wire  _GEN_16331 = 6'h25 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13500 = 6'h25 == _GEN_13430 | _GEN_6185; // @[decode.scala 891:{62,62}]
  wire  _GEN_16332 = 6'h26 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13501 = 6'h26 == _GEN_13430 | _GEN_6186; // @[decode.scala 891:{62,62}]
  wire  _GEN_16333 = 6'h27 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13502 = 6'h27 == _GEN_13430 | _GEN_6187; // @[decode.scala 891:{62,62}]
  wire  _GEN_16334 = 6'h28 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13503 = 6'h28 == _GEN_13430 | _GEN_6188; // @[decode.scala 891:{62,62}]
  wire  _GEN_16335 = 6'h29 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13504 = 6'h29 == _GEN_13430 | _GEN_6189; // @[decode.scala 891:{62,62}]
  wire  _GEN_16336 = 6'h2a == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13505 = 6'h2a == _GEN_13430 | _GEN_6190; // @[decode.scala 891:{62,62}]
  wire  _GEN_16337 = 6'h2b == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13506 = 6'h2b == _GEN_13430 | _GEN_6191; // @[decode.scala 891:{62,62}]
  wire  _GEN_16338 = 6'h2c == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13507 = 6'h2c == _GEN_13430 | _GEN_6192; // @[decode.scala 891:{62,62}]
  wire  _GEN_16339 = 6'h2d == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13508 = 6'h2d == _GEN_13430 | _GEN_6193; // @[decode.scala 891:{62,62}]
  wire  _GEN_16340 = 6'h2e == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13509 = 6'h2e == _GEN_13430 | _GEN_6194; // @[decode.scala 891:{62,62}]
  wire  _GEN_16341 = 6'h2f == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13510 = 6'h2f == _GEN_13430 | _GEN_6195; // @[decode.scala 891:{62,62}]
  wire  _GEN_16342 = 6'h30 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13511 = 6'h30 == _GEN_13430 | _GEN_6196; // @[decode.scala 891:{62,62}]
  wire  _GEN_16343 = 6'h31 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13512 = 6'h31 == _GEN_13430 | _GEN_6197; // @[decode.scala 891:{62,62}]
  wire  _GEN_16344 = 6'h32 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13513 = 6'h32 == _GEN_13430 | _GEN_6198; // @[decode.scala 891:{62,62}]
  wire  _GEN_16345 = 6'h33 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13514 = 6'h33 == _GEN_13430 | _GEN_6199; // @[decode.scala 891:{62,62}]
  wire  _GEN_16346 = 6'h34 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13515 = 6'h34 == _GEN_13430 | _GEN_6200; // @[decode.scala 891:{62,62}]
  wire  _GEN_16347 = 6'h35 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13516 = 6'h35 == _GEN_13430 | _GEN_6201; // @[decode.scala 891:{62,62}]
  wire  _GEN_16348 = 6'h36 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13517 = 6'h36 == _GEN_13430 | _GEN_6202; // @[decode.scala 891:{62,62}]
  wire  _GEN_16349 = 6'h37 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13518 = 6'h37 == _GEN_13430 | _GEN_6203; // @[decode.scala 891:{62,62}]
  wire  _GEN_16350 = 6'h38 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13519 = 6'h38 == _GEN_13430 | _GEN_6204; // @[decode.scala 891:{62,62}]
  wire  _GEN_16351 = 6'h39 == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13520 = 6'h39 == _GEN_13430 | _GEN_6205; // @[decode.scala 891:{62,62}]
  wire  _GEN_16352 = 6'h3a == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13521 = 6'h3a == _GEN_13430 | _GEN_6206; // @[decode.scala 891:{62,62}]
  wire  _GEN_16353 = 6'h3b == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13522 = 6'h3b == _GEN_13430 | _GEN_6207; // @[decode.scala 891:{62,62}]
  wire  _GEN_16354 = 6'h3c == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13523 = 6'h3c == _GEN_13430 | _GEN_6208; // @[decode.scala 891:{62,62}]
  wire  _GEN_16355 = 6'h3d == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13524 = 6'h3d == _GEN_13430 | _GEN_6209; // @[decode.scala 891:{62,62}]
  wire  _GEN_16356 = 6'h3e == _GEN_13430; // @[decode.scala 891:{62,62}]
  wire  _GEN_13525 = 6'h3e == _GEN_13430 | _GEN_6210; // @[decode.scala 891:{62,62}]
  wire  _GEN_13527 = _GEN_16294 | _GEN_10335; // @[decode.scala 892:{68,68}]
  wire  _GEN_13528 = _GEN_16295 | _GEN_10336; // @[decode.scala 892:{68,68}]
  wire  _GEN_13529 = _GEN_16296 | _GEN_10337; // @[decode.scala 892:{68,68}]
  wire  _GEN_13530 = _GEN_16297 | _GEN_10338; // @[decode.scala 892:{68,68}]
  wire  _GEN_13531 = _GEN_16298 | _GEN_10339; // @[decode.scala 892:{68,68}]
  wire  _GEN_13532 = _GEN_16299 | _GEN_10340; // @[decode.scala 892:{68,68}]
  wire  _GEN_13533 = _GEN_16300 | _GEN_10341; // @[decode.scala 892:{68,68}]
  wire  _GEN_13534 = _GEN_16301 | _GEN_10342; // @[decode.scala 892:{68,68}]
  wire  _GEN_13535 = _GEN_16302 | _GEN_10343; // @[decode.scala 892:{68,68}]
  wire  _GEN_13536 = _GEN_16303 | _GEN_10344; // @[decode.scala 892:{68,68}]
  wire  _GEN_13537 = _GEN_16304 | _GEN_10345; // @[decode.scala 892:{68,68}]
  wire  _GEN_13538 = _GEN_16305 | _GEN_10346; // @[decode.scala 892:{68,68}]
  wire  _GEN_13539 = _GEN_16306 | _GEN_10347; // @[decode.scala 892:{68,68}]
  wire  _GEN_13540 = _GEN_16307 | _GEN_10348; // @[decode.scala 892:{68,68}]
  wire  _GEN_13541 = _GEN_16308 | _GEN_10349; // @[decode.scala 892:{68,68}]
  wire  _GEN_13542 = _GEN_16309 | _GEN_10350; // @[decode.scala 892:{68,68}]
  wire  _GEN_13543 = _GEN_16310 | _GEN_10351; // @[decode.scala 892:{68,68}]
  wire  _GEN_13544 = _GEN_16311 | _GEN_10352; // @[decode.scala 892:{68,68}]
  wire  _GEN_13545 = _GEN_16312 | _GEN_10353; // @[decode.scala 892:{68,68}]
  wire  _GEN_13546 = _GEN_16313 | _GEN_10354; // @[decode.scala 892:{68,68}]
  wire  _GEN_13547 = _GEN_16314 | _GEN_10355; // @[decode.scala 892:{68,68}]
  wire  _GEN_13548 = _GEN_16315 | _GEN_10356; // @[decode.scala 892:{68,68}]
  wire  _GEN_13549 = _GEN_16316 | _GEN_10357; // @[decode.scala 892:{68,68}]
  wire  _GEN_13550 = _GEN_16317 | _GEN_10358; // @[decode.scala 892:{68,68}]
  wire  _GEN_13551 = _GEN_16318 | _GEN_10359; // @[decode.scala 892:{68,68}]
  wire  _GEN_13552 = _GEN_16319 | _GEN_10360; // @[decode.scala 892:{68,68}]
  wire  _GEN_13553 = _GEN_16320 | _GEN_10361; // @[decode.scala 892:{68,68}]
  wire  _GEN_13554 = _GEN_16321 | _GEN_10362; // @[decode.scala 892:{68,68}]
  wire  _GEN_13555 = _GEN_16322 | _GEN_10363; // @[decode.scala 892:{68,68}]
  wire  _GEN_13556 = _GEN_16323 | _GEN_10364; // @[decode.scala 892:{68,68}]
  wire  _GEN_13557 = _GEN_16324 | _GEN_10365; // @[decode.scala 892:{68,68}]
  wire  _GEN_13558 = _GEN_16325 | _GEN_10366; // @[decode.scala 892:{68,68}]
  wire  _GEN_13559 = _GEN_16326 | _GEN_10367; // @[decode.scala 892:{68,68}]
  wire  _GEN_13560 = _GEN_16327 | _GEN_10368; // @[decode.scala 892:{68,68}]
  wire  _GEN_13561 = _GEN_16328 | _GEN_10369; // @[decode.scala 892:{68,68}]
  wire  _GEN_13562 = _GEN_16329 | _GEN_10370; // @[decode.scala 892:{68,68}]
  wire  _GEN_13563 = _GEN_16330 | _GEN_10371; // @[decode.scala 892:{68,68}]
  wire  _GEN_13564 = _GEN_16331 | _GEN_10372; // @[decode.scala 892:{68,68}]
  wire  _GEN_13565 = _GEN_16332 | _GEN_10373; // @[decode.scala 892:{68,68}]
  wire  _GEN_13566 = _GEN_16333 | _GEN_10374; // @[decode.scala 892:{68,68}]
  wire  _GEN_13567 = _GEN_16334 | _GEN_10375; // @[decode.scala 892:{68,68}]
  wire  _GEN_13568 = _GEN_16335 | _GEN_10376; // @[decode.scala 892:{68,68}]
  wire  _GEN_13569 = _GEN_16336 | _GEN_10377; // @[decode.scala 892:{68,68}]
  wire  _GEN_13570 = _GEN_16337 | _GEN_10378; // @[decode.scala 892:{68,68}]
  wire  _GEN_13571 = _GEN_16338 | _GEN_10379; // @[decode.scala 892:{68,68}]
  wire  _GEN_13572 = _GEN_16339 | _GEN_10380; // @[decode.scala 892:{68,68}]
  wire  _GEN_13573 = _GEN_16340 | _GEN_10381; // @[decode.scala 892:{68,68}]
  wire  _GEN_13574 = _GEN_16341 | _GEN_10382; // @[decode.scala 892:{68,68}]
  wire  _GEN_13575 = _GEN_16342 | _GEN_10383; // @[decode.scala 892:{68,68}]
  wire  _GEN_13576 = _GEN_16343 | _GEN_10384; // @[decode.scala 892:{68,68}]
  wire  _GEN_13577 = _GEN_16344 | _GEN_10385; // @[decode.scala 892:{68,68}]
  wire  _GEN_13578 = _GEN_16345 | _GEN_10386; // @[decode.scala 892:{68,68}]
  wire  _GEN_13579 = _GEN_16346 | _GEN_10387; // @[decode.scala 892:{68,68}]
  wire  _GEN_13580 = _GEN_16347 | _GEN_10388; // @[decode.scala 892:{68,68}]
  wire  _GEN_13581 = _GEN_16348 | _GEN_10389; // @[decode.scala 892:{68,68}]
  wire  _GEN_13582 = _GEN_16349 | _GEN_10390; // @[decode.scala 892:{68,68}]
  wire  _GEN_13583 = _GEN_16350 | _GEN_10391; // @[decode.scala 892:{68,68}]
  wire  _GEN_13584 = _GEN_16351 | _GEN_10392; // @[decode.scala 892:{68,68}]
  wire  _GEN_13585 = _GEN_16352 | _GEN_10393; // @[decode.scala 892:{68,68}]
  wire  _GEN_13586 = _GEN_16353 | _GEN_10394; // @[decode.scala 892:{68,68}]
  wire  _GEN_13587 = _GEN_16354 | _GEN_10395; // @[decode.scala 892:{68,68}]
  wire  _GEN_13588 = _GEN_16355 | _GEN_10396; // @[decode.scala 892:{68,68}]
  wire  _GEN_13589 = _GEN_16356 | _GEN_10397; // @[decode.scala 892:{68,68}]
  wire  _GEN_13591 = _GEN_16294 | _GEN_10495; // @[decode.scala 893:{68,68}]
  wire  _GEN_13592 = _GEN_16295 | _GEN_10496; // @[decode.scala 893:{68,68}]
  wire  _GEN_13593 = _GEN_16296 | _GEN_10497; // @[decode.scala 893:{68,68}]
  wire  _GEN_13594 = _GEN_16297 | _GEN_10498; // @[decode.scala 893:{68,68}]
  wire  _GEN_13595 = _GEN_16298 | _GEN_10499; // @[decode.scala 893:{68,68}]
  wire  _GEN_13596 = _GEN_16299 | _GEN_10500; // @[decode.scala 893:{68,68}]
  wire  _GEN_13597 = _GEN_16300 | _GEN_10501; // @[decode.scala 893:{68,68}]
  wire  _GEN_13598 = _GEN_16301 | _GEN_10502; // @[decode.scala 893:{68,68}]
  wire  _GEN_13599 = _GEN_16302 | _GEN_10503; // @[decode.scala 893:{68,68}]
  wire  _GEN_13600 = _GEN_16303 | _GEN_10504; // @[decode.scala 893:{68,68}]
  wire  _GEN_13601 = _GEN_16304 | _GEN_10505; // @[decode.scala 893:{68,68}]
  wire  _GEN_13602 = _GEN_16305 | _GEN_10506; // @[decode.scala 893:{68,68}]
  wire  _GEN_13603 = _GEN_16306 | _GEN_10507; // @[decode.scala 893:{68,68}]
  wire  _GEN_13604 = _GEN_16307 | _GEN_10508; // @[decode.scala 893:{68,68}]
  wire  _GEN_13605 = _GEN_16308 | _GEN_10509; // @[decode.scala 893:{68,68}]
  wire  _GEN_13606 = _GEN_16309 | _GEN_10510; // @[decode.scala 893:{68,68}]
  wire  _GEN_13607 = _GEN_16310 | _GEN_10511; // @[decode.scala 893:{68,68}]
  wire  _GEN_13608 = _GEN_16311 | _GEN_10512; // @[decode.scala 893:{68,68}]
  wire  _GEN_13609 = _GEN_16312 | _GEN_10513; // @[decode.scala 893:{68,68}]
  wire  _GEN_13610 = _GEN_16313 | _GEN_10514; // @[decode.scala 893:{68,68}]
  wire  _GEN_13611 = _GEN_16314 | _GEN_10515; // @[decode.scala 893:{68,68}]
  wire  _GEN_13612 = _GEN_16315 | _GEN_10516; // @[decode.scala 893:{68,68}]
  wire  _GEN_13613 = _GEN_16316 | _GEN_10517; // @[decode.scala 893:{68,68}]
  wire  _GEN_13614 = _GEN_16317 | _GEN_10518; // @[decode.scala 893:{68,68}]
  wire  _GEN_13615 = _GEN_16318 | _GEN_10519; // @[decode.scala 893:{68,68}]
  wire  _GEN_13616 = _GEN_16319 | _GEN_10520; // @[decode.scala 893:{68,68}]
  wire  _GEN_13617 = _GEN_16320 | _GEN_10521; // @[decode.scala 893:{68,68}]
  wire  _GEN_13618 = _GEN_16321 | _GEN_10522; // @[decode.scala 893:{68,68}]
  wire  _GEN_13619 = _GEN_16322 | _GEN_10523; // @[decode.scala 893:{68,68}]
  wire  _GEN_13620 = _GEN_16323 | _GEN_10524; // @[decode.scala 893:{68,68}]
  wire  _GEN_13621 = _GEN_16324 | _GEN_10525; // @[decode.scala 893:{68,68}]
  wire  _GEN_13622 = _GEN_16325 | _GEN_10526; // @[decode.scala 893:{68,68}]
  wire  _GEN_13623 = _GEN_16326 | _GEN_10527; // @[decode.scala 893:{68,68}]
  wire  _GEN_13624 = _GEN_16327 | _GEN_10528; // @[decode.scala 893:{68,68}]
  wire  _GEN_13625 = _GEN_16328 | _GEN_10529; // @[decode.scala 893:{68,68}]
  wire  _GEN_13626 = _GEN_16329 | _GEN_10530; // @[decode.scala 893:{68,68}]
  wire  _GEN_13627 = _GEN_16330 | _GEN_10531; // @[decode.scala 893:{68,68}]
  wire  _GEN_13628 = _GEN_16331 | _GEN_10532; // @[decode.scala 893:{68,68}]
  wire  _GEN_13629 = _GEN_16332 | _GEN_10533; // @[decode.scala 893:{68,68}]
  wire  _GEN_13630 = _GEN_16333 | _GEN_10534; // @[decode.scala 893:{68,68}]
  wire  _GEN_13631 = _GEN_16334 | _GEN_10535; // @[decode.scala 893:{68,68}]
  wire  _GEN_13632 = _GEN_16335 | _GEN_10536; // @[decode.scala 893:{68,68}]
  wire  _GEN_13633 = _GEN_16336 | _GEN_10537; // @[decode.scala 893:{68,68}]
  wire  _GEN_13634 = _GEN_16337 | _GEN_10538; // @[decode.scala 893:{68,68}]
  wire  _GEN_13635 = _GEN_16338 | _GEN_10539; // @[decode.scala 893:{68,68}]
  wire  _GEN_13636 = _GEN_16339 | _GEN_10540; // @[decode.scala 893:{68,68}]
  wire  _GEN_13637 = _GEN_16340 | _GEN_10541; // @[decode.scala 893:{68,68}]
  wire  _GEN_13638 = _GEN_16341 | _GEN_10542; // @[decode.scala 893:{68,68}]
  wire  _GEN_13639 = _GEN_16342 | _GEN_10543; // @[decode.scala 893:{68,68}]
  wire  _GEN_13640 = _GEN_16343 | _GEN_10544; // @[decode.scala 893:{68,68}]
  wire  _GEN_13641 = _GEN_16344 | _GEN_10545; // @[decode.scala 893:{68,68}]
  wire  _GEN_13642 = _GEN_16345 | _GEN_10546; // @[decode.scala 893:{68,68}]
  wire  _GEN_13643 = _GEN_16346 | _GEN_10547; // @[decode.scala 893:{68,68}]
  wire  _GEN_13644 = _GEN_16347 | _GEN_10548; // @[decode.scala 893:{68,68}]
  wire  _GEN_13645 = _GEN_16348 | _GEN_10549; // @[decode.scala 893:{68,68}]
  wire  _GEN_13646 = _GEN_16349 | _GEN_10550; // @[decode.scala 893:{68,68}]
  wire  _GEN_13647 = _GEN_16350 | _GEN_10551; // @[decode.scala 893:{68,68}]
  wire  _GEN_13648 = _GEN_16351 | _GEN_10552; // @[decode.scala 893:{68,68}]
  wire  _GEN_13649 = _GEN_16352 | _GEN_10553; // @[decode.scala 893:{68,68}]
  wire  _GEN_13650 = _GEN_16353 | _GEN_10554; // @[decode.scala 893:{68,68}]
  wire  _GEN_13651 = _GEN_16354 | _GEN_10555; // @[decode.scala 893:{68,68}]
  wire  _GEN_13652 = _GEN_16355 | _GEN_10556; // @[decode.scala 893:{68,68}]
  wire  _GEN_13653 = _GEN_16356 | _GEN_10557; // @[decode.scala 893:{68,68}]
  wire  _GEN_13655 = _GEN_16294 | _GEN_10655; // @[decode.scala 894:{68,68}]
  wire  _GEN_13656 = _GEN_16295 | _GEN_10656; // @[decode.scala 894:{68,68}]
  wire  _GEN_13657 = _GEN_16296 | _GEN_10657; // @[decode.scala 894:{68,68}]
  wire  _GEN_13658 = _GEN_16297 | _GEN_10658; // @[decode.scala 894:{68,68}]
  wire  _GEN_13659 = _GEN_16298 | _GEN_10659; // @[decode.scala 894:{68,68}]
  wire  _GEN_13660 = _GEN_16299 | _GEN_10660; // @[decode.scala 894:{68,68}]
  wire  _GEN_13661 = _GEN_16300 | _GEN_10661; // @[decode.scala 894:{68,68}]
  wire  _GEN_13662 = _GEN_16301 | _GEN_10662; // @[decode.scala 894:{68,68}]
  wire  _GEN_13663 = _GEN_16302 | _GEN_10663; // @[decode.scala 894:{68,68}]
  wire  _GEN_13664 = _GEN_16303 | _GEN_10664; // @[decode.scala 894:{68,68}]
  wire  _GEN_13665 = _GEN_16304 | _GEN_10665; // @[decode.scala 894:{68,68}]
  wire  _GEN_13666 = _GEN_16305 | _GEN_10666; // @[decode.scala 894:{68,68}]
  wire  _GEN_13667 = _GEN_16306 | _GEN_10667; // @[decode.scala 894:{68,68}]
  wire  _GEN_13668 = _GEN_16307 | _GEN_10668; // @[decode.scala 894:{68,68}]
  wire  _GEN_13669 = _GEN_16308 | _GEN_10669; // @[decode.scala 894:{68,68}]
  wire  _GEN_13670 = _GEN_16309 | _GEN_10670; // @[decode.scala 894:{68,68}]
  wire  _GEN_13671 = _GEN_16310 | _GEN_10671; // @[decode.scala 894:{68,68}]
  wire  _GEN_13672 = _GEN_16311 | _GEN_10672; // @[decode.scala 894:{68,68}]
  wire  _GEN_13673 = _GEN_16312 | _GEN_10673; // @[decode.scala 894:{68,68}]
  wire  _GEN_13674 = _GEN_16313 | _GEN_10674; // @[decode.scala 894:{68,68}]
  wire  _GEN_13675 = _GEN_16314 | _GEN_10675; // @[decode.scala 894:{68,68}]
  wire  _GEN_13676 = _GEN_16315 | _GEN_10676; // @[decode.scala 894:{68,68}]
  wire  _GEN_13677 = _GEN_16316 | _GEN_10677; // @[decode.scala 894:{68,68}]
  wire  _GEN_13678 = _GEN_16317 | _GEN_10678; // @[decode.scala 894:{68,68}]
  wire  _GEN_13679 = _GEN_16318 | _GEN_10679; // @[decode.scala 894:{68,68}]
  wire  _GEN_13680 = _GEN_16319 | _GEN_10680; // @[decode.scala 894:{68,68}]
  wire  _GEN_13681 = _GEN_16320 | _GEN_10681; // @[decode.scala 894:{68,68}]
  wire  _GEN_13682 = _GEN_16321 | _GEN_10682; // @[decode.scala 894:{68,68}]
  wire  _GEN_13683 = _GEN_16322 | _GEN_10683; // @[decode.scala 894:{68,68}]
  wire  _GEN_13684 = _GEN_16323 | _GEN_10684; // @[decode.scala 894:{68,68}]
  wire  _GEN_13685 = _GEN_16324 | _GEN_10685; // @[decode.scala 894:{68,68}]
  wire  _GEN_13686 = _GEN_16325 | _GEN_10686; // @[decode.scala 894:{68,68}]
  wire  _GEN_13687 = _GEN_16326 | _GEN_10687; // @[decode.scala 894:{68,68}]
  wire  _GEN_13688 = _GEN_16327 | _GEN_10688; // @[decode.scala 894:{68,68}]
  wire  _GEN_13689 = _GEN_16328 | _GEN_10689; // @[decode.scala 894:{68,68}]
  wire  _GEN_13690 = _GEN_16329 | _GEN_10690; // @[decode.scala 894:{68,68}]
  wire  _GEN_13691 = _GEN_16330 | _GEN_10691; // @[decode.scala 894:{68,68}]
  wire  _GEN_13692 = _GEN_16331 | _GEN_10692; // @[decode.scala 894:{68,68}]
  wire  _GEN_13693 = _GEN_16332 | _GEN_10693; // @[decode.scala 894:{68,68}]
  wire  _GEN_13694 = _GEN_16333 | _GEN_10694; // @[decode.scala 894:{68,68}]
  wire  _GEN_13695 = _GEN_16334 | _GEN_10695; // @[decode.scala 894:{68,68}]
  wire  _GEN_13696 = _GEN_16335 | _GEN_10696; // @[decode.scala 894:{68,68}]
  wire  _GEN_13697 = _GEN_16336 | _GEN_10697; // @[decode.scala 894:{68,68}]
  wire  _GEN_13698 = _GEN_16337 | _GEN_10698; // @[decode.scala 894:{68,68}]
  wire  _GEN_13699 = _GEN_16338 | _GEN_10699; // @[decode.scala 894:{68,68}]
  wire  _GEN_13700 = _GEN_16339 | _GEN_10700; // @[decode.scala 894:{68,68}]
  wire  _GEN_13701 = _GEN_16340 | _GEN_10701; // @[decode.scala 894:{68,68}]
  wire  _GEN_13702 = _GEN_16341 | _GEN_10702; // @[decode.scala 894:{68,68}]
  wire  _GEN_13703 = _GEN_16342 | _GEN_10703; // @[decode.scala 894:{68,68}]
  wire  _GEN_13704 = _GEN_16343 | _GEN_10704; // @[decode.scala 894:{68,68}]
  wire  _GEN_13705 = _GEN_16344 | _GEN_10705; // @[decode.scala 894:{68,68}]
  wire  _GEN_13706 = _GEN_16345 | _GEN_10706; // @[decode.scala 894:{68,68}]
  wire  _GEN_13707 = _GEN_16346 | _GEN_10707; // @[decode.scala 894:{68,68}]
  wire  _GEN_13708 = _GEN_16347 | _GEN_10708; // @[decode.scala 894:{68,68}]
  wire  _GEN_13709 = _GEN_16348 | _GEN_10709; // @[decode.scala 894:{68,68}]
  wire  _GEN_13710 = _GEN_16349 | _GEN_10710; // @[decode.scala 894:{68,68}]
  wire  _GEN_13711 = _GEN_16350 | _GEN_10711; // @[decode.scala 894:{68,68}]
  wire  _GEN_13712 = _GEN_16351 | _GEN_10712; // @[decode.scala 894:{68,68}]
  wire  _GEN_13713 = _GEN_16352 | _GEN_10713; // @[decode.scala 894:{68,68}]
  wire  _GEN_13714 = _GEN_16353 | _GEN_10714; // @[decode.scala 894:{68,68}]
  wire  _GEN_13715 = _GEN_16354 | _GEN_10715; // @[decode.scala 894:{68,68}]
  wire  _GEN_13716 = _GEN_16355 | _GEN_10716; // @[decode.scala 894:{68,68}]
  wire  _GEN_13717 = _GEN_16356 | _GEN_10717; // @[decode.scala 894:{68,68}]
  wire  _GEN_13719 = _GEN_16294 | _GEN_10815; // @[decode.scala 895:{68,68}]
  wire  _GEN_13720 = _GEN_16295 | _GEN_10816; // @[decode.scala 895:{68,68}]
  wire  _GEN_13721 = _GEN_16296 | _GEN_10817; // @[decode.scala 895:{68,68}]
  wire  _GEN_13722 = _GEN_16297 | _GEN_10818; // @[decode.scala 895:{68,68}]
  wire  _GEN_13723 = _GEN_16298 | _GEN_10819; // @[decode.scala 895:{68,68}]
  wire  _GEN_13724 = _GEN_16299 | _GEN_10820; // @[decode.scala 895:{68,68}]
  wire  _GEN_13725 = _GEN_16300 | _GEN_10821; // @[decode.scala 895:{68,68}]
  wire  _GEN_13726 = _GEN_16301 | _GEN_10822; // @[decode.scala 895:{68,68}]
  wire  _GEN_13727 = _GEN_16302 | _GEN_10823; // @[decode.scala 895:{68,68}]
  wire  _GEN_13728 = _GEN_16303 | _GEN_10824; // @[decode.scala 895:{68,68}]
  wire  _GEN_13729 = _GEN_16304 | _GEN_10825; // @[decode.scala 895:{68,68}]
  wire  _GEN_13730 = _GEN_16305 | _GEN_10826; // @[decode.scala 895:{68,68}]
  wire  _GEN_13731 = _GEN_16306 | _GEN_10827; // @[decode.scala 895:{68,68}]
  wire  _GEN_13732 = _GEN_16307 | _GEN_10828; // @[decode.scala 895:{68,68}]
  wire  _GEN_13733 = _GEN_16308 | _GEN_10829; // @[decode.scala 895:{68,68}]
  wire  _GEN_13734 = _GEN_16309 | _GEN_10830; // @[decode.scala 895:{68,68}]
  wire  _GEN_13735 = _GEN_16310 | _GEN_10831; // @[decode.scala 895:{68,68}]
  wire  _GEN_13736 = _GEN_16311 | _GEN_10832; // @[decode.scala 895:{68,68}]
  wire  _GEN_13737 = _GEN_16312 | _GEN_10833; // @[decode.scala 895:{68,68}]
  wire  _GEN_13738 = _GEN_16313 | _GEN_10834; // @[decode.scala 895:{68,68}]
  wire  _GEN_13739 = _GEN_16314 | _GEN_10835; // @[decode.scala 895:{68,68}]
  wire  _GEN_13740 = _GEN_16315 | _GEN_10836; // @[decode.scala 895:{68,68}]
  wire  _GEN_13741 = _GEN_16316 | _GEN_10837; // @[decode.scala 895:{68,68}]
  wire  _GEN_13742 = _GEN_16317 | _GEN_10838; // @[decode.scala 895:{68,68}]
  wire  _GEN_13743 = _GEN_16318 | _GEN_10839; // @[decode.scala 895:{68,68}]
  wire  _GEN_13744 = _GEN_16319 | _GEN_10840; // @[decode.scala 895:{68,68}]
  wire  _GEN_13745 = _GEN_16320 | _GEN_10841; // @[decode.scala 895:{68,68}]
  wire  _GEN_13746 = _GEN_16321 | _GEN_10842; // @[decode.scala 895:{68,68}]
  wire  _GEN_13747 = _GEN_16322 | _GEN_10843; // @[decode.scala 895:{68,68}]
  wire  _GEN_13748 = _GEN_16323 | _GEN_10844; // @[decode.scala 895:{68,68}]
  wire  _GEN_13749 = _GEN_16324 | _GEN_10845; // @[decode.scala 895:{68,68}]
  wire  _GEN_13750 = _GEN_16325 | _GEN_10846; // @[decode.scala 895:{68,68}]
  wire  _GEN_13751 = _GEN_16326 | _GEN_10847; // @[decode.scala 895:{68,68}]
  wire  _GEN_13752 = _GEN_16327 | _GEN_10848; // @[decode.scala 895:{68,68}]
  wire  _GEN_13753 = _GEN_16328 | _GEN_10849; // @[decode.scala 895:{68,68}]
  wire  _GEN_13754 = _GEN_16329 | _GEN_10850; // @[decode.scala 895:{68,68}]
  wire  _GEN_13755 = _GEN_16330 | _GEN_10851; // @[decode.scala 895:{68,68}]
  wire  _GEN_13756 = _GEN_16331 | _GEN_10852; // @[decode.scala 895:{68,68}]
  wire  _GEN_13757 = _GEN_16332 | _GEN_10853; // @[decode.scala 895:{68,68}]
  wire  _GEN_13758 = _GEN_16333 | _GEN_10854; // @[decode.scala 895:{68,68}]
  wire  _GEN_13759 = _GEN_16334 | _GEN_10855; // @[decode.scala 895:{68,68}]
  wire  _GEN_13760 = _GEN_16335 | _GEN_10856; // @[decode.scala 895:{68,68}]
  wire  _GEN_13761 = _GEN_16336 | _GEN_10857; // @[decode.scala 895:{68,68}]
  wire  _GEN_13762 = _GEN_16337 | _GEN_10858; // @[decode.scala 895:{68,68}]
  wire  _GEN_13763 = _GEN_16338 | _GEN_10859; // @[decode.scala 895:{68,68}]
  wire  _GEN_13764 = _GEN_16339 | _GEN_10860; // @[decode.scala 895:{68,68}]
  wire  _GEN_13765 = _GEN_16340 | _GEN_10861; // @[decode.scala 895:{68,68}]
  wire  _GEN_13766 = _GEN_16341 | _GEN_10862; // @[decode.scala 895:{68,68}]
  wire  _GEN_13767 = _GEN_16342 | _GEN_10863; // @[decode.scala 895:{68,68}]
  wire  _GEN_13768 = _GEN_16343 | _GEN_10864; // @[decode.scala 895:{68,68}]
  wire  _GEN_13769 = _GEN_16344 | _GEN_10865; // @[decode.scala 895:{68,68}]
  wire  _GEN_13770 = _GEN_16345 | _GEN_10866; // @[decode.scala 895:{68,68}]
  wire  _GEN_13771 = _GEN_16346 | _GEN_10867; // @[decode.scala 895:{68,68}]
  wire  _GEN_13772 = _GEN_16347 | _GEN_10868; // @[decode.scala 895:{68,68}]
  wire  _GEN_13773 = _GEN_16348 | _GEN_10869; // @[decode.scala 895:{68,68}]
  wire  _GEN_13774 = _GEN_16349 | _GEN_10870; // @[decode.scala 895:{68,68}]
  wire  _GEN_13775 = _GEN_16350 | _GEN_10871; // @[decode.scala 895:{68,68}]
  wire  _GEN_13776 = _GEN_16351 | _GEN_10872; // @[decode.scala 895:{68,68}]
  wire  _GEN_13777 = _GEN_16352 | _GEN_10873; // @[decode.scala 895:{68,68}]
  wire  _GEN_13778 = _GEN_16353 | _GEN_10874; // @[decode.scala 895:{68,68}]
  wire  _GEN_13779 = _GEN_16354 | _GEN_10875; // @[decode.scala 895:{68,68}]
  wire  _GEN_13780 = _GEN_16355 | _GEN_10876; // @[decode.scala 895:{68,68}]
  wire  _GEN_13781 = _GEN_16356 | _GEN_10877; // @[decode.scala 895:{68,68}]
  wire  _GEN_13847 = _T_474 ? _GEN_13495 : _GEN_6180; // @[decode.scala 889:5]
  wire  _GEN_13848 = _T_474 ? _GEN_13496 : _GEN_6181; // @[decode.scala 889:5]
  wire  _GEN_13849 = _T_474 ? _GEN_13497 : _GEN_6182; // @[decode.scala 889:5]
  wire  _GEN_13850 = _T_474 ? _GEN_13498 : _GEN_6183; // @[decode.scala 889:5]
  wire  _GEN_13851 = _T_474 ? _GEN_13499 : _GEN_6184; // @[decode.scala 889:5]
  wire  _GEN_13852 = _T_474 ? _GEN_13500 : _GEN_6185; // @[decode.scala 889:5]
  wire  _GEN_13853 = _T_474 ? _GEN_13501 : _GEN_6186; // @[decode.scala 889:5]
  wire  _GEN_13854 = _T_474 ? _GEN_13502 : _GEN_6187; // @[decode.scala 889:5]
  wire  _GEN_13855 = _T_474 ? _GEN_13503 : _GEN_6188; // @[decode.scala 889:5]
  wire  _GEN_13856 = _T_474 ? _GEN_13504 : _GEN_6189; // @[decode.scala 889:5]
  wire  _GEN_13857 = _T_474 ? _GEN_13505 : _GEN_6190; // @[decode.scala 889:5]
  wire  _GEN_13858 = _T_474 ? _GEN_13506 : _GEN_6191; // @[decode.scala 889:5]
  wire  _GEN_13859 = _T_474 ? _GEN_13507 : _GEN_6192; // @[decode.scala 889:5]
  wire  _GEN_13860 = _T_474 ? _GEN_13508 : _GEN_6193; // @[decode.scala 889:5]
  wire  _GEN_13861 = _T_474 ? _GEN_13509 : _GEN_6194; // @[decode.scala 889:5]
  wire  _GEN_13862 = _T_474 ? _GEN_13510 : _GEN_6195; // @[decode.scala 889:5]
  wire  _GEN_13863 = _T_474 ? _GEN_13511 : _GEN_6196; // @[decode.scala 889:5]
  wire  _GEN_13864 = _T_474 ? _GEN_13512 : _GEN_6197; // @[decode.scala 889:5]
  wire  _GEN_13865 = _T_474 ? _GEN_13513 : _GEN_6198; // @[decode.scala 889:5]
  wire  _GEN_13866 = _T_474 ? _GEN_13514 : _GEN_6199; // @[decode.scala 889:5]
  wire  _GEN_13867 = _T_474 ? _GEN_13515 : _GEN_6200; // @[decode.scala 889:5]
  wire  _GEN_13868 = _T_474 ? _GEN_13516 : _GEN_6201; // @[decode.scala 889:5]
  wire  _GEN_13869 = _T_474 ? _GEN_13517 : _GEN_6202; // @[decode.scala 889:5]
  wire  _GEN_13870 = _T_474 ? _GEN_13518 : _GEN_6203; // @[decode.scala 889:5]
  wire  _GEN_13871 = _T_474 ? _GEN_13519 : _GEN_6204; // @[decode.scala 889:5]
  wire  _GEN_13872 = _T_474 ? _GEN_13520 : _GEN_6205; // @[decode.scala 889:5]
  wire  _GEN_13873 = _T_474 ? _GEN_13521 : _GEN_6206; // @[decode.scala 889:5]
  wire  _GEN_13874 = _T_474 ? _GEN_13522 : _GEN_6207; // @[decode.scala 889:5]
  wire  _GEN_13875 = _T_474 ? _GEN_13523 : _GEN_6208; // @[decode.scala 889:5]
  wire  _GEN_13876 = _T_474 ? _GEN_13524 : _GEN_6209; // @[decode.scala 889:5]
  wire  _GEN_13877 = _T_474 ? _GEN_13525 : _GEN_6210; // @[decode.scala 889:5]
  wire  _GEN_14135 = currentPrivilege == 64'h2200001800 ? mie[7] : mstatus[3] & mie[7]; // @[decode.scala 903:44 905:22 908:22]
  wire [63:0] _GEN_16609 = reset ? 64'h0 : _GEN_10951; // @[decode.scala 242:{27,27}]
  wire [126:0] _GEN_16610 = reset ? 127'h0 : _GEN_12932; // @[decode.scala 504:{28,28}]
  assign fromFetch_ready = ~stateRegInputBuf ? _GEN_13363 : stateRegInputBuf & _GEN_13374; // @[decode.scala 792:28]
  assign fromFetch_expected_valid = expectedPC != 64'h0; // @[decode.scala 261:42]
  assign fromFetch_expected_pc = expectedPC; // @[decode.scala 262:28]
  assign fromFetch_expected_coherency = coherency; // @[decode.scala 263:32]
  assign toExec_ready = ~stateRegOutputBuf ? 1'h0 : stateRegOutputBuf & _GEN_13361; // @[decode.scala 846:29]
  assign toExec_instruction = outputBuffer_instruction; // @[decode.scala 250:22]
  assign toExec_pc = outputBuffer_pc; // @[decode.scala 251:22]
  assign toExec_PRFDest = outputBuffer_PRFDest; // @[decode.scala 252:22]
  assign toExec_rs1Addr = outputBuffer_rs1Addr; // @[decode.scala 253:22]
  assign toExec_rs1Ready = 6'h3f == outputBuffer_rs1Addr ? PRFValidList_63 : _GEN_74; // @[decode.scala 254:{22,22}]
  assign toExec_rs2Addr = outputBuffer_rs2Addr; // @[decode.scala 255:22]
  assign toExec_rs2Ready = _GEN_181 | (3'h1 == toExec_rs2Ready_insType | 3'h4 == toExec_rs2Ready_insType | 3'h5 ==
    toExec_rs2Ready_insType); // @[decode.scala 256:60]
  assign toExec_branchMask = {toExec_branchMask_hi,toExec_branchMask_lo}; // @[decode.scala 258:49]
  assign jumpAddrWrite_ready = validOutputBuf & (unconditionalJumps | csrIns); // @[decode.scala 265:44]
  assign jumpAddrWrite_PRFDest = outputBuffer_PRFDest; // @[decode.scala 266:26]
  assign jumpAddrWrite_linkAddr = unconditionalJumps ? _GEN_185 : csrReadDataReg; // @[decode.scala 267:28 268:28 274:28]
  assign branchPCs_branchPCReady = branchBuffer_branchPCReady; // @[decode.scala 279:30]
  assign branchPCs_branchPC = branchBuffer_branchPC; // @[decode.scala 281:30]
  assign branchPCs_predictedPCReady = branchBuffer_predictedPCReady; // @[decode.scala 280:30]
  assign branchPCs_predictedPC = branchBuffer_predictedPC; // @[decode.scala 282:30]
  assign branchPCs_branchMask = branchPCMask; // @[decode.scala 283:30]
  assign canTakeInterrupt = stallReg ? 1'h0 : _GEN_14135; // @[decode.scala 899:18 902:22]
  always @(posedge clock) begin
    if (reset) begin // @[decode.scala 111:28]
      inputBuffer_pc <= 64'hffffffc; // @[decode.scala 111:28]
    end else if (fromFetch_fired & readyInputBuf) begin // @[decode.scala 202:42]
      inputBuffer_pc <= fromFetch_pc; // @[decode.scala 204:29]
    end
    if (reset) begin // @[decode.scala 111:28]
      inputBuffer_instruction <= 32'h0; // @[decode.scala 111:28]
    end else if (fromFetch_fired & readyInputBuf) begin // @[decode.scala 202:42]
      inputBuffer_instruction <= fromFetch_instruction; // @[decode.scala 203:29]
    end
    if (reset) begin // @[decode.scala 120:29]
      outputBuffer_instruction <= 32'h0; // @[decode.scala 120:29]
    end else if (validInputBuf & readyOutputBuf) begin // @[decode.scala 212:41]
      outputBuffer_instruction <= inputBuffer_instruction; // @[decode.scala 213:30]
    end
    if (reset) begin // @[decode.scala 120:29]
      outputBuffer_pc <= 64'h0; // @[decode.scala 120:29]
    end else if (validInputBuf & readyOutputBuf) begin // @[decode.scala 212:41]
      outputBuffer_pc <= inputBuffer_pc; // @[decode.scala 214:30]
    end
    if (reset) begin // @[decode.scala 120:29]
      outputBuffer_PRFDest <= 6'h0; // @[decode.scala 120:29]
    end else if (validInputBuf & readyOutputBuf) begin // @[decode.scala 212:41]
      if (PRFFreeList_0) begin // @[Mux.scala 47:70]
        outputBuffer_PRFDest <= 6'h0;
      end else if (PRFFreeList_1) begin // @[Mux.scala 47:70]
        outputBuffer_PRFDest <= 6'h1;
      end else begin
        outputBuffer_PRFDest <= _freeRegAddr_T_60;
      end
    end
    if (reset) begin // @[decode.scala 120:29]
      outputBuffer_rs1Addr <= 6'h0; // @[decode.scala 120:29]
    end else if (validInputBuf & readyOutputBuf) begin // @[decode.scala 212:41]
      if (5'h1f == rs1) begin // @[decode.scala 332:12]
        outputBuffer_rs1Addr <= frontEndRegMap_31; // @[decode.scala 332:12]
      end else if (5'h1e == rs1) begin // @[decode.scala 332:12]
        outputBuffer_rs1Addr <= frontEndRegMap_30; // @[decode.scala 332:12]
      end else begin
        outputBuffer_rs1Addr <= _GEN_237;
      end
    end
    if (reset) begin // @[decode.scala 120:29]
      outputBuffer_rs2Addr <= 6'h0; // @[decode.scala 120:29]
    end else if (validInputBuf & readyOutputBuf) begin // @[decode.scala 212:41]
      if (5'h1f == rs2) begin // @[decode.scala 333:12]
        outputBuffer_rs2Addr <= frontEndRegMap_31; // @[decode.scala 333:12]
      end else if (5'h1e == rs2) begin // @[decode.scala 333:12]
        outputBuffer_rs2Addr <= frontEndRegMap_30; // @[decode.scala 333:12]
      end else begin
        outputBuffer_rs2Addr <= _GEN_269;
      end
    end
    if (reset) begin // @[decode.scala 120:29]
      outputBuffer_immediate <= 64'h0; // @[decode.scala 120:29]
    end else if (validInputBuf & readyOutputBuf) begin // @[decode.scala 212:41]
      outputBuffer_immediate <= immediate_immediate; // @[decode.scala 218:30]
    end
    if (reset) begin // @[decode.scala 142:29]
      branchBuffer_branchPCReady <= 1'h0; // @[decode.scala 142:29]
    end else begin
      branchBuffer_branchPCReady <= _T_445 & validInputBuf & readyOutputBuf; // @[decode.scala 484:30]
    end
    if (reset) begin // @[decode.scala 142:29]
      branchBuffer_predictedPCReady <= 1'h0; // @[decode.scala 142:29]
    end else begin
      branchBuffer_predictedPCReady <= branchReg & validInputBuf & readyOutputBuf; // @[decode.scala 485:33]
    end
    if (reset) begin // @[decode.scala 142:29]
      branchBuffer_branchPC <= 64'h0; // @[decode.scala 142:29]
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        branchBuffer_branchPC <= inputBuffer_pc; // @[decode.scala 422:29]
      end
    end
    if (reset) begin // @[decode.scala 142:29]
      branchBuffer_predictedPC <= 64'h0; // @[decode.scala 142:29]
    end else if (_toExec_branchMask_T != 5'h0 & validInputBuf & readyOutputBuf) begin // @[decode.scala 480:83]
      branchBuffer_predictedPC <= inputBuffer_pc; // @[decode.scala 481:30]
    end
    if (reset) begin // @[decode.scala 142:29]
      branchBuffer_branchMask_0 <= 1'h0; // @[decode.scala 142:29]
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        branchBuffer_branchMask_0 <= _GEN_6757;
      end else begin
        branchBuffer_branchMask_0 <= _GEN_6109;
      end
    end else begin
      branchBuffer_branchMask_0 <= _GEN_6109;
    end
    if (reset) begin // @[decode.scala 142:29]
      branchBuffer_branchMask_1 <= 1'h0; // @[decode.scala 142:29]
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        branchBuffer_branchMask_1 <= _GEN_6758;
      end else begin
        branchBuffer_branchMask_1 <= _GEN_6110;
      end
    end else begin
      branchBuffer_branchMask_1 <= _GEN_6110;
    end
    if (reset) begin // @[decode.scala 142:29]
      branchBuffer_branchMask_2 <= 1'h0; // @[decode.scala 142:29]
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        branchBuffer_branchMask_2 <= _GEN_6759;
      end else begin
        branchBuffer_branchMask_2 <= _GEN_6111;
      end
    end else begin
      branchBuffer_branchMask_2 <= _GEN_6111;
    end
    if (reset) begin // @[decode.scala 142:29]
      branchBuffer_branchMask_3 <= 1'h0; // @[decode.scala 142:29]
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        branchBuffer_branchMask_3 <= _GEN_6760;
      end else begin
        branchBuffer_branchMask_3 <= _GEN_6112;
      end
    end else begin
      branchBuffer_branchMask_3 <= _GEN_6112;
    end
    branchBuffer_branchMask_4 <= reset | _GEN_10301; // @[decode.scala 142:{29,29}]
    if (reset) begin // @[decode.scala 178:30]
      branchTracker <= 3'h0; // @[decode.scala 178:30]
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        branchTracker <= _branchTracker_T_3; // @[decode.scala 473:21]
      end else begin
        branchTracker <= _GEN_6108;
      end
    end else begin
      branchTracker <= _GEN_6108;
    end
    if (reset) begin // @[decode.scala 188:27]
      expectedPC <= 64'h10000000; // @[decode.scala 188:27]
    end else if (_T_256 & writeBackResult_instruction[14:12] == 3'h0) begin // @[decode.scala 744:126]
      if (writeBackResult_instruction[31:20] == 12'h302) begin // @[decode.scala 745:60]
        expectedPC <= mepc; // @[decode.scala 748:18]
      end else if (~(|writeBackResult_instruction[31:20])) begin // @[decode.scala 750:58]
        expectedPC <= mtvec; // @[decode.scala 756:18]
      end else begin
        expectedPC <= _GEN_12955;
      end
    end else if (_fromFetch_expected_valid_T & fromFetch_fired & fromFetch_expected_pc == fromFetch_pc) begin // @[decode.scala 487:89]
      expectedPC <= 64'h0; // @[decode.scala 488:16]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      expectedPC <= _GEN_5465;
    end
    if (reset) begin // @[decode.scala 189:26]
      coherency <= 1'h0; // @[decode.scala 189:26]
    end else if (_fromFetch_expected_valid_T & fromFetch_fired & fromFetch_expected_pc == fromFetch_pc) begin // @[decode.scala 487:89]
      coherency <= 1'h0; // @[decode.scala 489:15]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        coherency <= _GEN_5458;
      end
    end
    if (reset) begin // @[decode.scala 193:34]
      stateRegInputBuf <= 1'h0; // @[decode.scala 193:34]
    end else if (~stateRegInputBuf) begin // @[decode.scala 792:28]
      if (branchEvalIn_fired & ~branchEvalIn_passFail) begin // @[decode.scala 794:58]
        stateRegInputBuf <= 1'h0; // @[decode.scala 795:26]
      end else if (fromFetch_fired) begin // @[decode.scala 802:31]
        stateRegInputBuf <= _GEN_13357;
      end
    end else if (stateRegInputBuf) begin // @[decode.scala 792:28]
      if (_T_435) begin // @[decode.scala 817:58]
        stateRegInputBuf <= 1'h0; // @[decode.scala 818:26]
      end else begin
        stateRegInputBuf <= _GEN_13369;
      end
    end
    if (reset) begin // @[decode.scala 194:34]
      stateRegOutputBuf <= 1'h0; // @[decode.scala 194:34]
    end else if (~stateRegOutputBuf) begin // @[decode.scala 846:29]
      if (_T_435) begin // @[decode.scala 848:58]
        stateRegOutputBuf <= 1'h0; // @[decode.scala 849:27]
      end else begin
        stateRegOutputBuf <= _GEN_13383;
      end
    end else if (stateRegOutputBuf) begin // @[decode.scala 846:29]
      if (_T_435) begin // @[decode.scala 861:58]
        stateRegOutputBuf <= 1'h0; // @[decode.scala 862:27]
      end else begin
        stateRegOutputBuf <= _GEN_13389;
      end
    end
    if (reset) begin // @[decode.scala 196:25]
      stallReg <= 1'h0; // @[decode.scala 196:25]
    end else if (~stateRegInputBuf) begin // @[decode.scala 792:28]
      stallReg <= _GEN_13362;
    end else if (stateRegInputBuf) begin // @[decode.scala 792:28]
      stallReg <= _GEN_13362;
    end else begin
      stallReg <= _GEN_10979;
    end
    if (fromFetch_fired & readyInputBuf) begin // @[decode.scala 202:42]
      if (fromFetch_instruction[6:0] == 7'h73) begin // @[decode.scala 205:97]
        ecallPC <= fromFetch_pc; // @[decode.scala 207:15]
      end
    end
    PRFValidList_0 <= reset | _GEN_13292; // @[decode.scala 199:{29,29}]
    PRFValidList_1 <= reset | _GEN_13293; // @[decode.scala 199:{29,29}]
    PRFValidList_2 <= reset | _GEN_13294; // @[decode.scala 199:{29,29}]
    PRFValidList_3 <= reset | _GEN_13295; // @[decode.scala 199:{29,29}]
    PRFValidList_4 <= reset | _GEN_13296; // @[decode.scala 199:{29,29}]
    PRFValidList_5 <= reset | _GEN_13297; // @[decode.scala 199:{29,29}]
    PRFValidList_6 <= reset | _GEN_13298; // @[decode.scala 199:{29,29}]
    PRFValidList_7 <= reset | _GEN_13299; // @[decode.scala 199:{29,29}]
    PRFValidList_8 <= reset | _GEN_13300; // @[decode.scala 199:{29,29}]
    PRFValidList_9 <= reset | _GEN_13301; // @[decode.scala 199:{29,29}]
    PRFValidList_10 <= reset | _GEN_13302; // @[decode.scala 199:{29,29}]
    PRFValidList_11 <= reset | _GEN_13303; // @[decode.scala 199:{29,29}]
    PRFValidList_12 <= reset | _GEN_13304; // @[decode.scala 199:{29,29}]
    PRFValidList_13 <= reset | _GEN_13305; // @[decode.scala 199:{29,29}]
    PRFValidList_14 <= reset | _GEN_13306; // @[decode.scala 199:{29,29}]
    PRFValidList_15 <= reset | _GEN_13307; // @[decode.scala 199:{29,29}]
    PRFValidList_16 <= reset | _GEN_13308; // @[decode.scala 199:{29,29}]
    PRFValidList_17 <= reset | _GEN_13309; // @[decode.scala 199:{29,29}]
    PRFValidList_18 <= reset | _GEN_13310; // @[decode.scala 199:{29,29}]
    PRFValidList_19 <= reset | _GEN_13311; // @[decode.scala 199:{29,29}]
    PRFValidList_20 <= reset | _GEN_13312; // @[decode.scala 199:{29,29}]
    PRFValidList_21 <= reset | _GEN_13313; // @[decode.scala 199:{29,29}]
    PRFValidList_22 <= reset | _GEN_13314; // @[decode.scala 199:{29,29}]
    PRFValidList_23 <= reset | _GEN_13315; // @[decode.scala 199:{29,29}]
    PRFValidList_24 <= reset | _GEN_13316; // @[decode.scala 199:{29,29}]
    PRFValidList_25 <= reset | _GEN_13317; // @[decode.scala 199:{29,29}]
    PRFValidList_26 <= reset | _GEN_13318; // @[decode.scala 199:{29,29}]
    PRFValidList_27 <= reset | _GEN_13319; // @[decode.scala 199:{29,29}]
    PRFValidList_28 <= reset | _GEN_13320; // @[decode.scala 199:{29,29}]
    PRFValidList_29 <= reset | _GEN_13321; // @[decode.scala 199:{29,29}]
    PRFValidList_30 <= reset | _GEN_13322; // @[decode.scala 199:{29,29}]
    PRFValidList_31 <= reset | _GEN_13323; // @[decode.scala 199:{29,29}]
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_32 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_32 <= 6'h20 == writeAddrPRF_exec3Addr | _GEN_13196;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_32 <= 6'h20 == writeAddrPRF_exec2Addr | _GEN_13068;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_32 <= 6'h20 == writeAddrPRF_exec1Addr | _GEN_6244;
    end else begin
      PRFValidList_32 <= _GEN_6244;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_33 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_33 <= 6'h21 == writeAddrPRF_exec3Addr | _GEN_13197;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_33 <= 6'h21 == writeAddrPRF_exec2Addr | _GEN_13069;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_33 <= 6'h21 == writeAddrPRF_exec1Addr | _GEN_6245;
    end else begin
      PRFValidList_33 <= _GEN_6245;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_34 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_34 <= 6'h22 == writeAddrPRF_exec3Addr | _GEN_13198;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_34 <= 6'h22 == writeAddrPRF_exec2Addr | _GEN_13070;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_34 <= 6'h22 == writeAddrPRF_exec1Addr | _GEN_6246;
    end else begin
      PRFValidList_34 <= _GEN_6246;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_35 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_35 <= 6'h23 == writeAddrPRF_exec3Addr | _GEN_13199;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_35 <= 6'h23 == writeAddrPRF_exec2Addr | _GEN_13071;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_35 <= 6'h23 == writeAddrPRF_exec1Addr | _GEN_6247;
    end else begin
      PRFValidList_35 <= _GEN_6247;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_36 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_36 <= 6'h24 == writeAddrPRF_exec3Addr | _GEN_13200;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_36 <= 6'h24 == writeAddrPRF_exec2Addr | _GEN_13072;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_36 <= 6'h24 == writeAddrPRF_exec1Addr | _GEN_6248;
    end else begin
      PRFValidList_36 <= _GEN_6248;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_37 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_37 <= 6'h25 == writeAddrPRF_exec3Addr | _GEN_13201;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_37 <= 6'h25 == writeAddrPRF_exec2Addr | _GEN_13073;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_37 <= 6'h25 == writeAddrPRF_exec1Addr | _GEN_6249;
    end else begin
      PRFValidList_37 <= _GEN_6249;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_38 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_38 <= 6'h26 == writeAddrPRF_exec3Addr | _GEN_13202;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_38 <= 6'h26 == writeAddrPRF_exec2Addr | _GEN_13074;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_38 <= 6'h26 == writeAddrPRF_exec1Addr | _GEN_6250;
    end else begin
      PRFValidList_38 <= _GEN_6250;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_39 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_39 <= 6'h27 == writeAddrPRF_exec3Addr | _GEN_13203;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_39 <= 6'h27 == writeAddrPRF_exec2Addr | _GEN_13075;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_39 <= 6'h27 == writeAddrPRF_exec1Addr | _GEN_6251;
    end else begin
      PRFValidList_39 <= _GEN_6251;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_40 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_40 <= 6'h28 == writeAddrPRF_exec3Addr | _GEN_13204;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_40 <= 6'h28 == writeAddrPRF_exec2Addr | _GEN_13076;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_40 <= 6'h28 == writeAddrPRF_exec1Addr | _GEN_6252;
    end else begin
      PRFValidList_40 <= _GEN_6252;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_41 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_41 <= 6'h29 == writeAddrPRF_exec3Addr | _GEN_13205;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_41 <= 6'h29 == writeAddrPRF_exec2Addr | _GEN_13077;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_41 <= 6'h29 == writeAddrPRF_exec1Addr | _GEN_6253;
    end else begin
      PRFValidList_41 <= _GEN_6253;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_42 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_42 <= 6'h2a == writeAddrPRF_exec3Addr | _GEN_13206;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_42 <= 6'h2a == writeAddrPRF_exec2Addr | _GEN_13078;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_42 <= 6'h2a == writeAddrPRF_exec1Addr | _GEN_6254;
    end else begin
      PRFValidList_42 <= _GEN_6254;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_43 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_43 <= 6'h2b == writeAddrPRF_exec3Addr | _GEN_13207;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_43 <= 6'h2b == writeAddrPRF_exec2Addr | _GEN_13079;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_43 <= 6'h2b == writeAddrPRF_exec1Addr | _GEN_6255;
    end else begin
      PRFValidList_43 <= _GEN_6255;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_44 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_44 <= 6'h2c == writeAddrPRF_exec3Addr | _GEN_13208;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_44 <= 6'h2c == writeAddrPRF_exec2Addr | _GEN_13080;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_44 <= 6'h2c == writeAddrPRF_exec1Addr | _GEN_6256;
    end else begin
      PRFValidList_44 <= _GEN_6256;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_45 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_45 <= 6'h2d == writeAddrPRF_exec3Addr | _GEN_13209;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_45 <= 6'h2d == writeAddrPRF_exec2Addr | _GEN_13081;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_45 <= 6'h2d == writeAddrPRF_exec1Addr | _GEN_6257;
    end else begin
      PRFValidList_45 <= _GEN_6257;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_46 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_46 <= 6'h2e == writeAddrPRF_exec3Addr | _GEN_13210;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_46 <= 6'h2e == writeAddrPRF_exec2Addr | _GEN_13082;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_46 <= 6'h2e == writeAddrPRF_exec1Addr | _GEN_6258;
    end else begin
      PRFValidList_46 <= _GEN_6258;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_47 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_47 <= 6'h2f == writeAddrPRF_exec3Addr | _GEN_13211;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_47 <= 6'h2f == writeAddrPRF_exec2Addr | _GEN_13083;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_47 <= 6'h2f == writeAddrPRF_exec1Addr | _GEN_6259;
    end else begin
      PRFValidList_47 <= _GEN_6259;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_48 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_48 <= 6'h30 == writeAddrPRF_exec3Addr | _GEN_13212;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_48 <= 6'h30 == writeAddrPRF_exec2Addr | _GEN_13084;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_48 <= 6'h30 == writeAddrPRF_exec1Addr | _GEN_6260;
    end else begin
      PRFValidList_48 <= _GEN_6260;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_49 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_49 <= 6'h31 == writeAddrPRF_exec3Addr | _GEN_13213;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_49 <= 6'h31 == writeAddrPRF_exec2Addr | _GEN_13085;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_49 <= 6'h31 == writeAddrPRF_exec1Addr | _GEN_6261;
    end else begin
      PRFValidList_49 <= _GEN_6261;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_50 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_50 <= 6'h32 == writeAddrPRF_exec3Addr | _GEN_13214;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_50 <= 6'h32 == writeAddrPRF_exec2Addr | _GEN_13086;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_50 <= 6'h32 == writeAddrPRF_exec1Addr | _GEN_6262;
    end else begin
      PRFValidList_50 <= _GEN_6262;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_51 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_51 <= 6'h33 == writeAddrPRF_exec3Addr | _GEN_13215;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_51 <= 6'h33 == writeAddrPRF_exec2Addr | _GEN_13087;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_51 <= 6'h33 == writeAddrPRF_exec1Addr | _GEN_6263;
    end else begin
      PRFValidList_51 <= _GEN_6263;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_52 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_52 <= 6'h34 == writeAddrPRF_exec3Addr | _GEN_13216;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_52 <= 6'h34 == writeAddrPRF_exec2Addr | _GEN_13088;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_52 <= 6'h34 == writeAddrPRF_exec1Addr | _GEN_6264;
    end else begin
      PRFValidList_52 <= _GEN_6264;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_53 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_53 <= 6'h35 == writeAddrPRF_exec3Addr | _GEN_13217;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_53 <= 6'h35 == writeAddrPRF_exec2Addr | _GEN_13089;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_53 <= 6'h35 == writeAddrPRF_exec1Addr | _GEN_6265;
    end else begin
      PRFValidList_53 <= _GEN_6265;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_54 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_54 <= 6'h36 == writeAddrPRF_exec3Addr | _GEN_13218;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_54 <= 6'h36 == writeAddrPRF_exec2Addr | _GEN_13090;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_54 <= 6'h36 == writeAddrPRF_exec1Addr | _GEN_6266;
    end else begin
      PRFValidList_54 <= _GEN_6266;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_55 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_55 <= 6'h37 == writeAddrPRF_exec3Addr | _GEN_13219;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_55 <= 6'h37 == writeAddrPRF_exec2Addr | _GEN_13091;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_55 <= 6'h37 == writeAddrPRF_exec1Addr | _GEN_6267;
    end else begin
      PRFValidList_55 <= _GEN_6267;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_56 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_56 <= 6'h38 == writeAddrPRF_exec3Addr | _GEN_13220;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_56 <= 6'h38 == writeAddrPRF_exec2Addr | _GEN_13092;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_56 <= 6'h38 == writeAddrPRF_exec1Addr | _GEN_6268;
    end else begin
      PRFValidList_56 <= _GEN_6268;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_57 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_57 <= 6'h39 == writeAddrPRF_exec3Addr | _GEN_13221;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_57 <= 6'h39 == writeAddrPRF_exec2Addr | _GEN_13093;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_57 <= 6'h39 == writeAddrPRF_exec1Addr | _GEN_6269;
    end else begin
      PRFValidList_57 <= _GEN_6269;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_58 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_58 <= 6'h3a == writeAddrPRF_exec3Addr | _GEN_13222;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_58 <= 6'h3a == writeAddrPRF_exec2Addr | _GEN_13094;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_58 <= 6'h3a == writeAddrPRF_exec1Addr | _GEN_6270;
    end else begin
      PRFValidList_58 <= _GEN_6270;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_59 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_59 <= 6'h3b == writeAddrPRF_exec3Addr | _GEN_13223;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_59 <= 6'h3b == writeAddrPRF_exec2Addr | _GEN_13095;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_59 <= 6'h3b == writeAddrPRF_exec1Addr | _GEN_6271;
    end else begin
      PRFValidList_59 <= _GEN_6271;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_60 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_60 <= 6'h3c == writeAddrPRF_exec3Addr | _GEN_13224;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_60 <= 6'h3c == writeAddrPRF_exec2Addr | _GEN_13096;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_60 <= 6'h3c == writeAddrPRF_exec1Addr | _GEN_6272;
    end else begin
      PRFValidList_60 <= _GEN_6272;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_61 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_61 <= 6'h3d == writeAddrPRF_exec3Addr | _GEN_13225;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_61 <= 6'h3d == writeAddrPRF_exec2Addr | _GEN_13097;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_61 <= 6'h3d == writeAddrPRF_exec1Addr | _GEN_6273;
    end else begin
      PRFValidList_61 <= _GEN_6273;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_62 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_62 <= 6'h3e == writeAddrPRF_exec3Addr | _GEN_13226;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_62 <= 6'h3e == writeAddrPRF_exec2Addr | _GEN_13098;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_62 <= 6'h3e == writeAddrPRF_exec1Addr | _GEN_6274;
    end else begin
      PRFValidList_62 <= _GEN_6274;
    end
    if (reset) begin // @[decode.scala 199:29]
      PRFValidList_63 <= 1'h0; // @[decode.scala 199:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 786:33]
      PRFValidList_63 <= 6'h3f == writeAddrPRF_exec3Addr | _GEN_13227;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 785:33]
      PRFValidList_63 <= 6'h3f == writeAddrPRF_exec2Addr | _GEN_13099;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 784:33]
      PRFValidList_63 <= 6'h3f == writeAddrPRF_exec1Addr | _GEN_6275;
    end else begin
      PRFValidList_63 <= _GEN_6275;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_31 <= 6'h1f; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_31 <= reservedRegMap1_31; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_31 <= architecturalRegMap_31; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_31 <= _GEN_1201;
      end
    end else begin
      frontEndRegMap_31 <= _GEN_1201;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_30 <= 6'h1e; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_30 <= reservedRegMap1_30; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_30 <= architecturalRegMap_30; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_30 <= _GEN_1200;
      end
    end else begin
      frontEndRegMap_30 <= _GEN_1200;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_29 <= 6'h1d; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_29 <= reservedRegMap1_29; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_29 <= architecturalRegMap_29; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_29 <= _GEN_1199;
      end
    end else begin
      frontEndRegMap_29 <= _GEN_1199;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_28 <= 6'h1c; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_28 <= reservedRegMap1_28; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_28 <= architecturalRegMap_28; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_28 <= _GEN_1198;
      end
    end else begin
      frontEndRegMap_28 <= _GEN_1198;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_27 <= 6'h1b; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_27 <= reservedRegMap1_27; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_27 <= architecturalRegMap_27; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_27 <= _GEN_1197;
      end
    end else begin
      frontEndRegMap_27 <= _GEN_1197;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_26 <= 6'h1a; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_26 <= reservedRegMap1_26; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_26 <= architecturalRegMap_26; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_26 <= _GEN_1196;
      end
    end else begin
      frontEndRegMap_26 <= _GEN_1196;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_25 <= 6'h19; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_25 <= reservedRegMap1_25; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_25 <= architecturalRegMap_25; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_25 <= _GEN_1195;
      end
    end else begin
      frontEndRegMap_25 <= _GEN_1195;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_24 <= 6'h18; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_24 <= reservedRegMap1_24; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_24 <= architecturalRegMap_24; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_24 <= _GEN_1194;
      end
    end else begin
      frontEndRegMap_24 <= _GEN_1194;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_23 <= 6'h17; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_23 <= reservedRegMap1_23; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_23 <= architecturalRegMap_23; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_23 <= _GEN_1193;
      end
    end else begin
      frontEndRegMap_23 <= _GEN_1193;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_22 <= 6'h16; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_22 <= reservedRegMap1_22; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_22 <= architecturalRegMap_22; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_22 <= _GEN_1192;
      end
    end else begin
      frontEndRegMap_22 <= _GEN_1192;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_21 <= 6'h15; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_21 <= reservedRegMap1_21; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_21 <= architecturalRegMap_21; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_21 <= _GEN_1191;
      end
    end else begin
      frontEndRegMap_21 <= _GEN_1191;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_20 <= 6'h14; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_20 <= reservedRegMap1_20; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_20 <= architecturalRegMap_20; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_20 <= _GEN_1190;
      end
    end else begin
      frontEndRegMap_20 <= _GEN_1190;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_19 <= 6'h13; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_19 <= reservedRegMap1_19; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_19 <= architecturalRegMap_19; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_19 <= _GEN_1189;
      end
    end else begin
      frontEndRegMap_19 <= _GEN_1189;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_18 <= 6'h12; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_18 <= reservedRegMap1_18; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_18 <= architecturalRegMap_18; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_18 <= _GEN_1188;
      end
    end else begin
      frontEndRegMap_18 <= _GEN_1188;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_17 <= 6'h11; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_17 <= reservedRegMap1_17; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_17 <= architecturalRegMap_17; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_17 <= _GEN_1187;
      end
    end else begin
      frontEndRegMap_17 <= _GEN_1187;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_16 <= 6'h10; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_16 <= reservedRegMap1_16; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_16 <= architecturalRegMap_16; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_16 <= _GEN_1186;
      end
    end else begin
      frontEndRegMap_16 <= _GEN_1186;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_15 <= 6'hf; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_15 <= reservedRegMap1_15; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_15 <= architecturalRegMap_15; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_15 <= _GEN_1185;
      end
    end else begin
      frontEndRegMap_15 <= _GEN_1185;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_14 <= 6'he; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_14 <= reservedRegMap1_14; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_14 <= architecturalRegMap_14; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_14 <= _GEN_1184;
      end
    end else begin
      frontEndRegMap_14 <= _GEN_1184;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_13 <= 6'hd; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_13 <= reservedRegMap1_13; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_13 <= architecturalRegMap_13; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_13 <= _GEN_1183;
      end
    end else begin
      frontEndRegMap_13 <= _GEN_1183;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_12 <= 6'hc; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_12 <= reservedRegMap1_12; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_12 <= architecturalRegMap_12; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_12 <= _GEN_1182;
      end
    end else begin
      frontEndRegMap_12 <= _GEN_1182;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_11 <= 6'hb; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_11 <= reservedRegMap1_11; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_11 <= architecturalRegMap_11; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_11 <= _GEN_1181;
      end
    end else begin
      frontEndRegMap_11 <= _GEN_1181;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_10 <= 6'ha; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_10 <= reservedRegMap1_10; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_10 <= architecturalRegMap_10; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_10 <= _GEN_1180;
      end
    end else begin
      frontEndRegMap_10 <= _GEN_1180;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_9 <= 6'h9; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_9 <= reservedRegMap1_9; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_9 <= architecturalRegMap_9; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_9 <= _GEN_1179;
      end
    end else begin
      frontEndRegMap_9 <= _GEN_1179;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_8 <= 6'h8; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_8 <= reservedRegMap1_8; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_8 <= architecturalRegMap_8; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_8 <= _GEN_1178;
      end
    end else begin
      frontEndRegMap_8 <= _GEN_1178;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_7 <= 6'h7; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_7 <= reservedRegMap1_7; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_7 <= architecturalRegMap_7; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_7 <= _GEN_1177;
      end
    end else begin
      frontEndRegMap_7 <= _GEN_1177;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_6 <= 6'h6; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_6 <= reservedRegMap1_6; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_6 <= architecturalRegMap_6; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_6 <= _GEN_1176;
      end
    end else begin
      frontEndRegMap_6 <= _GEN_1176;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_5 <= 6'h5; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_5 <= reservedRegMap1_5; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_5 <= architecturalRegMap_5; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_5 <= _GEN_1175;
      end
    end else begin
      frontEndRegMap_5 <= _GEN_1175;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_4 <= 6'h4; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_4 <= reservedRegMap1_4; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_4 <= architecturalRegMap_4; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_4 <= _GEN_1174;
      end
    end else begin
      frontEndRegMap_4 <= _GEN_1174;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_3 <= 6'h3; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_3 <= reservedRegMap1_3; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_3 <= architecturalRegMap_3; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_3 <= _GEN_1173;
      end
    end else begin
      frontEndRegMap_3 <= _GEN_1173;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_2 <= 6'h2; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_2 <= reservedRegMap1_2; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_2 <= architecturalRegMap_2; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_2 <= _GEN_1172;
      end
    end else begin
      frontEndRegMap_2 <= _GEN_1172;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_1 <= 6'h1; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_1 <= reservedRegMap1_1; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_1 <= architecturalRegMap_1; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_1 <= _GEN_1171;
      end
    end else begin
      frontEndRegMap_1 <= _GEN_1171;
    end
    if (reset) begin // @[decode.scala 308:36]
      frontEndRegMap_0 <= 6'h0; // @[decode.scala 308:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        if (|branchEvalIn_branchMask[3:0]) begin // @[decode.scala 381:45]
          frontEndRegMap_0 <= reservedRegMap1_0; // @[decode.scala 382:22]
        end else begin
          frontEndRegMap_0 <= architecturalRegMap_0; // @[decode.scala 386:24]
        end
      end else begin
        frontEndRegMap_0 <= _GEN_1170;
      end
    end else begin
      frontEndRegMap_0 <= _GEN_1170;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_0 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_0 <= _GEN_13463;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_0 <= _GEN_5330;
      end else begin
        PRFFreeList_0 <= _GEN_1042;
      end
    end else begin
      PRFFreeList_0 <= _GEN_1042;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_1 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_1 <= _GEN_13464;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_1 <= _GEN_5331;
      end else begin
        PRFFreeList_1 <= _GEN_1043;
      end
    end else begin
      PRFFreeList_1 <= _GEN_1043;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_2 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_2 <= _GEN_13465;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_2 <= _GEN_5332;
      end else begin
        PRFFreeList_2 <= _GEN_1044;
      end
    end else begin
      PRFFreeList_2 <= _GEN_1044;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_3 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_3 <= _GEN_13466;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_3 <= _GEN_5333;
      end else begin
        PRFFreeList_3 <= _GEN_1045;
      end
    end else begin
      PRFFreeList_3 <= _GEN_1045;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_4 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_4 <= _GEN_13467;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_4 <= _GEN_5334;
      end else begin
        PRFFreeList_4 <= _GEN_1046;
      end
    end else begin
      PRFFreeList_4 <= _GEN_1046;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_5 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_5 <= _GEN_13468;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_5 <= _GEN_5335;
      end else begin
        PRFFreeList_5 <= _GEN_1047;
      end
    end else begin
      PRFFreeList_5 <= _GEN_1047;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_6 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_6 <= _GEN_13469;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_6 <= _GEN_5336;
      end else begin
        PRFFreeList_6 <= _GEN_1048;
      end
    end else begin
      PRFFreeList_6 <= _GEN_1048;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_7 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_7 <= _GEN_13470;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_7 <= _GEN_5337;
      end else begin
        PRFFreeList_7 <= _GEN_1049;
      end
    end else begin
      PRFFreeList_7 <= _GEN_1049;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_8 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_8 <= _GEN_13471;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_8 <= _GEN_5338;
      end else begin
        PRFFreeList_8 <= _GEN_1050;
      end
    end else begin
      PRFFreeList_8 <= _GEN_1050;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_9 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_9 <= _GEN_13472;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_9 <= _GEN_5339;
      end else begin
        PRFFreeList_9 <= _GEN_1051;
      end
    end else begin
      PRFFreeList_9 <= _GEN_1051;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_10 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_10 <= _GEN_13473;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_10 <= _GEN_5340;
      end else begin
        PRFFreeList_10 <= _GEN_1052;
      end
    end else begin
      PRFFreeList_10 <= _GEN_1052;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_11 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_11 <= _GEN_13474;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_11 <= _GEN_5341;
      end else begin
        PRFFreeList_11 <= _GEN_1053;
      end
    end else begin
      PRFFreeList_11 <= _GEN_1053;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_12 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_12 <= _GEN_13475;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_12 <= _GEN_5342;
      end else begin
        PRFFreeList_12 <= _GEN_1054;
      end
    end else begin
      PRFFreeList_12 <= _GEN_1054;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_13 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_13 <= _GEN_13476;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_13 <= _GEN_5343;
      end else begin
        PRFFreeList_13 <= _GEN_1055;
      end
    end else begin
      PRFFreeList_13 <= _GEN_1055;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_14 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_14 <= _GEN_13477;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_14 <= _GEN_5344;
      end else begin
        PRFFreeList_14 <= _GEN_1056;
      end
    end else begin
      PRFFreeList_14 <= _GEN_1056;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_15 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_15 <= _GEN_13478;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_15 <= _GEN_5345;
      end else begin
        PRFFreeList_15 <= _GEN_1057;
      end
    end else begin
      PRFFreeList_15 <= _GEN_1057;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_16 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_16 <= _GEN_13479;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_16 <= _GEN_5346;
      end else begin
        PRFFreeList_16 <= _GEN_1058;
      end
    end else begin
      PRFFreeList_16 <= _GEN_1058;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_17 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_17 <= _GEN_13480;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_17 <= _GEN_5347;
      end else begin
        PRFFreeList_17 <= _GEN_1059;
      end
    end else begin
      PRFFreeList_17 <= _GEN_1059;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_18 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_18 <= _GEN_13481;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_18 <= _GEN_5348;
      end else begin
        PRFFreeList_18 <= _GEN_1060;
      end
    end else begin
      PRFFreeList_18 <= _GEN_1060;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_19 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_19 <= _GEN_13482;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_19 <= _GEN_5349;
      end else begin
        PRFFreeList_19 <= _GEN_1061;
      end
    end else begin
      PRFFreeList_19 <= _GEN_1061;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_20 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_20 <= _GEN_13483;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_20 <= _GEN_5350;
      end else begin
        PRFFreeList_20 <= _GEN_1062;
      end
    end else begin
      PRFFreeList_20 <= _GEN_1062;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_21 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_21 <= _GEN_13484;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_21 <= _GEN_5351;
      end else begin
        PRFFreeList_21 <= _GEN_1063;
      end
    end else begin
      PRFFreeList_21 <= _GEN_1063;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_22 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_22 <= _GEN_13485;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_22 <= _GEN_5352;
      end else begin
        PRFFreeList_22 <= _GEN_1064;
      end
    end else begin
      PRFFreeList_22 <= _GEN_1064;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_23 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_23 <= _GEN_13486;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_23 <= _GEN_5353;
      end else begin
        PRFFreeList_23 <= _GEN_1065;
      end
    end else begin
      PRFFreeList_23 <= _GEN_1065;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_24 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_24 <= _GEN_13487;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_24 <= _GEN_5354;
      end else begin
        PRFFreeList_24 <= _GEN_1066;
      end
    end else begin
      PRFFreeList_24 <= _GEN_1066;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_25 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_25 <= _GEN_13488;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_25 <= _GEN_5355;
      end else begin
        PRFFreeList_25 <= _GEN_1067;
      end
    end else begin
      PRFFreeList_25 <= _GEN_1067;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_26 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_26 <= _GEN_13489;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_26 <= _GEN_5356;
      end else begin
        PRFFreeList_26 <= _GEN_1068;
      end
    end else begin
      PRFFreeList_26 <= _GEN_1068;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_27 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_27 <= _GEN_13490;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_27 <= _GEN_5357;
      end else begin
        PRFFreeList_27 <= _GEN_1069;
      end
    end else begin
      PRFFreeList_27 <= _GEN_1069;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_28 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_28 <= _GEN_13491;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_28 <= _GEN_5358;
      end else begin
        PRFFreeList_28 <= _GEN_1070;
      end
    end else begin
      PRFFreeList_28 <= _GEN_1070;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_29 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_29 <= _GEN_13492;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_29 <= _GEN_5359;
      end else begin
        PRFFreeList_29 <= _GEN_1071;
      end
    end else begin
      PRFFreeList_29 <= _GEN_1071;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_30 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_30 <= _GEN_13493;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_30 <= _GEN_5360;
      end else begin
        PRFFreeList_30 <= _GEN_1072;
      end
    end else begin
      PRFFreeList_30 <= _GEN_1072;
    end
    if (reset) begin // @[decode.scala 310:36]
      PRFFreeList_31 <= 1'h0; // @[decode.scala 310:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      PRFFreeList_31 <= _GEN_13494;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        PRFFreeList_31 <= _GEN_5361;
      end else begin
        PRFFreeList_31 <= _GEN_1073;
      end
    end else begin
      PRFFreeList_31 <= _GEN_1073;
    end
    PRFFreeList_32 <= reset | _GEN_13847; // @[decode.scala 310:{36,36}]
    PRFFreeList_33 <= reset | _GEN_13848; // @[decode.scala 310:{36,36}]
    PRFFreeList_34 <= reset | _GEN_13849; // @[decode.scala 310:{36,36}]
    PRFFreeList_35 <= reset | _GEN_13850; // @[decode.scala 310:{36,36}]
    PRFFreeList_36 <= reset | _GEN_13851; // @[decode.scala 310:{36,36}]
    PRFFreeList_37 <= reset | _GEN_13852; // @[decode.scala 310:{36,36}]
    PRFFreeList_38 <= reset | _GEN_13853; // @[decode.scala 310:{36,36}]
    PRFFreeList_39 <= reset | _GEN_13854; // @[decode.scala 310:{36,36}]
    PRFFreeList_40 <= reset | _GEN_13855; // @[decode.scala 310:{36,36}]
    PRFFreeList_41 <= reset | _GEN_13856; // @[decode.scala 310:{36,36}]
    PRFFreeList_42 <= reset | _GEN_13857; // @[decode.scala 310:{36,36}]
    PRFFreeList_43 <= reset | _GEN_13858; // @[decode.scala 310:{36,36}]
    PRFFreeList_44 <= reset | _GEN_13859; // @[decode.scala 310:{36,36}]
    PRFFreeList_45 <= reset | _GEN_13860; // @[decode.scala 310:{36,36}]
    PRFFreeList_46 <= reset | _GEN_13861; // @[decode.scala 310:{36,36}]
    PRFFreeList_47 <= reset | _GEN_13862; // @[decode.scala 310:{36,36}]
    PRFFreeList_48 <= reset | _GEN_13863; // @[decode.scala 310:{36,36}]
    PRFFreeList_49 <= reset | _GEN_13864; // @[decode.scala 310:{36,36}]
    PRFFreeList_50 <= reset | _GEN_13865; // @[decode.scala 310:{36,36}]
    PRFFreeList_51 <= reset | _GEN_13866; // @[decode.scala 310:{36,36}]
    PRFFreeList_52 <= reset | _GEN_13867; // @[decode.scala 310:{36,36}]
    PRFFreeList_53 <= reset | _GEN_13868; // @[decode.scala 310:{36,36}]
    PRFFreeList_54 <= reset | _GEN_13869; // @[decode.scala 310:{36,36}]
    PRFFreeList_55 <= reset | _GEN_13870; // @[decode.scala 310:{36,36}]
    PRFFreeList_56 <= reset | _GEN_13871; // @[decode.scala 310:{36,36}]
    PRFFreeList_57 <= reset | _GEN_13872; // @[decode.scala 310:{36,36}]
    PRFFreeList_58 <= reset | _GEN_13873; // @[decode.scala 310:{36,36}]
    PRFFreeList_59 <= reset | _GEN_13874; // @[decode.scala 310:{36,36}]
    PRFFreeList_60 <= reset | _GEN_13875; // @[decode.scala 310:{36,36}]
    PRFFreeList_61 <= reset | _GEN_13876; // @[decode.scala 310:{36,36}]
    PRFFreeList_62 <= reset | _GEN_13877; // @[decode.scala 310:{36,36}]
    if (reset) begin // @[decode.scala 225:29]
      branchPCMask <= 5'h0; // @[decode.scala 225:29]
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (_GEN_16095) begin // @[decode.scala 424:27]
          branchPCMask <= 5'h1; // @[decode.scala 425:32]
        end else begin
          branchPCMask <= _GEN_6764;
        end
      end
    end
    if (reset) begin // @[decode.scala 226:29]
      branchReg <= 1'h0; // @[decode.scala 226:29]
    end else if (_T_3) begin // @[decode.scala 419:41]
      branchReg <= _T_191;
    end else if (branchEvalIn_fired) begin // @[decode.scala 363:28]
      if (_T_434) begin // @[decode.scala 369:34]
        branchReg <= 1'h0; // @[decode.scala 370:17]
      end
    end
    if (reset) begin // @[decode.scala 240:31]
      csrReadDataReg <= 64'h0; // @[decode.scala 240:31]
    end else if (opcode == 7'h73 & fun3 != 3'h0 & validInputBuf & readyOutputBuf) begin // @[decode.scala 534:80]
      if (64'h0 == _T_229) begin // @[decode.scala 535:34]
        csrReadDataReg <= ustatus; // @[decode.scala 536:37]
      end else if (64'h5 == _T_229) begin // @[decode.scala 535:34]
        csrReadDataReg <= utvec; // @[decode.scala 537:37]
      end else begin
        csrReadDataReg <= _GEN_10975;
      end
    end
    csrAddrReg <= _GEN_16609[11:0]; // @[decode.scala 242:{27,27}]
    if (reset) begin // @[decode.scala 243:26]
      csrImmReg <= 64'h0; // @[decode.scala 243:26]
    end else if (isCSR) begin // @[decode.scala 525:15]
      csrImmReg <= {{59'd0}, outputBuffer_instruction[19:15]}; // @[decode.scala 529:19]
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_0 <= 6'h0; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h0 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_0 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_1 <= 6'h1; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h1 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_1 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_2 <= 6'h2; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h2 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_2 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_3 <= 6'h3; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h3 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_3 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_4 <= 6'h4; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h4 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_4 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_5 <= 6'h5; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h5 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_5 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_6 <= 6'h6; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h6 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_6 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_7 <= 6'h7; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h7 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_7 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_8 <= 6'h8; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h8 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_8 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_9 <= 6'h9; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h9 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_9 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_10 <= 6'ha; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'ha == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_10 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_11 <= 6'hb; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'hb == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_11 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_12 <= 6'hc; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'hc == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_12 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_13 <= 6'hd; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'hd == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_13 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_14 <= 6'he; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'he == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_14 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_15 <= 6'hf; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'hf == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_15 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_16 <= 6'h10; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h10 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_16 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_17 <= 6'h11; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h11 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_17 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_18 <= 6'h12; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h12 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_18 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_19 <= 6'h13; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h13 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_19 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_20 <= 6'h14; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h14 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_20 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_21 <= 6'h15; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h15 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_21 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_22 <= 6'h16; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h16 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_22 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_23 <= 6'h17; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h17 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_23 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_24 <= 6'h18; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h18 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_24 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_25 <= 6'h19; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h19 == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_25 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_26 <= 6'h1a; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h1a == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_26 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_27 <= 6'h1b; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h1b == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_27 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_28 <= 6'h1c; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h1c == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_28 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_29 <= 6'h1d; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h1d == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_29 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_30 <= 6'h1e; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h1e == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_30 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (reset) begin // @[decode.scala 309:36]
      architecturalRegMap_31 <= 6'h1f; // @[decode.scala 309:36]
    end else if (_T_474) begin // @[decode.scala 889:5]
      if (5'h1f == writeBackResult_rdAddr) begin // @[decode.scala 890:62]
        architecturalRegMap_31 <= writeBackResult_PRFDest; // @[decode.scala 890:62]
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_0 <= _GEN_850;
          end else begin
            reservedRegMap1_0 <= frontEndRegMap_0; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_0 <= _GEN_6277;
        end
      end else begin
        reservedRegMap1_0 <= _GEN_6277;
      end
    end else begin
      reservedRegMap1_0 <= _GEN_6277;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_1 <= _GEN_851;
          end else begin
            reservedRegMap1_1 <= frontEndRegMap_1; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_1 <= _GEN_6278;
        end
      end else begin
        reservedRegMap1_1 <= _GEN_6278;
      end
    end else begin
      reservedRegMap1_1 <= _GEN_6278;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_2 <= _GEN_852;
          end else begin
            reservedRegMap1_2 <= frontEndRegMap_2; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_2 <= _GEN_6279;
        end
      end else begin
        reservedRegMap1_2 <= _GEN_6279;
      end
    end else begin
      reservedRegMap1_2 <= _GEN_6279;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_3 <= _GEN_853;
          end else begin
            reservedRegMap1_3 <= frontEndRegMap_3; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_3 <= _GEN_6280;
        end
      end else begin
        reservedRegMap1_3 <= _GEN_6280;
      end
    end else begin
      reservedRegMap1_3 <= _GEN_6280;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_4 <= _GEN_854;
          end else begin
            reservedRegMap1_4 <= frontEndRegMap_4; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_4 <= _GEN_6281;
        end
      end else begin
        reservedRegMap1_4 <= _GEN_6281;
      end
    end else begin
      reservedRegMap1_4 <= _GEN_6281;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_5 <= _GEN_855;
          end else begin
            reservedRegMap1_5 <= frontEndRegMap_5; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_5 <= _GEN_6282;
        end
      end else begin
        reservedRegMap1_5 <= _GEN_6282;
      end
    end else begin
      reservedRegMap1_5 <= _GEN_6282;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_6 <= _GEN_856;
          end else begin
            reservedRegMap1_6 <= frontEndRegMap_6; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_6 <= _GEN_6283;
        end
      end else begin
        reservedRegMap1_6 <= _GEN_6283;
      end
    end else begin
      reservedRegMap1_6 <= _GEN_6283;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_7 <= _GEN_857;
          end else begin
            reservedRegMap1_7 <= frontEndRegMap_7; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_7 <= _GEN_6284;
        end
      end else begin
        reservedRegMap1_7 <= _GEN_6284;
      end
    end else begin
      reservedRegMap1_7 <= _GEN_6284;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_8 <= _GEN_858;
          end else begin
            reservedRegMap1_8 <= frontEndRegMap_8; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_8 <= _GEN_6285;
        end
      end else begin
        reservedRegMap1_8 <= _GEN_6285;
      end
    end else begin
      reservedRegMap1_8 <= _GEN_6285;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_9 <= _GEN_859;
          end else begin
            reservedRegMap1_9 <= frontEndRegMap_9; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_9 <= _GEN_6286;
        end
      end else begin
        reservedRegMap1_9 <= _GEN_6286;
      end
    end else begin
      reservedRegMap1_9 <= _GEN_6286;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_10 <= _GEN_860;
          end else begin
            reservedRegMap1_10 <= frontEndRegMap_10; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_10 <= _GEN_6287;
        end
      end else begin
        reservedRegMap1_10 <= _GEN_6287;
      end
    end else begin
      reservedRegMap1_10 <= _GEN_6287;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_11 <= _GEN_861;
          end else begin
            reservedRegMap1_11 <= frontEndRegMap_11; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_11 <= _GEN_6288;
        end
      end else begin
        reservedRegMap1_11 <= _GEN_6288;
      end
    end else begin
      reservedRegMap1_11 <= _GEN_6288;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_12 <= _GEN_862;
          end else begin
            reservedRegMap1_12 <= frontEndRegMap_12; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_12 <= _GEN_6289;
        end
      end else begin
        reservedRegMap1_12 <= _GEN_6289;
      end
    end else begin
      reservedRegMap1_12 <= _GEN_6289;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_13 <= _GEN_863;
          end else begin
            reservedRegMap1_13 <= frontEndRegMap_13; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_13 <= _GEN_6290;
        end
      end else begin
        reservedRegMap1_13 <= _GEN_6290;
      end
    end else begin
      reservedRegMap1_13 <= _GEN_6290;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_14 <= _GEN_864;
          end else begin
            reservedRegMap1_14 <= frontEndRegMap_14; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_14 <= _GEN_6291;
        end
      end else begin
        reservedRegMap1_14 <= _GEN_6291;
      end
    end else begin
      reservedRegMap1_14 <= _GEN_6291;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_15 <= _GEN_865;
          end else begin
            reservedRegMap1_15 <= frontEndRegMap_15; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_15 <= _GEN_6292;
        end
      end else begin
        reservedRegMap1_15 <= _GEN_6292;
      end
    end else begin
      reservedRegMap1_15 <= _GEN_6292;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_16 <= _GEN_866;
          end else begin
            reservedRegMap1_16 <= frontEndRegMap_16; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_16 <= _GEN_6293;
        end
      end else begin
        reservedRegMap1_16 <= _GEN_6293;
      end
    end else begin
      reservedRegMap1_16 <= _GEN_6293;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_17 <= _GEN_867;
          end else begin
            reservedRegMap1_17 <= frontEndRegMap_17; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_17 <= _GEN_6294;
        end
      end else begin
        reservedRegMap1_17 <= _GEN_6294;
      end
    end else begin
      reservedRegMap1_17 <= _GEN_6294;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_18 <= _GEN_868;
          end else begin
            reservedRegMap1_18 <= frontEndRegMap_18; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_18 <= _GEN_6295;
        end
      end else begin
        reservedRegMap1_18 <= _GEN_6295;
      end
    end else begin
      reservedRegMap1_18 <= _GEN_6295;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_19 <= _GEN_869;
          end else begin
            reservedRegMap1_19 <= frontEndRegMap_19; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_19 <= _GEN_6296;
        end
      end else begin
        reservedRegMap1_19 <= _GEN_6296;
      end
    end else begin
      reservedRegMap1_19 <= _GEN_6296;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_20 <= _GEN_870;
          end else begin
            reservedRegMap1_20 <= frontEndRegMap_20; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_20 <= _GEN_6297;
        end
      end else begin
        reservedRegMap1_20 <= _GEN_6297;
      end
    end else begin
      reservedRegMap1_20 <= _GEN_6297;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_21 <= _GEN_871;
          end else begin
            reservedRegMap1_21 <= frontEndRegMap_21; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_21 <= _GEN_6298;
        end
      end else begin
        reservedRegMap1_21 <= _GEN_6298;
      end
    end else begin
      reservedRegMap1_21 <= _GEN_6298;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_22 <= _GEN_872;
          end else begin
            reservedRegMap1_22 <= frontEndRegMap_22; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_22 <= _GEN_6299;
        end
      end else begin
        reservedRegMap1_22 <= _GEN_6299;
      end
    end else begin
      reservedRegMap1_22 <= _GEN_6299;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_23 <= _GEN_873;
          end else begin
            reservedRegMap1_23 <= frontEndRegMap_23; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_23 <= _GEN_6300;
        end
      end else begin
        reservedRegMap1_23 <= _GEN_6300;
      end
    end else begin
      reservedRegMap1_23 <= _GEN_6300;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_24 <= _GEN_874;
          end else begin
            reservedRegMap1_24 <= frontEndRegMap_24; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_24 <= _GEN_6301;
        end
      end else begin
        reservedRegMap1_24 <= _GEN_6301;
      end
    end else begin
      reservedRegMap1_24 <= _GEN_6301;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_25 <= _GEN_875;
          end else begin
            reservedRegMap1_25 <= frontEndRegMap_25; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_25 <= _GEN_6302;
        end
      end else begin
        reservedRegMap1_25 <= _GEN_6302;
      end
    end else begin
      reservedRegMap1_25 <= _GEN_6302;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_26 <= _GEN_876;
          end else begin
            reservedRegMap1_26 <= frontEndRegMap_26; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_26 <= _GEN_6303;
        end
      end else begin
        reservedRegMap1_26 <= _GEN_6303;
      end
    end else begin
      reservedRegMap1_26 <= _GEN_6303;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_27 <= _GEN_877;
          end else begin
            reservedRegMap1_27 <= frontEndRegMap_27; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_27 <= _GEN_6304;
        end
      end else begin
        reservedRegMap1_27 <= _GEN_6304;
      end
    end else begin
      reservedRegMap1_27 <= _GEN_6304;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_28 <= _GEN_878;
          end else begin
            reservedRegMap1_28 <= frontEndRegMap_28; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_28 <= _GEN_6305;
        end
      end else begin
        reservedRegMap1_28 <= _GEN_6305;
      end
    end else begin
      reservedRegMap1_28 <= _GEN_6305;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_29 <= _GEN_879;
          end else begin
            reservedRegMap1_29 <= frontEndRegMap_29; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_29 <= _GEN_6306;
        end
      end else begin
        reservedRegMap1_29 <= _GEN_6306;
      end
    end else begin
      reservedRegMap1_29 <= _GEN_6306;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_30 <= _GEN_880;
          end else begin
            reservedRegMap1_30 <= frontEndRegMap_30; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_30 <= _GEN_6307;
        end
      end else begin
        reservedRegMap1_30 <= _GEN_6307;
      end
    end else begin
      reservedRegMap1_30 <= _GEN_6307;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedRegMap1_31 <= _GEN_881;
          end else begin
            reservedRegMap1_31 <= frontEndRegMap_31; // @[decode.scala 433:30]
          end
        end else begin
          reservedRegMap1_31 <= _GEN_6308;
        end
      end else begin
        reservedRegMap1_31 <= _GEN_6308;
      end
    end else begin
      reservedRegMap1_31 <= _GEN_6308;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_0 <= _GEN_6309;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_0 <= _GEN_6926;
        end else begin
          reservedRegMap2_0 <= _GEN_6309;
        end
      end else begin
        reservedRegMap2_0 <= _GEN_6309;
      end
    end else begin
      reservedRegMap2_0 <= _GEN_6309;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_1 <= _GEN_6310;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_1 <= _GEN_6927;
        end else begin
          reservedRegMap2_1 <= _GEN_6310;
        end
      end else begin
        reservedRegMap2_1 <= _GEN_6310;
      end
    end else begin
      reservedRegMap2_1 <= _GEN_6310;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_2 <= _GEN_6311;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_2 <= _GEN_6928;
        end else begin
          reservedRegMap2_2 <= _GEN_6311;
        end
      end else begin
        reservedRegMap2_2 <= _GEN_6311;
      end
    end else begin
      reservedRegMap2_2 <= _GEN_6311;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_3 <= _GEN_6312;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_3 <= _GEN_6929;
        end else begin
          reservedRegMap2_3 <= _GEN_6312;
        end
      end else begin
        reservedRegMap2_3 <= _GEN_6312;
      end
    end else begin
      reservedRegMap2_3 <= _GEN_6312;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_4 <= _GEN_6313;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_4 <= _GEN_6930;
        end else begin
          reservedRegMap2_4 <= _GEN_6313;
        end
      end else begin
        reservedRegMap2_4 <= _GEN_6313;
      end
    end else begin
      reservedRegMap2_4 <= _GEN_6313;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_5 <= _GEN_6314;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_5 <= _GEN_6931;
        end else begin
          reservedRegMap2_5 <= _GEN_6314;
        end
      end else begin
        reservedRegMap2_5 <= _GEN_6314;
      end
    end else begin
      reservedRegMap2_5 <= _GEN_6314;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_6 <= _GEN_6315;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_6 <= _GEN_6932;
        end else begin
          reservedRegMap2_6 <= _GEN_6315;
        end
      end else begin
        reservedRegMap2_6 <= _GEN_6315;
      end
    end else begin
      reservedRegMap2_6 <= _GEN_6315;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_7 <= _GEN_6316;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_7 <= _GEN_6933;
        end else begin
          reservedRegMap2_7 <= _GEN_6316;
        end
      end else begin
        reservedRegMap2_7 <= _GEN_6316;
      end
    end else begin
      reservedRegMap2_7 <= _GEN_6316;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_8 <= _GEN_6317;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_8 <= _GEN_6934;
        end else begin
          reservedRegMap2_8 <= _GEN_6317;
        end
      end else begin
        reservedRegMap2_8 <= _GEN_6317;
      end
    end else begin
      reservedRegMap2_8 <= _GEN_6317;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_9 <= _GEN_6318;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_9 <= _GEN_6935;
        end else begin
          reservedRegMap2_9 <= _GEN_6318;
        end
      end else begin
        reservedRegMap2_9 <= _GEN_6318;
      end
    end else begin
      reservedRegMap2_9 <= _GEN_6318;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_10 <= _GEN_6319;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_10 <= _GEN_6936;
        end else begin
          reservedRegMap2_10 <= _GEN_6319;
        end
      end else begin
        reservedRegMap2_10 <= _GEN_6319;
      end
    end else begin
      reservedRegMap2_10 <= _GEN_6319;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_11 <= _GEN_6320;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_11 <= _GEN_6937;
        end else begin
          reservedRegMap2_11 <= _GEN_6320;
        end
      end else begin
        reservedRegMap2_11 <= _GEN_6320;
      end
    end else begin
      reservedRegMap2_11 <= _GEN_6320;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_12 <= _GEN_6321;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_12 <= _GEN_6938;
        end else begin
          reservedRegMap2_12 <= _GEN_6321;
        end
      end else begin
        reservedRegMap2_12 <= _GEN_6321;
      end
    end else begin
      reservedRegMap2_12 <= _GEN_6321;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_13 <= _GEN_6322;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_13 <= _GEN_6939;
        end else begin
          reservedRegMap2_13 <= _GEN_6322;
        end
      end else begin
        reservedRegMap2_13 <= _GEN_6322;
      end
    end else begin
      reservedRegMap2_13 <= _GEN_6322;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_14 <= _GEN_6323;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_14 <= _GEN_6940;
        end else begin
          reservedRegMap2_14 <= _GEN_6323;
        end
      end else begin
        reservedRegMap2_14 <= _GEN_6323;
      end
    end else begin
      reservedRegMap2_14 <= _GEN_6323;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_15 <= _GEN_6324;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_15 <= _GEN_6941;
        end else begin
          reservedRegMap2_15 <= _GEN_6324;
        end
      end else begin
        reservedRegMap2_15 <= _GEN_6324;
      end
    end else begin
      reservedRegMap2_15 <= _GEN_6324;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_16 <= _GEN_6325;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_16 <= _GEN_6942;
        end else begin
          reservedRegMap2_16 <= _GEN_6325;
        end
      end else begin
        reservedRegMap2_16 <= _GEN_6325;
      end
    end else begin
      reservedRegMap2_16 <= _GEN_6325;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_17 <= _GEN_6326;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_17 <= _GEN_6943;
        end else begin
          reservedRegMap2_17 <= _GEN_6326;
        end
      end else begin
        reservedRegMap2_17 <= _GEN_6326;
      end
    end else begin
      reservedRegMap2_17 <= _GEN_6326;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_18 <= _GEN_6327;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_18 <= _GEN_6944;
        end else begin
          reservedRegMap2_18 <= _GEN_6327;
        end
      end else begin
        reservedRegMap2_18 <= _GEN_6327;
      end
    end else begin
      reservedRegMap2_18 <= _GEN_6327;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_19 <= _GEN_6328;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_19 <= _GEN_6945;
        end else begin
          reservedRegMap2_19 <= _GEN_6328;
        end
      end else begin
        reservedRegMap2_19 <= _GEN_6328;
      end
    end else begin
      reservedRegMap2_19 <= _GEN_6328;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_20 <= _GEN_6329;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_20 <= _GEN_6946;
        end else begin
          reservedRegMap2_20 <= _GEN_6329;
        end
      end else begin
        reservedRegMap2_20 <= _GEN_6329;
      end
    end else begin
      reservedRegMap2_20 <= _GEN_6329;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_21 <= _GEN_6330;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_21 <= _GEN_6947;
        end else begin
          reservedRegMap2_21 <= _GEN_6330;
        end
      end else begin
        reservedRegMap2_21 <= _GEN_6330;
      end
    end else begin
      reservedRegMap2_21 <= _GEN_6330;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_22 <= _GEN_6331;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_22 <= _GEN_6948;
        end else begin
          reservedRegMap2_22 <= _GEN_6331;
        end
      end else begin
        reservedRegMap2_22 <= _GEN_6331;
      end
    end else begin
      reservedRegMap2_22 <= _GEN_6331;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_23 <= _GEN_6332;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_23 <= _GEN_6949;
        end else begin
          reservedRegMap2_23 <= _GEN_6332;
        end
      end else begin
        reservedRegMap2_23 <= _GEN_6332;
      end
    end else begin
      reservedRegMap2_23 <= _GEN_6332;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_24 <= _GEN_6333;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_24 <= _GEN_6950;
        end else begin
          reservedRegMap2_24 <= _GEN_6333;
        end
      end else begin
        reservedRegMap2_24 <= _GEN_6333;
      end
    end else begin
      reservedRegMap2_24 <= _GEN_6333;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_25 <= _GEN_6334;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_25 <= _GEN_6951;
        end else begin
          reservedRegMap2_25 <= _GEN_6334;
        end
      end else begin
        reservedRegMap2_25 <= _GEN_6334;
      end
    end else begin
      reservedRegMap2_25 <= _GEN_6334;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_26 <= _GEN_6335;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_26 <= _GEN_6952;
        end else begin
          reservedRegMap2_26 <= _GEN_6335;
        end
      end else begin
        reservedRegMap2_26 <= _GEN_6335;
      end
    end else begin
      reservedRegMap2_26 <= _GEN_6335;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_27 <= _GEN_6336;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_27 <= _GEN_6953;
        end else begin
          reservedRegMap2_27 <= _GEN_6336;
        end
      end else begin
        reservedRegMap2_27 <= _GEN_6336;
      end
    end else begin
      reservedRegMap2_27 <= _GEN_6336;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_28 <= _GEN_6337;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_28 <= _GEN_6954;
        end else begin
          reservedRegMap2_28 <= _GEN_6337;
        end
      end else begin
        reservedRegMap2_28 <= _GEN_6337;
      end
    end else begin
      reservedRegMap2_28 <= _GEN_6337;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_29 <= _GEN_6338;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_29 <= _GEN_6955;
        end else begin
          reservedRegMap2_29 <= _GEN_6338;
        end
      end else begin
        reservedRegMap2_29 <= _GEN_6338;
      end
    end else begin
      reservedRegMap2_29 <= _GEN_6338;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_30 <= _GEN_6339;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_30 <= _GEN_6956;
        end else begin
          reservedRegMap2_30 <= _GEN_6339;
        end
      end else begin
        reservedRegMap2_30 <= _GEN_6339;
      end
    end else begin
      reservedRegMap2_30 <= _GEN_6339;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_31 <= _GEN_6340;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap2_31 <= _GEN_6957;
        end else begin
          reservedRegMap2_31 <= _GEN_6340;
        end
      end else begin
        reservedRegMap2_31 <= _GEN_6340;
      end
    end else begin
      reservedRegMap2_31 <= _GEN_6340;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_0 <= _GEN_6341;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_0 <= _GEN_6341;
        end else begin
          reservedRegMap3_0 <= _GEN_8206;
        end
      end else begin
        reservedRegMap3_0 <= _GEN_6341;
      end
    end else begin
      reservedRegMap3_0 <= _GEN_6341;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_1 <= _GEN_6342;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_1 <= _GEN_6342;
        end else begin
          reservedRegMap3_1 <= _GEN_8207;
        end
      end else begin
        reservedRegMap3_1 <= _GEN_6342;
      end
    end else begin
      reservedRegMap3_1 <= _GEN_6342;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_2 <= _GEN_6343;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_2 <= _GEN_6343;
        end else begin
          reservedRegMap3_2 <= _GEN_8208;
        end
      end else begin
        reservedRegMap3_2 <= _GEN_6343;
      end
    end else begin
      reservedRegMap3_2 <= _GEN_6343;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_3 <= _GEN_6344;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_3 <= _GEN_6344;
        end else begin
          reservedRegMap3_3 <= _GEN_8209;
        end
      end else begin
        reservedRegMap3_3 <= _GEN_6344;
      end
    end else begin
      reservedRegMap3_3 <= _GEN_6344;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_4 <= _GEN_6345;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_4 <= _GEN_6345;
        end else begin
          reservedRegMap3_4 <= _GEN_8210;
        end
      end else begin
        reservedRegMap3_4 <= _GEN_6345;
      end
    end else begin
      reservedRegMap3_4 <= _GEN_6345;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_5 <= _GEN_6346;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_5 <= _GEN_6346;
        end else begin
          reservedRegMap3_5 <= _GEN_8211;
        end
      end else begin
        reservedRegMap3_5 <= _GEN_6346;
      end
    end else begin
      reservedRegMap3_5 <= _GEN_6346;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_6 <= _GEN_6347;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_6 <= _GEN_6347;
        end else begin
          reservedRegMap3_6 <= _GEN_8212;
        end
      end else begin
        reservedRegMap3_6 <= _GEN_6347;
      end
    end else begin
      reservedRegMap3_6 <= _GEN_6347;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_7 <= _GEN_6348;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_7 <= _GEN_6348;
        end else begin
          reservedRegMap3_7 <= _GEN_8213;
        end
      end else begin
        reservedRegMap3_7 <= _GEN_6348;
      end
    end else begin
      reservedRegMap3_7 <= _GEN_6348;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_8 <= _GEN_6349;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_8 <= _GEN_6349;
        end else begin
          reservedRegMap3_8 <= _GEN_8214;
        end
      end else begin
        reservedRegMap3_8 <= _GEN_6349;
      end
    end else begin
      reservedRegMap3_8 <= _GEN_6349;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_9 <= _GEN_6350;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_9 <= _GEN_6350;
        end else begin
          reservedRegMap3_9 <= _GEN_8215;
        end
      end else begin
        reservedRegMap3_9 <= _GEN_6350;
      end
    end else begin
      reservedRegMap3_9 <= _GEN_6350;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_10 <= _GEN_6351;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_10 <= _GEN_6351;
        end else begin
          reservedRegMap3_10 <= _GEN_8216;
        end
      end else begin
        reservedRegMap3_10 <= _GEN_6351;
      end
    end else begin
      reservedRegMap3_10 <= _GEN_6351;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_11 <= _GEN_6352;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_11 <= _GEN_6352;
        end else begin
          reservedRegMap3_11 <= _GEN_8217;
        end
      end else begin
        reservedRegMap3_11 <= _GEN_6352;
      end
    end else begin
      reservedRegMap3_11 <= _GEN_6352;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_12 <= _GEN_6353;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_12 <= _GEN_6353;
        end else begin
          reservedRegMap3_12 <= _GEN_8218;
        end
      end else begin
        reservedRegMap3_12 <= _GEN_6353;
      end
    end else begin
      reservedRegMap3_12 <= _GEN_6353;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_13 <= _GEN_6354;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_13 <= _GEN_6354;
        end else begin
          reservedRegMap3_13 <= _GEN_8219;
        end
      end else begin
        reservedRegMap3_13 <= _GEN_6354;
      end
    end else begin
      reservedRegMap3_13 <= _GEN_6354;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_14 <= _GEN_6355;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_14 <= _GEN_6355;
        end else begin
          reservedRegMap3_14 <= _GEN_8220;
        end
      end else begin
        reservedRegMap3_14 <= _GEN_6355;
      end
    end else begin
      reservedRegMap3_14 <= _GEN_6355;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_15 <= _GEN_6356;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_15 <= _GEN_6356;
        end else begin
          reservedRegMap3_15 <= _GEN_8221;
        end
      end else begin
        reservedRegMap3_15 <= _GEN_6356;
      end
    end else begin
      reservedRegMap3_15 <= _GEN_6356;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_16 <= _GEN_6357;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_16 <= _GEN_6357;
        end else begin
          reservedRegMap3_16 <= _GEN_8222;
        end
      end else begin
        reservedRegMap3_16 <= _GEN_6357;
      end
    end else begin
      reservedRegMap3_16 <= _GEN_6357;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_17 <= _GEN_6358;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_17 <= _GEN_6358;
        end else begin
          reservedRegMap3_17 <= _GEN_8223;
        end
      end else begin
        reservedRegMap3_17 <= _GEN_6358;
      end
    end else begin
      reservedRegMap3_17 <= _GEN_6358;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_18 <= _GEN_6359;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_18 <= _GEN_6359;
        end else begin
          reservedRegMap3_18 <= _GEN_8224;
        end
      end else begin
        reservedRegMap3_18 <= _GEN_6359;
      end
    end else begin
      reservedRegMap3_18 <= _GEN_6359;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_19 <= _GEN_6360;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_19 <= _GEN_6360;
        end else begin
          reservedRegMap3_19 <= _GEN_8225;
        end
      end else begin
        reservedRegMap3_19 <= _GEN_6360;
      end
    end else begin
      reservedRegMap3_19 <= _GEN_6360;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_20 <= _GEN_6361;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_20 <= _GEN_6361;
        end else begin
          reservedRegMap3_20 <= _GEN_8226;
        end
      end else begin
        reservedRegMap3_20 <= _GEN_6361;
      end
    end else begin
      reservedRegMap3_20 <= _GEN_6361;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_21 <= _GEN_6362;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_21 <= _GEN_6362;
        end else begin
          reservedRegMap3_21 <= _GEN_8227;
        end
      end else begin
        reservedRegMap3_21 <= _GEN_6362;
      end
    end else begin
      reservedRegMap3_21 <= _GEN_6362;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_22 <= _GEN_6363;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_22 <= _GEN_6363;
        end else begin
          reservedRegMap3_22 <= _GEN_8228;
        end
      end else begin
        reservedRegMap3_22 <= _GEN_6363;
      end
    end else begin
      reservedRegMap3_22 <= _GEN_6363;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_23 <= _GEN_6364;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_23 <= _GEN_6364;
        end else begin
          reservedRegMap3_23 <= _GEN_8229;
        end
      end else begin
        reservedRegMap3_23 <= _GEN_6364;
      end
    end else begin
      reservedRegMap3_23 <= _GEN_6364;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_24 <= _GEN_6365;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_24 <= _GEN_6365;
        end else begin
          reservedRegMap3_24 <= _GEN_8230;
        end
      end else begin
        reservedRegMap3_24 <= _GEN_6365;
      end
    end else begin
      reservedRegMap3_24 <= _GEN_6365;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_25 <= _GEN_6366;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_25 <= _GEN_6366;
        end else begin
          reservedRegMap3_25 <= _GEN_8231;
        end
      end else begin
        reservedRegMap3_25 <= _GEN_6366;
      end
    end else begin
      reservedRegMap3_25 <= _GEN_6366;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_26 <= _GEN_6367;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_26 <= _GEN_6367;
        end else begin
          reservedRegMap3_26 <= _GEN_8232;
        end
      end else begin
        reservedRegMap3_26 <= _GEN_6367;
      end
    end else begin
      reservedRegMap3_26 <= _GEN_6367;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_27 <= _GEN_6368;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_27 <= _GEN_6368;
        end else begin
          reservedRegMap3_27 <= _GEN_8233;
        end
      end else begin
        reservedRegMap3_27 <= _GEN_6368;
      end
    end else begin
      reservedRegMap3_27 <= _GEN_6368;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_28 <= _GEN_6369;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_28 <= _GEN_6369;
        end else begin
          reservedRegMap3_28 <= _GEN_8234;
        end
      end else begin
        reservedRegMap3_28 <= _GEN_6369;
      end
    end else begin
      reservedRegMap3_28 <= _GEN_6369;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_29 <= _GEN_6370;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_29 <= _GEN_6370;
        end else begin
          reservedRegMap3_29 <= _GEN_8235;
        end
      end else begin
        reservedRegMap3_29 <= _GEN_6370;
      end
    end else begin
      reservedRegMap3_29 <= _GEN_6370;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_30 <= _GEN_6371;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_30 <= _GEN_6371;
        end else begin
          reservedRegMap3_30 <= _GEN_8236;
        end
      end else begin
        reservedRegMap3_30 <= _GEN_6371;
      end
    end else begin
      reservedRegMap3_30 <= _GEN_6371;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_31 <= _GEN_6372;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedRegMap3_31 <= _GEN_6372;
        end else begin
          reservedRegMap3_31 <= _GEN_8237;
        end
      end else begin
        reservedRegMap3_31 <= _GEN_6372;
      end
    end else begin
      reservedRegMap3_31 <= _GEN_6372;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_0 <= _GEN_8366;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_1 <= _GEN_8367;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_2 <= _GEN_8368;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_3 <= _GEN_8369;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_4 <= _GEN_8370;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_5 <= _GEN_8371;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_6 <= _GEN_8372;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_7 <= _GEN_8373;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_8 <= _GEN_8374;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_9 <= _GEN_8375;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_10 <= _GEN_8376;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_11 <= _GEN_8377;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_12 <= _GEN_8378;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_13 <= _GEN_8379;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_14 <= _GEN_8380;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_15 <= _GEN_8381;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_16 <= _GEN_8382;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_17 <= _GEN_8383;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_18 <= _GEN_8384;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_19 <= _GEN_8385;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_20 <= _GEN_8386;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_21 <= _GEN_8387;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_22 <= _GEN_8388;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_23 <= _GEN_8389;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_24 <= _GEN_8390;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_25 <= _GEN_8391;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_26 <= _GEN_8392;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_27 <= _GEN_8393;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_28 <= _GEN_8394;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_29 <= _GEN_8395;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_30 <= _GEN_8396;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedRegMap4_31 <= _GEN_8397;
          end
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_0 <= _GEN_13527;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_0 <= _GEN_6958;
        end else begin
          reservedFreeList1_0 <= _GEN_6373;
        end
      end else begin
        reservedFreeList1_0 <= _GEN_6373;
      end
    end else begin
      reservedFreeList1_0 <= _GEN_6373;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_1 <= _GEN_13528;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_1 <= _GEN_6959;
        end else begin
          reservedFreeList1_1 <= _GEN_6374;
        end
      end else begin
        reservedFreeList1_1 <= _GEN_6374;
      end
    end else begin
      reservedFreeList1_1 <= _GEN_6374;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_2 <= _GEN_13529;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_2 <= _GEN_6960;
        end else begin
          reservedFreeList1_2 <= _GEN_6375;
        end
      end else begin
        reservedFreeList1_2 <= _GEN_6375;
      end
    end else begin
      reservedFreeList1_2 <= _GEN_6375;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_3 <= _GEN_13530;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_3 <= _GEN_6961;
        end else begin
          reservedFreeList1_3 <= _GEN_6376;
        end
      end else begin
        reservedFreeList1_3 <= _GEN_6376;
      end
    end else begin
      reservedFreeList1_3 <= _GEN_6376;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_4 <= _GEN_13531;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_4 <= _GEN_6962;
        end else begin
          reservedFreeList1_4 <= _GEN_6377;
        end
      end else begin
        reservedFreeList1_4 <= _GEN_6377;
      end
    end else begin
      reservedFreeList1_4 <= _GEN_6377;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_5 <= _GEN_13532;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_5 <= _GEN_6963;
        end else begin
          reservedFreeList1_5 <= _GEN_6378;
        end
      end else begin
        reservedFreeList1_5 <= _GEN_6378;
      end
    end else begin
      reservedFreeList1_5 <= _GEN_6378;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_6 <= _GEN_13533;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_6 <= _GEN_6964;
        end else begin
          reservedFreeList1_6 <= _GEN_6379;
        end
      end else begin
        reservedFreeList1_6 <= _GEN_6379;
      end
    end else begin
      reservedFreeList1_6 <= _GEN_6379;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_7 <= _GEN_13534;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_7 <= _GEN_6965;
        end else begin
          reservedFreeList1_7 <= _GEN_6380;
        end
      end else begin
        reservedFreeList1_7 <= _GEN_6380;
      end
    end else begin
      reservedFreeList1_7 <= _GEN_6380;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_8 <= _GEN_13535;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_8 <= _GEN_6966;
        end else begin
          reservedFreeList1_8 <= _GEN_6381;
        end
      end else begin
        reservedFreeList1_8 <= _GEN_6381;
      end
    end else begin
      reservedFreeList1_8 <= _GEN_6381;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_9 <= _GEN_13536;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_9 <= _GEN_6967;
        end else begin
          reservedFreeList1_9 <= _GEN_6382;
        end
      end else begin
        reservedFreeList1_9 <= _GEN_6382;
      end
    end else begin
      reservedFreeList1_9 <= _GEN_6382;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_10 <= _GEN_13537;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_10 <= _GEN_6968;
        end else begin
          reservedFreeList1_10 <= _GEN_6383;
        end
      end else begin
        reservedFreeList1_10 <= _GEN_6383;
      end
    end else begin
      reservedFreeList1_10 <= _GEN_6383;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_11 <= _GEN_13538;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_11 <= _GEN_6969;
        end else begin
          reservedFreeList1_11 <= _GEN_6384;
        end
      end else begin
        reservedFreeList1_11 <= _GEN_6384;
      end
    end else begin
      reservedFreeList1_11 <= _GEN_6384;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_12 <= _GEN_13539;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_12 <= _GEN_6970;
        end else begin
          reservedFreeList1_12 <= _GEN_6385;
        end
      end else begin
        reservedFreeList1_12 <= _GEN_6385;
      end
    end else begin
      reservedFreeList1_12 <= _GEN_6385;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_13 <= _GEN_13540;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_13 <= _GEN_6971;
        end else begin
          reservedFreeList1_13 <= _GEN_6386;
        end
      end else begin
        reservedFreeList1_13 <= _GEN_6386;
      end
    end else begin
      reservedFreeList1_13 <= _GEN_6386;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_14 <= _GEN_13541;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_14 <= _GEN_6972;
        end else begin
          reservedFreeList1_14 <= _GEN_6387;
        end
      end else begin
        reservedFreeList1_14 <= _GEN_6387;
      end
    end else begin
      reservedFreeList1_14 <= _GEN_6387;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_15 <= _GEN_13542;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_15 <= _GEN_6973;
        end else begin
          reservedFreeList1_15 <= _GEN_6388;
        end
      end else begin
        reservedFreeList1_15 <= _GEN_6388;
      end
    end else begin
      reservedFreeList1_15 <= _GEN_6388;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_16 <= _GEN_13543;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_16 <= _GEN_6974;
        end else begin
          reservedFreeList1_16 <= _GEN_6389;
        end
      end else begin
        reservedFreeList1_16 <= _GEN_6389;
      end
    end else begin
      reservedFreeList1_16 <= _GEN_6389;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_17 <= _GEN_13544;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_17 <= _GEN_6975;
        end else begin
          reservedFreeList1_17 <= _GEN_6390;
        end
      end else begin
        reservedFreeList1_17 <= _GEN_6390;
      end
    end else begin
      reservedFreeList1_17 <= _GEN_6390;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_18 <= _GEN_13545;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_18 <= _GEN_6976;
        end else begin
          reservedFreeList1_18 <= _GEN_6391;
        end
      end else begin
        reservedFreeList1_18 <= _GEN_6391;
      end
    end else begin
      reservedFreeList1_18 <= _GEN_6391;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_19 <= _GEN_13546;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_19 <= _GEN_6977;
        end else begin
          reservedFreeList1_19 <= _GEN_6392;
        end
      end else begin
        reservedFreeList1_19 <= _GEN_6392;
      end
    end else begin
      reservedFreeList1_19 <= _GEN_6392;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_20 <= _GEN_13547;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_20 <= _GEN_6978;
        end else begin
          reservedFreeList1_20 <= _GEN_6393;
        end
      end else begin
        reservedFreeList1_20 <= _GEN_6393;
      end
    end else begin
      reservedFreeList1_20 <= _GEN_6393;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_21 <= _GEN_13548;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_21 <= _GEN_6979;
        end else begin
          reservedFreeList1_21 <= _GEN_6394;
        end
      end else begin
        reservedFreeList1_21 <= _GEN_6394;
      end
    end else begin
      reservedFreeList1_21 <= _GEN_6394;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_22 <= _GEN_13549;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_22 <= _GEN_6980;
        end else begin
          reservedFreeList1_22 <= _GEN_6395;
        end
      end else begin
        reservedFreeList1_22 <= _GEN_6395;
      end
    end else begin
      reservedFreeList1_22 <= _GEN_6395;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_23 <= _GEN_13550;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_23 <= _GEN_6981;
        end else begin
          reservedFreeList1_23 <= _GEN_6396;
        end
      end else begin
        reservedFreeList1_23 <= _GEN_6396;
      end
    end else begin
      reservedFreeList1_23 <= _GEN_6396;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_24 <= _GEN_13551;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_24 <= _GEN_6982;
        end else begin
          reservedFreeList1_24 <= _GEN_6397;
        end
      end else begin
        reservedFreeList1_24 <= _GEN_6397;
      end
    end else begin
      reservedFreeList1_24 <= _GEN_6397;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_25 <= _GEN_13552;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_25 <= _GEN_6983;
        end else begin
          reservedFreeList1_25 <= _GEN_6398;
        end
      end else begin
        reservedFreeList1_25 <= _GEN_6398;
      end
    end else begin
      reservedFreeList1_25 <= _GEN_6398;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_26 <= _GEN_13553;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_26 <= _GEN_6984;
        end else begin
          reservedFreeList1_26 <= _GEN_6399;
        end
      end else begin
        reservedFreeList1_26 <= _GEN_6399;
      end
    end else begin
      reservedFreeList1_26 <= _GEN_6399;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_27 <= _GEN_13554;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_27 <= _GEN_6985;
        end else begin
          reservedFreeList1_27 <= _GEN_6400;
        end
      end else begin
        reservedFreeList1_27 <= _GEN_6400;
      end
    end else begin
      reservedFreeList1_27 <= _GEN_6400;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_28 <= _GEN_13555;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_28 <= _GEN_6986;
        end else begin
          reservedFreeList1_28 <= _GEN_6401;
        end
      end else begin
        reservedFreeList1_28 <= _GEN_6401;
      end
    end else begin
      reservedFreeList1_28 <= _GEN_6401;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_29 <= _GEN_13556;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_29 <= _GEN_6987;
        end else begin
          reservedFreeList1_29 <= _GEN_6402;
        end
      end else begin
        reservedFreeList1_29 <= _GEN_6402;
      end
    end else begin
      reservedFreeList1_29 <= _GEN_6402;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_30 <= _GEN_13557;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_30 <= _GEN_6988;
        end else begin
          reservedFreeList1_30 <= _GEN_6403;
        end
      end else begin
        reservedFreeList1_30 <= _GEN_6403;
      end
    end else begin
      reservedFreeList1_30 <= _GEN_6403;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_31 <= _GEN_13558;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_31 <= _GEN_6989;
        end else begin
          reservedFreeList1_31 <= _GEN_6404;
        end
      end else begin
        reservedFreeList1_31 <= _GEN_6404;
      end
    end else begin
      reservedFreeList1_31 <= _GEN_6404;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_32 <= _GEN_13559;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_32 <= _GEN_6990;
        end else begin
          reservedFreeList1_32 <= _GEN_6405;
        end
      end else begin
        reservedFreeList1_32 <= _GEN_6405;
      end
    end else begin
      reservedFreeList1_32 <= _GEN_6405;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_33 <= _GEN_13560;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_33 <= _GEN_6991;
        end else begin
          reservedFreeList1_33 <= _GEN_6406;
        end
      end else begin
        reservedFreeList1_33 <= _GEN_6406;
      end
    end else begin
      reservedFreeList1_33 <= _GEN_6406;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_34 <= _GEN_13561;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_34 <= _GEN_6992;
        end else begin
          reservedFreeList1_34 <= _GEN_6407;
        end
      end else begin
        reservedFreeList1_34 <= _GEN_6407;
      end
    end else begin
      reservedFreeList1_34 <= _GEN_6407;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_35 <= _GEN_13562;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_35 <= _GEN_6993;
        end else begin
          reservedFreeList1_35 <= _GEN_6408;
        end
      end else begin
        reservedFreeList1_35 <= _GEN_6408;
      end
    end else begin
      reservedFreeList1_35 <= _GEN_6408;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_36 <= _GEN_13563;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_36 <= _GEN_6994;
        end else begin
          reservedFreeList1_36 <= _GEN_6409;
        end
      end else begin
        reservedFreeList1_36 <= _GEN_6409;
      end
    end else begin
      reservedFreeList1_36 <= _GEN_6409;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_37 <= _GEN_13564;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_37 <= _GEN_6995;
        end else begin
          reservedFreeList1_37 <= _GEN_6410;
        end
      end else begin
        reservedFreeList1_37 <= _GEN_6410;
      end
    end else begin
      reservedFreeList1_37 <= _GEN_6410;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_38 <= _GEN_13565;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_38 <= _GEN_6996;
        end else begin
          reservedFreeList1_38 <= _GEN_6411;
        end
      end else begin
        reservedFreeList1_38 <= _GEN_6411;
      end
    end else begin
      reservedFreeList1_38 <= _GEN_6411;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_39 <= _GEN_13566;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_39 <= _GEN_6997;
        end else begin
          reservedFreeList1_39 <= _GEN_6412;
        end
      end else begin
        reservedFreeList1_39 <= _GEN_6412;
      end
    end else begin
      reservedFreeList1_39 <= _GEN_6412;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_40 <= _GEN_13567;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_40 <= _GEN_6998;
        end else begin
          reservedFreeList1_40 <= _GEN_6413;
        end
      end else begin
        reservedFreeList1_40 <= _GEN_6413;
      end
    end else begin
      reservedFreeList1_40 <= _GEN_6413;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_41 <= _GEN_13568;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_41 <= _GEN_6999;
        end else begin
          reservedFreeList1_41 <= _GEN_6414;
        end
      end else begin
        reservedFreeList1_41 <= _GEN_6414;
      end
    end else begin
      reservedFreeList1_41 <= _GEN_6414;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_42 <= _GEN_13569;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_42 <= _GEN_7000;
        end else begin
          reservedFreeList1_42 <= _GEN_6415;
        end
      end else begin
        reservedFreeList1_42 <= _GEN_6415;
      end
    end else begin
      reservedFreeList1_42 <= _GEN_6415;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_43 <= _GEN_13570;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_43 <= _GEN_7001;
        end else begin
          reservedFreeList1_43 <= _GEN_6416;
        end
      end else begin
        reservedFreeList1_43 <= _GEN_6416;
      end
    end else begin
      reservedFreeList1_43 <= _GEN_6416;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_44 <= _GEN_13571;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_44 <= _GEN_7002;
        end else begin
          reservedFreeList1_44 <= _GEN_6417;
        end
      end else begin
        reservedFreeList1_44 <= _GEN_6417;
      end
    end else begin
      reservedFreeList1_44 <= _GEN_6417;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_45 <= _GEN_13572;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_45 <= _GEN_7003;
        end else begin
          reservedFreeList1_45 <= _GEN_6418;
        end
      end else begin
        reservedFreeList1_45 <= _GEN_6418;
      end
    end else begin
      reservedFreeList1_45 <= _GEN_6418;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_46 <= _GEN_13573;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_46 <= _GEN_7004;
        end else begin
          reservedFreeList1_46 <= _GEN_6419;
        end
      end else begin
        reservedFreeList1_46 <= _GEN_6419;
      end
    end else begin
      reservedFreeList1_46 <= _GEN_6419;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_47 <= _GEN_13574;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_47 <= _GEN_7005;
        end else begin
          reservedFreeList1_47 <= _GEN_6420;
        end
      end else begin
        reservedFreeList1_47 <= _GEN_6420;
      end
    end else begin
      reservedFreeList1_47 <= _GEN_6420;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_48 <= _GEN_13575;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_48 <= _GEN_7006;
        end else begin
          reservedFreeList1_48 <= _GEN_6421;
        end
      end else begin
        reservedFreeList1_48 <= _GEN_6421;
      end
    end else begin
      reservedFreeList1_48 <= _GEN_6421;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_49 <= _GEN_13576;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_49 <= _GEN_7007;
        end else begin
          reservedFreeList1_49 <= _GEN_6422;
        end
      end else begin
        reservedFreeList1_49 <= _GEN_6422;
      end
    end else begin
      reservedFreeList1_49 <= _GEN_6422;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_50 <= _GEN_13577;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_50 <= _GEN_7008;
        end else begin
          reservedFreeList1_50 <= _GEN_6423;
        end
      end else begin
        reservedFreeList1_50 <= _GEN_6423;
      end
    end else begin
      reservedFreeList1_50 <= _GEN_6423;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_51 <= _GEN_13578;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_51 <= _GEN_7009;
        end else begin
          reservedFreeList1_51 <= _GEN_6424;
        end
      end else begin
        reservedFreeList1_51 <= _GEN_6424;
      end
    end else begin
      reservedFreeList1_51 <= _GEN_6424;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_52 <= _GEN_13579;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_52 <= _GEN_7010;
        end else begin
          reservedFreeList1_52 <= _GEN_6425;
        end
      end else begin
        reservedFreeList1_52 <= _GEN_6425;
      end
    end else begin
      reservedFreeList1_52 <= _GEN_6425;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_53 <= _GEN_13580;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_53 <= _GEN_7011;
        end else begin
          reservedFreeList1_53 <= _GEN_6426;
        end
      end else begin
        reservedFreeList1_53 <= _GEN_6426;
      end
    end else begin
      reservedFreeList1_53 <= _GEN_6426;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_54 <= _GEN_13581;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_54 <= _GEN_7012;
        end else begin
          reservedFreeList1_54 <= _GEN_6427;
        end
      end else begin
        reservedFreeList1_54 <= _GEN_6427;
      end
    end else begin
      reservedFreeList1_54 <= _GEN_6427;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_55 <= _GEN_13582;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_55 <= _GEN_7013;
        end else begin
          reservedFreeList1_55 <= _GEN_6428;
        end
      end else begin
        reservedFreeList1_55 <= _GEN_6428;
      end
    end else begin
      reservedFreeList1_55 <= _GEN_6428;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_56 <= _GEN_13583;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_56 <= _GEN_7014;
        end else begin
          reservedFreeList1_56 <= _GEN_6429;
        end
      end else begin
        reservedFreeList1_56 <= _GEN_6429;
      end
    end else begin
      reservedFreeList1_56 <= _GEN_6429;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_57 <= _GEN_13584;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_57 <= _GEN_7015;
        end else begin
          reservedFreeList1_57 <= _GEN_6430;
        end
      end else begin
        reservedFreeList1_57 <= _GEN_6430;
      end
    end else begin
      reservedFreeList1_57 <= _GEN_6430;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_58 <= _GEN_13585;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_58 <= _GEN_7016;
        end else begin
          reservedFreeList1_58 <= _GEN_6431;
        end
      end else begin
        reservedFreeList1_58 <= _GEN_6431;
      end
    end else begin
      reservedFreeList1_58 <= _GEN_6431;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_59 <= _GEN_13586;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_59 <= _GEN_7017;
        end else begin
          reservedFreeList1_59 <= _GEN_6432;
        end
      end else begin
        reservedFreeList1_59 <= _GEN_6432;
      end
    end else begin
      reservedFreeList1_59 <= _GEN_6432;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_60 <= _GEN_13587;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_60 <= _GEN_7018;
        end else begin
          reservedFreeList1_60 <= _GEN_6433;
        end
      end else begin
        reservedFreeList1_60 <= _GEN_6433;
      end
    end else begin
      reservedFreeList1_60 <= _GEN_6433;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_61 <= _GEN_13588;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_61 <= _GEN_7019;
        end else begin
          reservedFreeList1_61 <= _GEN_6434;
        end
      end else begin
        reservedFreeList1_61 <= _GEN_6434;
      end
    end else begin
      reservedFreeList1_61 <= _GEN_6434;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList1_62 <= _GEN_13589;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList1_62 <= _GEN_7020;
        end else begin
          reservedFreeList1_62 <= _GEN_6435;
        end
      end else begin
        reservedFreeList1_62 <= _GEN_6435;
      end
    end else begin
      reservedFreeList1_62 <= _GEN_6435;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_0 <= _GEN_13591;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_0 <= _GEN_6437;
        end else begin
          reservedFreeList2_0 <= _GEN_8558;
        end
      end else begin
        reservedFreeList2_0 <= _GEN_6437;
      end
    end else begin
      reservedFreeList2_0 <= _GEN_6437;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_1 <= _GEN_13592;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_1 <= _GEN_6438;
        end else begin
          reservedFreeList2_1 <= _GEN_8559;
        end
      end else begin
        reservedFreeList2_1 <= _GEN_6438;
      end
    end else begin
      reservedFreeList2_1 <= _GEN_6438;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_2 <= _GEN_13593;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_2 <= _GEN_6439;
        end else begin
          reservedFreeList2_2 <= _GEN_8560;
        end
      end else begin
        reservedFreeList2_2 <= _GEN_6439;
      end
    end else begin
      reservedFreeList2_2 <= _GEN_6439;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_3 <= _GEN_13594;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_3 <= _GEN_6440;
        end else begin
          reservedFreeList2_3 <= _GEN_8561;
        end
      end else begin
        reservedFreeList2_3 <= _GEN_6440;
      end
    end else begin
      reservedFreeList2_3 <= _GEN_6440;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_4 <= _GEN_13595;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_4 <= _GEN_6441;
        end else begin
          reservedFreeList2_4 <= _GEN_8562;
        end
      end else begin
        reservedFreeList2_4 <= _GEN_6441;
      end
    end else begin
      reservedFreeList2_4 <= _GEN_6441;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_5 <= _GEN_13596;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_5 <= _GEN_6442;
        end else begin
          reservedFreeList2_5 <= _GEN_8563;
        end
      end else begin
        reservedFreeList2_5 <= _GEN_6442;
      end
    end else begin
      reservedFreeList2_5 <= _GEN_6442;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_6 <= _GEN_13597;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_6 <= _GEN_6443;
        end else begin
          reservedFreeList2_6 <= _GEN_8564;
        end
      end else begin
        reservedFreeList2_6 <= _GEN_6443;
      end
    end else begin
      reservedFreeList2_6 <= _GEN_6443;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_7 <= _GEN_13598;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_7 <= _GEN_6444;
        end else begin
          reservedFreeList2_7 <= _GEN_8565;
        end
      end else begin
        reservedFreeList2_7 <= _GEN_6444;
      end
    end else begin
      reservedFreeList2_7 <= _GEN_6444;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_8 <= _GEN_13599;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_8 <= _GEN_6445;
        end else begin
          reservedFreeList2_8 <= _GEN_8566;
        end
      end else begin
        reservedFreeList2_8 <= _GEN_6445;
      end
    end else begin
      reservedFreeList2_8 <= _GEN_6445;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_9 <= _GEN_13600;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_9 <= _GEN_6446;
        end else begin
          reservedFreeList2_9 <= _GEN_8567;
        end
      end else begin
        reservedFreeList2_9 <= _GEN_6446;
      end
    end else begin
      reservedFreeList2_9 <= _GEN_6446;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_10 <= _GEN_13601;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_10 <= _GEN_6447;
        end else begin
          reservedFreeList2_10 <= _GEN_8568;
        end
      end else begin
        reservedFreeList2_10 <= _GEN_6447;
      end
    end else begin
      reservedFreeList2_10 <= _GEN_6447;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_11 <= _GEN_13602;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_11 <= _GEN_6448;
        end else begin
          reservedFreeList2_11 <= _GEN_8569;
        end
      end else begin
        reservedFreeList2_11 <= _GEN_6448;
      end
    end else begin
      reservedFreeList2_11 <= _GEN_6448;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_12 <= _GEN_13603;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_12 <= _GEN_6449;
        end else begin
          reservedFreeList2_12 <= _GEN_8570;
        end
      end else begin
        reservedFreeList2_12 <= _GEN_6449;
      end
    end else begin
      reservedFreeList2_12 <= _GEN_6449;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_13 <= _GEN_13604;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_13 <= _GEN_6450;
        end else begin
          reservedFreeList2_13 <= _GEN_8571;
        end
      end else begin
        reservedFreeList2_13 <= _GEN_6450;
      end
    end else begin
      reservedFreeList2_13 <= _GEN_6450;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_14 <= _GEN_13605;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_14 <= _GEN_6451;
        end else begin
          reservedFreeList2_14 <= _GEN_8572;
        end
      end else begin
        reservedFreeList2_14 <= _GEN_6451;
      end
    end else begin
      reservedFreeList2_14 <= _GEN_6451;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_15 <= _GEN_13606;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_15 <= _GEN_6452;
        end else begin
          reservedFreeList2_15 <= _GEN_8573;
        end
      end else begin
        reservedFreeList2_15 <= _GEN_6452;
      end
    end else begin
      reservedFreeList2_15 <= _GEN_6452;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_16 <= _GEN_13607;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_16 <= _GEN_6453;
        end else begin
          reservedFreeList2_16 <= _GEN_8574;
        end
      end else begin
        reservedFreeList2_16 <= _GEN_6453;
      end
    end else begin
      reservedFreeList2_16 <= _GEN_6453;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_17 <= _GEN_13608;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_17 <= _GEN_6454;
        end else begin
          reservedFreeList2_17 <= _GEN_8575;
        end
      end else begin
        reservedFreeList2_17 <= _GEN_6454;
      end
    end else begin
      reservedFreeList2_17 <= _GEN_6454;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_18 <= _GEN_13609;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_18 <= _GEN_6455;
        end else begin
          reservedFreeList2_18 <= _GEN_8576;
        end
      end else begin
        reservedFreeList2_18 <= _GEN_6455;
      end
    end else begin
      reservedFreeList2_18 <= _GEN_6455;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_19 <= _GEN_13610;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_19 <= _GEN_6456;
        end else begin
          reservedFreeList2_19 <= _GEN_8577;
        end
      end else begin
        reservedFreeList2_19 <= _GEN_6456;
      end
    end else begin
      reservedFreeList2_19 <= _GEN_6456;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_20 <= _GEN_13611;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_20 <= _GEN_6457;
        end else begin
          reservedFreeList2_20 <= _GEN_8578;
        end
      end else begin
        reservedFreeList2_20 <= _GEN_6457;
      end
    end else begin
      reservedFreeList2_20 <= _GEN_6457;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_21 <= _GEN_13612;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_21 <= _GEN_6458;
        end else begin
          reservedFreeList2_21 <= _GEN_8579;
        end
      end else begin
        reservedFreeList2_21 <= _GEN_6458;
      end
    end else begin
      reservedFreeList2_21 <= _GEN_6458;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_22 <= _GEN_13613;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_22 <= _GEN_6459;
        end else begin
          reservedFreeList2_22 <= _GEN_8580;
        end
      end else begin
        reservedFreeList2_22 <= _GEN_6459;
      end
    end else begin
      reservedFreeList2_22 <= _GEN_6459;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_23 <= _GEN_13614;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_23 <= _GEN_6460;
        end else begin
          reservedFreeList2_23 <= _GEN_8581;
        end
      end else begin
        reservedFreeList2_23 <= _GEN_6460;
      end
    end else begin
      reservedFreeList2_23 <= _GEN_6460;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_24 <= _GEN_13615;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_24 <= _GEN_6461;
        end else begin
          reservedFreeList2_24 <= _GEN_8582;
        end
      end else begin
        reservedFreeList2_24 <= _GEN_6461;
      end
    end else begin
      reservedFreeList2_24 <= _GEN_6461;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_25 <= _GEN_13616;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_25 <= _GEN_6462;
        end else begin
          reservedFreeList2_25 <= _GEN_8583;
        end
      end else begin
        reservedFreeList2_25 <= _GEN_6462;
      end
    end else begin
      reservedFreeList2_25 <= _GEN_6462;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_26 <= _GEN_13617;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_26 <= _GEN_6463;
        end else begin
          reservedFreeList2_26 <= _GEN_8584;
        end
      end else begin
        reservedFreeList2_26 <= _GEN_6463;
      end
    end else begin
      reservedFreeList2_26 <= _GEN_6463;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_27 <= _GEN_13618;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_27 <= _GEN_6464;
        end else begin
          reservedFreeList2_27 <= _GEN_8585;
        end
      end else begin
        reservedFreeList2_27 <= _GEN_6464;
      end
    end else begin
      reservedFreeList2_27 <= _GEN_6464;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_28 <= _GEN_13619;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_28 <= _GEN_6465;
        end else begin
          reservedFreeList2_28 <= _GEN_8586;
        end
      end else begin
        reservedFreeList2_28 <= _GEN_6465;
      end
    end else begin
      reservedFreeList2_28 <= _GEN_6465;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_29 <= _GEN_13620;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_29 <= _GEN_6466;
        end else begin
          reservedFreeList2_29 <= _GEN_8587;
        end
      end else begin
        reservedFreeList2_29 <= _GEN_6466;
      end
    end else begin
      reservedFreeList2_29 <= _GEN_6466;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_30 <= _GEN_13621;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_30 <= _GEN_6467;
        end else begin
          reservedFreeList2_30 <= _GEN_8588;
        end
      end else begin
        reservedFreeList2_30 <= _GEN_6467;
      end
    end else begin
      reservedFreeList2_30 <= _GEN_6467;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_31 <= _GEN_13622;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_31 <= _GEN_6468;
        end else begin
          reservedFreeList2_31 <= _GEN_8589;
        end
      end else begin
        reservedFreeList2_31 <= _GEN_6468;
      end
    end else begin
      reservedFreeList2_31 <= _GEN_6468;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_32 <= _GEN_13623;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_32 <= _GEN_6469;
        end else begin
          reservedFreeList2_32 <= _GEN_8590;
        end
      end else begin
        reservedFreeList2_32 <= _GEN_6469;
      end
    end else begin
      reservedFreeList2_32 <= _GEN_6469;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_33 <= _GEN_13624;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_33 <= _GEN_6470;
        end else begin
          reservedFreeList2_33 <= _GEN_8591;
        end
      end else begin
        reservedFreeList2_33 <= _GEN_6470;
      end
    end else begin
      reservedFreeList2_33 <= _GEN_6470;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_34 <= _GEN_13625;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_34 <= _GEN_6471;
        end else begin
          reservedFreeList2_34 <= _GEN_8592;
        end
      end else begin
        reservedFreeList2_34 <= _GEN_6471;
      end
    end else begin
      reservedFreeList2_34 <= _GEN_6471;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_35 <= _GEN_13626;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_35 <= _GEN_6472;
        end else begin
          reservedFreeList2_35 <= _GEN_8593;
        end
      end else begin
        reservedFreeList2_35 <= _GEN_6472;
      end
    end else begin
      reservedFreeList2_35 <= _GEN_6472;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_36 <= _GEN_13627;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_36 <= _GEN_6473;
        end else begin
          reservedFreeList2_36 <= _GEN_8594;
        end
      end else begin
        reservedFreeList2_36 <= _GEN_6473;
      end
    end else begin
      reservedFreeList2_36 <= _GEN_6473;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_37 <= _GEN_13628;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_37 <= _GEN_6474;
        end else begin
          reservedFreeList2_37 <= _GEN_8595;
        end
      end else begin
        reservedFreeList2_37 <= _GEN_6474;
      end
    end else begin
      reservedFreeList2_37 <= _GEN_6474;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_38 <= _GEN_13629;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_38 <= _GEN_6475;
        end else begin
          reservedFreeList2_38 <= _GEN_8596;
        end
      end else begin
        reservedFreeList2_38 <= _GEN_6475;
      end
    end else begin
      reservedFreeList2_38 <= _GEN_6475;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_39 <= _GEN_13630;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_39 <= _GEN_6476;
        end else begin
          reservedFreeList2_39 <= _GEN_8597;
        end
      end else begin
        reservedFreeList2_39 <= _GEN_6476;
      end
    end else begin
      reservedFreeList2_39 <= _GEN_6476;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_40 <= _GEN_13631;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_40 <= _GEN_6477;
        end else begin
          reservedFreeList2_40 <= _GEN_8598;
        end
      end else begin
        reservedFreeList2_40 <= _GEN_6477;
      end
    end else begin
      reservedFreeList2_40 <= _GEN_6477;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_41 <= _GEN_13632;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_41 <= _GEN_6478;
        end else begin
          reservedFreeList2_41 <= _GEN_8599;
        end
      end else begin
        reservedFreeList2_41 <= _GEN_6478;
      end
    end else begin
      reservedFreeList2_41 <= _GEN_6478;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_42 <= _GEN_13633;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_42 <= _GEN_6479;
        end else begin
          reservedFreeList2_42 <= _GEN_8600;
        end
      end else begin
        reservedFreeList2_42 <= _GEN_6479;
      end
    end else begin
      reservedFreeList2_42 <= _GEN_6479;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_43 <= _GEN_13634;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_43 <= _GEN_6480;
        end else begin
          reservedFreeList2_43 <= _GEN_8601;
        end
      end else begin
        reservedFreeList2_43 <= _GEN_6480;
      end
    end else begin
      reservedFreeList2_43 <= _GEN_6480;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_44 <= _GEN_13635;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_44 <= _GEN_6481;
        end else begin
          reservedFreeList2_44 <= _GEN_8602;
        end
      end else begin
        reservedFreeList2_44 <= _GEN_6481;
      end
    end else begin
      reservedFreeList2_44 <= _GEN_6481;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_45 <= _GEN_13636;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_45 <= _GEN_6482;
        end else begin
          reservedFreeList2_45 <= _GEN_8603;
        end
      end else begin
        reservedFreeList2_45 <= _GEN_6482;
      end
    end else begin
      reservedFreeList2_45 <= _GEN_6482;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_46 <= _GEN_13637;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_46 <= _GEN_6483;
        end else begin
          reservedFreeList2_46 <= _GEN_8604;
        end
      end else begin
        reservedFreeList2_46 <= _GEN_6483;
      end
    end else begin
      reservedFreeList2_46 <= _GEN_6483;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_47 <= _GEN_13638;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_47 <= _GEN_6484;
        end else begin
          reservedFreeList2_47 <= _GEN_8605;
        end
      end else begin
        reservedFreeList2_47 <= _GEN_6484;
      end
    end else begin
      reservedFreeList2_47 <= _GEN_6484;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_48 <= _GEN_13639;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_48 <= _GEN_6485;
        end else begin
          reservedFreeList2_48 <= _GEN_8606;
        end
      end else begin
        reservedFreeList2_48 <= _GEN_6485;
      end
    end else begin
      reservedFreeList2_48 <= _GEN_6485;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_49 <= _GEN_13640;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_49 <= _GEN_6486;
        end else begin
          reservedFreeList2_49 <= _GEN_8607;
        end
      end else begin
        reservedFreeList2_49 <= _GEN_6486;
      end
    end else begin
      reservedFreeList2_49 <= _GEN_6486;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_50 <= _GEN_13641;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_50 <= _GEN_6487;
        end else begin
          reservedFreeList2_50 <= _GEN_8608;
        end
      end else begin
        reservedFreeList2_50 <= _GEN_6487;
      end
    end else begin
      reservedFreeList2_50 <= _GEN_6487;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_51 <= _GEN_13642;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_51 <= _GEN_6488;
        end else begin
          reservedFreeList2_51 <= _GEN_8609;
        end
      end else begin
        reservedFreeList2_51 <= _GEN_6488;
      end
    end else begin
      reservedFreeList2_51 <= _GEN_6488;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_52 <= _GEN_13643;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_52 <= _GEN_6489;
        end else begin
          reservedFreeList2_52 <= _GEN_8610;
        end
      end else begin
        reservedFreeList2_52 <= _GEN_6489;
      end
    end else begin
      reservedFreeList2_52 <= _GEN_6489;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_53 <= _GEN_13644;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_53 <= _GEN_6490;
        end else begin
          reservedFreeList2_53 <= _GEN_8611;
        end
      end else begin
        reservedFreeList2_53 <= _GEN_6490;
      end
    end else begin
      reservedFreeList2_53 <= _GEN_6490;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_54 <= _GEN_13645;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_54 <= _GEN_6491;
        end else begin
          reservedFreeList2_54 <= _GEN_8612;
        end
      end else begin
        reservedFreeList2_54 <= _GEN_6491;
      end
    end else begin
      reservedFreeList2_54 <= _GEN_6491;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_55 <= _GEN_13646;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_55 <= _GEN_6492;
        end else begin
          reservedFreeList2_55 <= _GEN_8613;
        end
      end else begin
        reservedFreeList2_55 <= _GEN_6492;
      end
    end else begin
      reservedFreeList2_55 <= _GEN_6492;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_56 <= _GEN_13647;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_56 <= _GEN_6493;
        end else begin
          reservedFreeList2_56 <= _GEN_8614;
        end
      end else begin
        reservedFreeList2_56 <= _GEN_6493;
      end
    end else begin
      reservedFreeList2_56 <= _GEN_6493;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_57 <= _GEN_13648;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_57 <= _GEN_6494;
        end else begin
          reservedFreeList2_57 <= _GEN_8615;
        end
      end else begin
        reservedFreeList2_57 <= _GEN_6494;
      end
    end else begin
      reservedFreeList2_57 <= _GEN_6494;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_58 <= _GEN_13649;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_58 <= _GEN_6495;
        end else begin
          reservedFreeList2_58 <= _GEN_8616;
        end
      end else begin
        reservedFreeList2_58 <= _GEN_6495;
      end
    end else begin
      reservedFreeList2_58 <= _GEN_6495;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_59 <= _GEN_13650;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_59 <= _GEN_6496;
        end else begin
          reservedFreeList2_59 <= _GEN_8617;
        end
      end else begin
        reservedFreeList2_59 <= _GEN_6496;
      end
    end else begin
      reservedFreeList2_59 <= _GEN_6496;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_60 <= _GEN_13651;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_60 <= _GEN_6497;
        end else begin
          reservedFreeList2_60 <= _GEN_8618;
        end
      end else begin
        reservedFreeList2_60 <= _GEN_6497;
      end
    end else begin
      reservedFreeList2_60 <= _GEN_6497;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_61 <= _GEN_13652;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_61 <= _GEN_6498;
        end else begin
          reservedFreeList2_61 <= _GEN_8619;
        end
      end else begin
        reservedFreeList2_61 <= _GEN_6498;
      end
    end else begin
      reservedFreeList2_61 <= _GEN_6498;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList2_62 <= _GEN_13653;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList2_62 <= _GEN_6499;
        end else begin
          reservedFreeList2_62 <= _GEN_8620;
        end
      end else begin
        reservedFreeList2_62 <= _GEN_6499;
      end
    end else begin
      reservedFreeList2_62 <= _GEN_6499;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_0 <= _GEN_13655;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_0 <= _GEN_6501;
        end else begin
          reservedFreeList3_0 <= _GEN_8718;
        end
      end else begin
        reservedFreeList3_0 <= _GEN_6501;
      end
    end else begin
      reservedFreeList3_0 <= _GEN_6501;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_1 <= _GEN_13656;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_1 <= _GEN_6502;
        end else begin
          reservedFreeList3_1 <= _GEN_8719;
        end
      end else begin
        reservedFreeList3_1 <= _GEN_6502;
      end
    end else begin
      reservedFreeList3_1 <= _GEN_6502;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_2 <= _GEN_13657;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_2 <= _GEN_6503;
        end else begin
          reservedFreeList3_2 <= _GEN_8720;
        end
      end else begin
        reservedFreeList3_2 <= _GEN_6503;
      end
    end else begin
      reservedFreeList3_2 <= _GEN_6503;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_3 <= _GEN_13658;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_3 <= _GEN_6504;
        end else begin
          reservedFreeList3_3 <= _GEN_8721;
        end
      end else begin
        reservedFreeList3_3 <= _GEN_6504;
      end
    end else begin
      reservedFreeList3_3 <= _GEN_6504;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_4 <= _GEN_13659;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_4 <= _GEN_6505;
        end else begin
          reservedFreeList3_4 <= _GEN_8722;
        end
      end else begin
        reservedFreeList3_4 <= _GEN_6505;
      end
    end else begin
      reservedFreeList3_4 <= _GEN_6505;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_5 <= _GEN_13660;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_5 <= _GEN_6506;
        end else begin
          reservedFreeList3_5 <= _GEN_8723;
        end
      end else begin
        reservedFreeList3_5 <= _GEN_6506;
      end
    end else begin
      reservedFreeList3_5 <= _GEN_6506;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_6 <= _GEN_13661;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_6 <= _GEN_6507;
        end else begin
          reservedFreeList3_6 <= _GEN_8724;
        end
      end else begin
        reservedFreeList3_6 <= _GEN_6507;
      end
    end else begin
      reservedFreeList3_6 <= _GEN_6507;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_7 <= _GEN_13662;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_7 <= _GEN_6508;
        end else begin
          reservedFreeList3_7 <= _GEN_8725;
        end
      end else begin
        reservedFreeList3_7 <= _GEN_6508;
      end
    end else begin
      reservedFreeList3_7 <= _GEN_6508;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_8 <= _GEN_13663;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_8 <= _GEN_6509;
        end else begin
          reservedFreeList3_8 <= _GEN_8726;
        end
      end else begin
        reservedFreeList3_8 <= _GEN_6509;
      end
    end else begin
      reservedFreeList3_8 <= _GEN_6509;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_9 <= _GEN_13664;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_9 <= _GEN_6510;
        end else begin
          reservedFreeList3_9 <= _GEN_8727;
        end
      end else begin
        reservedFreeList3_9 <= _GEN_6510;
      end
    end else begin
      reservedFreeList3_9 <= _GEN_6510;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_10 <= _GEN_13665;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_10 <= _GEN_6511;
        end else begin
          reservedFreeList3_10 <= _GEN_8728;
        end
      end else begin
        reservedFreeList3_10 <= _GEN_6511;
      end
    end else begin
      reservedFreeList3_10 <= _GEN_6511;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_11 <= _GEN_13666;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_11 <= _GEN_6512;
        end else begin
          reservedFreeList3_11 <= _GEN_8729;
        end
      end else begin
        reservedFreeList3_11 <= _GEN_6512;
      end
    end else begin
      reservedFreeList3_11 <= _GEN_6512;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_12 <= _GEN_13667;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_12 <= _GEN_6513;
        end else begin
          reservedFreeList3_12 <= _GEN_8730;
        end
      end else begin
        reservedFreeList3_12 <= _GEN_6513;
      end
    end else begin
      reservedFreeList3_12 <= _GEN_6513;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_13 <= _GEN_13668;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_13 <= _GEN_6514;
        end else begin
          reservedFreeList3_13 <= _GEN_8731;
        end
      end else begin
        reservedFreeList3_13 <= _GEN_6514;
      end
    end else begin
      reservedFreeList3_13 <= _GEN_6514;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_14 <= _GEN_13669;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_14 <= _GEN_6515;
        end else begin
          reservedFreeList3_14 <= _GEN_8732;
        end
      end else begin
        reservedFreeList3_14 <= _GEN_6515;
      end
    end else begin
      reservedFreeList3_14 <= _GEN_6515;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_15 <= _GEN_13670;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_15 <= _GEN_6516;
        end else begin
          reservedFreeList3_15 <= _GEN_8733;
        end
      end else begin
        reservedFreeList3_15 <= _GEN_6516;
      end
    end else begin
      reservedFreeList3_15 <= _GEN_6516;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_16 <= _GEN_13671;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_16 <= _GEN_6517;
        end else begin
          reservedFreeList3_16 <= _GEN_8734;
        end
      end else begin
        reservedFreeList3_16 <= _GEN_6517;
      end
    end else begin
      reservedFreeList3_16 <= _GEN_6517;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_17 <= _GEN_13672;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_17 <= _GEN_6518;
        end else begin
          reservedFreeList3_17 <= _GEN_8735;
        end
      end else begin
        reservedFreeList3_17 <= _GEN_6518;
      end
    end else begin
      reservedFreeList3_17 <= _GEN_6518;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_18 <= _GEN_13673;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_18 <= _GEN_6519;
        end else begin
          reservedFreeList3_18 <= _GEN_8736;
        end
      end else begin
        reservedFreeList3_18 <= _GEN_6519;
      end
    end else begin
      reservedFreeList3_18 <= _GEN_6519;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_19 <= _GEN_13674;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_19 <= _GEN_6520;
        end else begin
          reservedFreeList3_19 <= _GEN_8737;
        end
      end else begin
        reservedFreeList3_19 <= _GEN_6520;
      end
    end else begin
      reservedFreeList3_19 <= _GEN_6520;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_20 <= _GEN_13675;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_20 <= _GEN_6521;
        end else begin
          reservedFreeList3_20 <= _GEN_8738;
        end
      end else begin
        reservedFreeList3_20 <= _GEN_6521;
      end
    end else begin
      reservedFreeList3_20 <= _GEN_6521;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_21 <= _GEN_13676;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_21 <= _GEN_6522;
        end else begin
          reservedFreeList3_21 <= _GEN_8739;
        end
      end else begin
        reservedFreeList3_21 <= _GEN_6522;
      end
    end else begin
      reservedFreeList3_21 <= _GEN_6522;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_22 <= _GEN_13677;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_22 <= _GEN_6523;
        end else begin
          reservedFreeList3_22 <= _GEN_8740;
        end
      end else begin
        reservedFreeList3_22 <= _GEN_6523;
      end
    end else begin
      reservedFreeList3_22 <= _GEN_6523;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_23 <= _GEN_13678;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_23 <= _GEN_6524;
        end else begin
          reservedFreeList3_23 <= _GEN_8741;
        end
      end else begin
        reservedFreeList3_23 <= _GEN_6524;
      end
    end else begin
      reservedFreeList3_23 <= _GEN_6524;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_24 <= _GEN_13679;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_24 <= _GEN_6525;
        end else begin
          reservedFreeList3_24 <= _GEN_8742;
        end
      end else begin
        reservedFreeList3_24 <= _GEN_6525;
      end
    end else begin
      reservedFreeList3_24 <= _GEN_6525;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_25 <= _GEN_13680;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_25 <= _GEN_6526;
        end else begin
          reservedFreeList3_25 <= _GEN_8743;
        end
      end else begin
        reservedFreeList3_25 <= _GEN_6526;
      end
    end else begin
      reservedFreeList3_25 <= _GEN_6526;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_26 <= _GEN_13681;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_26 <= _GEN_6527;
        end else begin
          reservedFreeList3_26 <= _GEN_8744;
        end
      end else begin
        reservedFreeList3_26 <= _GEN_6527;
      end
    end else begin
      reservedFreeList3_26 <= _GEN_6527;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_27 <= _GEN_13682;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_27 <= _GEN_6528;
        end else begin
          reservedFreeList3_27 <= _GEN_8745;
        end
      end else begin
        reservedFreeList3_27 <= _GEN_6528;
      end
    end else begin
      reservedFreeList3_27 <= _GEN_6528;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_28 <= _GEN_13683;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_28 <= _GEN_6529;
        end else begin
          reservedFreeList3_28 <= _GEN_8746;
        end
      end else begin
        reservedFreeList3_28 <= _GEN_6529;
      end
    end else begin
      reservedFreeList3_28 <= _GEN_6529;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_29 <= _GEN_13684;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_29 <= _GEN_6530;
        end else begin
          reservedFreeList3_29 <= _GEN_8747;
        end
      end else begin
        reservedFreeList3_29 <= _GEN_6530;
      end
    end else begin
      reservedFreeList3_29 <= _GEN_6530;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_30 <= _GEN_13685;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_30 <= _GEN_6531;
        end else begin
          reservedFreeList3_30 <= _GEN_8748;
        end
      end else begin
        reservedFreeList3_30 <= _GEN_6531;
      end
    end else begin
      reservedFreeList3_30 <= _GEN_6531;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_31 <= _GEN_13686;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_31 <= _GEN_6532;
        end else begin
          reservedFreeList3_31 <= _GEN_8749;
        end
      end else begin
        reservedFreeList3_31 <= _GEN_6532;
      end
    end else begin
      reservedFreeList3_31 <= _GEN_6532;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_32 <= _GEN_13687;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_32 <= _GEN_6533;
        end else begin
          reservedFreeList3_32 <= _GEN_8750;
        end
      end else begin
        reservedFreeList3_32 <= _GEN_6533;
      end
    end else begin
      reservedFreeList3_32 <= _GEN_6533;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_33 <= _GEN_13688;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_33 <= _GEN_6534;
        end else begin
          reservedFreeList3_33 <= _GEN_8751;
        end
      end else begin
        reservedFreeList3_33 <= _GEN_6534;
      end
    end else begin
      reservedFreeList3_33 <= _GEN_6534;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_34 <= _GEN_13689;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_34 <= _GEN_6535;
        end else begin
          reservedFreeList3_34 <= _GEN_8752;
        end
      end else begin
        reservedFreeList3_34 <= _GEN_6535;
      end
    end else begin
      reservedFreeList3_34 <= _GEN_6535;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_35 <= _GEN_13690;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_35 <= _GEN_6536;
        end else begin
          reservedFreeList3_35 <= _GEN_8753;
        end
      end else begin
        reservedFreeList3_35 <= _GEN_6536;
      end
    end else begin
      reservedFreeList3_35 <= _GEN_6536;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_36 <= _GEN_13691;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_36 <= _GEN_6537;
        end else begin
          reservedFreeList3_36 <= _GEN_8754;
        end
      end else begin
        reservedFreeList3_36 <= _GEN_6537;
      end
    end else begin
      reservedFreeList3_36 <= _GEN_6537;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_37 <= _GEN_13692;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_37 <= _GEN_6538;
        end else begin
          reservedFreeList3_37 <= _GEN_8755;
        end
      end else begin
        reservedFreeList3_37 <= _GEN_6538;
      end
    end else begin
      reservedFreeList3_37 <= _GEN_6538;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_38 <= _GEN_13693;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_38 <= _GEN_6539;
        end else begin
          reservedFreeList3_38 <= _GEN_8756;
        end
      end else begin
        reservedFreeList3_38 <= _GEN_6539;
      end
    end else begin
      reservedFreeList3_38 <= _GEN_6539;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_39 <= _GEN_13694;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_39 <= _GEN_6540;
        end else begin
          reservedFreeList3_39 <= _GEN_8757;
        end
      end else begin
        reservedFreeList3_39 <= _GEN_6540;
      end
    end else begin
      reservedFreeList3_39 <= _GEN_6540;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_40 <= _GEN_13695;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_40 <= _GEN_6541;
        end else begin
          reservedFreeList3_40 <= _GEN_8758;
        end
      end else begin
        reservedFreeList3_40 <= _GEN_6541;
      end
    end else begin
      reservedFreeList3_40 <= _GEN_6541;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_41 <= _GEN_13696;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_41 <= _GEN_6542;
        end else begin
          reservedFreeList3_41 <= _GEN_8759;
        end
      end else begin
        reservedFreeList3_41 <= _GEN_6542;
      end
    end else begin
      reservedFreeList3_41 <= _GEN_6542;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_42 <= _GEN_13697;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_42 <= _GEN_6543;
        end else begin
          reservedFreeList3_42 <= _GEN_8760;
        end
      end else begin
        reservedFreeList3_42 <= _GEN_6543;
      end
    end else begin
      reservedFreeList3_42 <= _GEN_6543;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_43 <= _GEN_13698;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_43 <= _GEN_6544;
        end else begin
          reservedFreeList3_43 <= _GEN_8761;
        end
      end else begin
        reservedFreeList3_43 <= _GEN_6544;
      end
    end else begin
      reservedFreeList3_43 <= _GEN_6544;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_44 <= _GEN_13699;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_44 <= _GEN_6545;
        end else begin
          reservedFreeList3_44 <= _GEN_8762;
        end
      end else begin
        reservedFreeList3_44 <= _GEN_6545;
      end
    end else begin
      reservedFreeList3_44 <= _GEN_6545;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_45 <= _GEN_13700;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_45 <= _GEN_6546;
        end else begin
          reservedFreeList3_45 <= _GEN_8763;
        end
      end else begin
        reservedFreeList3_45 <= _GEN_6546;
      end
    end else begin
      reservedFreeList3_45 <= _GEN_6546;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_46 <= _GEN_13701;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_46 <= _GEN_6547;
        end else begin
          reservedFreeList3_46 <= _GEN_8764;
        end
      end else begin
        reservedFreeList3_46 <= _GEN_6547;
      end
    end else begin
      reservedFreeList3_46 <= _GEN_6547;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_47 <= _GEN_13702;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_47 <= _GEN_6548;
        end else begin
          reservedFreeList3_47 <= _GEN_8765;
        end
      end else begin
        reservedFreeList3_47 <= _GEN_6548;
      end
    end else begin
      reservedFreeList3_47 <= _GEN_6548;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_48 <= _GEN_13703;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_48 <= _GEN_6549;
        end else begin
          reservedFreeList3_48 <= _GEN_8766;
        end
      end else begin
        reservedFreeList3_48 <= _GEN_6549;
      end
    end else begin
      reservedFreeList3_48 <= _GEN_6549;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_49 <= _GEN_13704;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_49 <= _GEN_6550;
        end else begin
          reservedFreeList3_49 <= _GEN_8767;
        end
      end else begin
        reservedFreeList3_49 <= _GEN_6550;
      end
    end else begin
      reservedFreeList3_49 <= _GEN_6550;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_50 <= _GEN_13705;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_50 <= _GEN_6551;
        end else begin
          reservedFreeList3_50 <= _GEN_8768;
        end
      end else begin
        reservedFreeList3_50 <= _GEN_6551;
      end
    end else begin
      reservedFreeList3_50 <= _GEN_6551;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_51 <= _GEN_13706;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_51 <= _GEN_6552;
        end else begin
          reservedFreeList3_51 <= _GEN_8769;
        end
      end else begin
        reservedFreeList3_51 <= _GEN_6552;
      end
    end else begin
      reservedFreeList3_51 <= _GEN_6552;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_52 <= _GEN_13707;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_52 <= _GEN_6553;
        end else begin
          reservedFreeList3_52 <= _GEN_8770;
        end
      end else begin
        reservedFreeList3_52 <= _GEN_6553;
      end
    end else begin
      reservedFreeList3_52 <= _GEN_6553;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_53 <= _GEN_13708;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_53 <= _GEN_6554;
        end else begin
          reservedFreeList3_53 <= _GEN_8771;
        end
      end else begin
        reservedFreeList3_53 <= _GEN_6554;
      end
    end else begin
      reservedFreeList3_53 <= _GEN_6554;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_54 <= _GEN_13709;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_54 <= _GEN_6555;
        end else begin
          reservedFreeList3_54 <= _GEN_8772;
        end
      end else begin
        reservedFreeList3_54 <= _GEN_6555;
      end
    end else begin
      reservedFreeList3_54 <= _GEN_6555;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_55 <= _GEN_13710;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_55 <= _GEN_6556;
        end else begin
          reservedFreeList3_55 <= _GEN_8773;
        end
      end else begin
        reservedFreeList3_55 <= _GEN_6556;
      end
    end else begin
      reservedFreeList3_55 <= _GEN_6556;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_56 <= _GEN_13711;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_56 <= _GEN_6557;
        end else begin
          reservedFreeList3_56 <= _GEN_8774;
        end
      end else begin
        reservedFreeList3_56 <= _GEN_6557;
      end
    end else begin
      reservedFreeList3_56 <= _GEN_6557;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_57 <= _GEN_13712;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_57 <= _GEN_6558;
        end else begin
          reservedFreeList3_57 <= _GEN_8775;
        end
      end else begin
        reservedFreeList3_57 <= _GEN_6558;
      end
    end else begin
      reservedFreeList3_57 <= _GEN_6558;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_58 <= _GEN_13713;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_58 <= _GEN_6559;
        end else begin
          reservedFreeList3_58 <= _GEN_8776;
        end
      end else begin
        reservedFreeList3_58 <= _GEN_6559;
      end
    end else begin
      reservedFreeList3_58 <= _GEN_6559;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_59 <= _GEN_13714;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_59 <= _GEN_6560;
        end else begin
          reservedFreeList3_59 <= _GEN_8777;
        end
      end else begin
        reservedFreeList3_59 <= _GEN_6560;
      end
    end else begin
      reservedFreeList3_59 <= _GEN_6560;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_60 <= _GEN_13715;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_60 <= _GEN_6561;
        end else begin
          reservedFreeList3_60 <= _GEN_8778;
        end
      end else begin
        reservedFreeList3_60 <= _GEN_6561;
      end
    end else begin
      reservedFreeList3_60 <= _GEN_6561;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_61 <= _GEN_13716;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_61 <= _GEN_6562;
        end else begin
          reservedFreeList3_61 <= _GEN_8779;
        end
      end else begin
        reservedFreeList3_61 <= _GEN_6562;
      end
    end else begin
      reservedFreeList3_61 <= _GEN_6562;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList3_62 <= _GEN_13717;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedFreeList3_62 <= _GEN_6563;
        end else begin
          reservedFreeList3_62 <= _GEN_8780;
        end
      end else begin
        reservedFreeList3_62 <= _GEN_6563;
      end
    end else begin
      reservedFreeList3_62 <= _GEN_6563;
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_0 <= _GEN_13719;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_0 <= _GEN_8878;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_1 <= _GEN_13720;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_1 <= _GEN_8879;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_2 <= _GEN_13721;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_2 <= _GEN_8880;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_3 <= _GEN_13722;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_3 <= _GEN_8881;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_4 <= _GEN_13723;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_4 <= _GEN_8882;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_5 <= _GEN_13724;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_5 <= _GEN_8883;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_6 <= _GEN_13725;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_6 <= _GEN_8884;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_7 <= _GEN_13726;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_7 <= _GEN_8885;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_8 <= _GEN_13727;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_8 <= _GEN_8886;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_9 <= _GEN_13728;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_9 <= _GEN_8887;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_10 <= _GEN_13729;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_10 <= _GEN_8888;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_11 <= _GEN_13730;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_11 <= _GEN_8889;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_12 <= _GEN_13731;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_12 <= _GEN_8890;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_13 <= _GEN_13732;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_13 <= _GEN_8891;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_14 <= _GEN_13733;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_14 <= _GEN_8892;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_15 <= _GEN_13734;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_15 <= _GEN_8893;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_16 <= _GEN_13735;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_16 <= _GEN_8894;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_17 <= _GEN_13736;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_17 <= _GEN_8895;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_18 <= _GEN_13737;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_18 <= _GEN_8896;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_19 <= _GEN_13738;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_19 <= _GEN_8897;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_20 <= _GEN_13739;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_20 <= _GEN_8898;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_21 <= _GEN_13740;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_21 <= _GEN_8899;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_22 <= _GEN_13741;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_22 <= _GEN_8900;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_23 <= _GEN_13742;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_23 <= _GEN_8901;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_24 <= _GEN_13743;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_24 <= _GEN_8902;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_25 <= _GEN_13744;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_25 <= _GEN_8903;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_26 <= _GEN_13745;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_26 <= _GEN_8904;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_27 <= _GEN_13746;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_27 <= _GEN_8905;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_28 <= _GEN_13747;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_28 <= _GEN_8906;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_29 <= _GEN_13748;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_29 <= _GEN_8907;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_30 <= _GEN_13749;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_30 <= _GEN_8908;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_31 <= _GEN_13750;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_31 <= _GEN_8909;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_32 <= _GEN_13751;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_32 <= _GEN_8910;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_33 <= _GEN_13752;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_33 <= _GEN_8911;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_34 <= _GEN_13753;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_34 <= _GEN_8912;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_35 <= _GEN_13754;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_35 <= _GEN_8913;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_36 <= _GEN_13755;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_36 <= _GEN_8914;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_37 <= _GEN_13756;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_37 <= _GEN_8915;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_38 <= _GEN_13757;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_38 <= _GEN_8916;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_39 <= _GEN_13758;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_39 <= _GEN_8917;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_40 <= _GEN_13759;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_40 <= _GEN_8918;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_41 <= _GEN_13760;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_41 <= _GEN_8919;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_42 <= _GEN_13761;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_42 <= _GEN_8920;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_43 <= _GEN_13762;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_43 <= _GEN_8921;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_44 <= _GEN_13763;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_44 <= _GEN_8922;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_45 <= _GEN_13764;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_45 <= _GEN_8923;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_46 <= _GEN_13765;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_46 <= _GEN_8924;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_47 <= _GEN_13766;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_47 <= _GEN_8925;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_48 <= _GEN_13767;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_48 <= _GEN_8926;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_49 <= _GEN_13768;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_49 <= _GEN_8927;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_50 <= _GEN_13769;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_50 <= _GEN_8928;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_51 <= _GEN_13770;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_51 <= _GEN_8929;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_52 <= _GEN_13771;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_52 <= _GEN_8930;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_53 <= _GEN_13772;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_53 <= _GEN_8931;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_54 <= _GEN_13773;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_54 <= _GEN_8932;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_55 <= _GEN_13774;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_55 <= _GEN_8933;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_56 <= _GEN_13775;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_56 <= _GEN_8934;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_57 <= _GEN_13776;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_57 <= _GEN_8935;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_58 <= _GEN_13777;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_58 <= _GEN_8936;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_59 <= _GEN_13778;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_59 <= _GEN_8937;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_60 <= _GEN_13779;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_60 <= _GEN_8938;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_61 <= _GEN_13780;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_61 <= _GEN_8939;
        end
      end
    end
    if (_T_474) begin // @[decode.scala 889:5]
      reservedFreeList4_62 <= _GEN_13781;
    end else if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          reservedFreeList4_62 <= _GEN_8940;
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_0 <= _GEN_6862;
          end else begin
            reservedValidList1_0 <= PRFValidList_0; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_0 <= _GEN_6565;
        end
      end else begin
        reservedValidList1_0 <= _GEN_6565;
      end
    end else begin
      reservedValidList1_0 <= _GEN_6565;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_1 <= _GEN_6863;
          end else begin
            reservedValidList1_1 <= PRFValidList_1; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_1 <= _GEN_6566;
        end
      end else begin
        reservedValidList1_1 <= _GEN_6566;
      end
    end else begin
      reservedValidList1_1 <= _GEN_6566;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_2 <= _GEN_6864;
          end else begin
            reservedValidList1_2 <= PRFValidList_2; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_2 <= _GEN_6567;
        end
      end else begin
        reservedValidList1_2 <= _GEN_6567;
      end
    end else begin
      reservedValidList1_2 <= _GEN_6567;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_3 <= _GEN_6865;
          end else begin
            reservedValidList1_3 <= PRFValidList_3; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_3 <= _GEN_6568;
        end
      end else begin
        reservedValidList1_3 <= _GEN_6568;
      end
    end else begin
      reservedValidList1_3 <= _GEN_6568;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_4 <= _GEN_6866;
          end else begin
            reservedValidList1_4 <= PRFValidList_4; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_4 <= _GEN_6569;
        end
      end else begin
        reservedValidList1_4 <= _GEN_6569;
      end
    end else begin
      reservedValidList1_4 <= _GEN_6569;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_5 <= _GEN_6867;
          end else begin
            reservedValidList1_5 <= PRFValidList_5; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_5 <= _GEN_6570;
        end
      end else begin
        reservedValidList1_5 <= _GEN_6570;
      end
    end else begin
      reservedValidList1_5 <= _GEN_6570;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_6 <= _GEN_6868;
          end else begin
            reservedValidList1_6 <= PRFValidList_6; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_6 <= _GEN_6571;
        end
      end else begin
        reservedValidList1_6 <= _GEN_6571;
      end
    end else begin
      reservedValidList1_6 <= _GEN_6571;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_7 <= _GEN_6869;
          end else begin
            reservedValidList1_7 <= PRFValidList_7; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_7 <= _GEN_6572;
        end
      end else begin
        reservedValidList1_7 <= _GEN_6572;
      end
    end else begin
      reservedValidList1_7 <= _GEN_6572;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_8 <= _GEN_6870;
          end else begin
            reservedValidList1_8 <= PRFValidList_8; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_8 <= _GEN_6573;
        end
      end else begin
        reservedValidList1_8 <= _GEN_6573;
      end
    end else begin
      reservedValidList1_8 <= _GEN_6573;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_9 <= _GEN_6871;
          end else begin
            reservedValidList1_9 <= PRFValidList_9; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_9 <= _GEN_6574;
        end
      end else begin
        reservedValidList1_9 <= _GEN_6574;
      end
    end else begin
      reservedValidList1_9 <= _GEN_6574;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_10 <= _GEN_6872;
          end else begin
            reservedValidList1_10 <= PRFValidList_10; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_10 <= _GEN_6575;
        end
      end else begin
        reservedValidList1_10 <= _GEN_6575;
      end
    end else begin
      reservedValidList1_10 <= _GEN_6575;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_11 <= _GEN_6873;
          end else begin
            reservedValidList1_11 <= PRFValidList_11; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_11 <= _GEN_6576;
        end
      end else begin
        reservedValidList1_11 <= _GEN_6576;
      end
    end else begin
      reservedValidList1_11 <= _GEN_6576;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_12 <= _GEN_6874;
          end else begin
            reservedValidList1_12 <= PRFValidList_12; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_12 <= _GEN_6577;
        end
      end else begin
        reservedValidList1_12 <= _GEN_6577;
      end
    end else begin
      reservedValidList1_12 <= _GEN_6577;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_13 <= _GEN_6875;
          end else begin
            reservedValidList1_13 <= PRFValidList_13; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_13 <= _GEN_6578;
        end
      end else begin
        reservedValidList1_13 <= _GEN_6578;
      end
    end else begin
      reservedValidList1_13 <= _GEN_6578;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_14 <= _GEN_6876;
          end else begin
            reservedValidList1_14 <= PRFValidList_14; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_14 <= _GEN_6579;
        end
      end else begin
        reservedValidList1_14 <= _GEN_6579;
      end
    end else begin
      reservedValidList1_14 <= _GEN_6579;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_15 <= _GEN_6877;
          end else begin
            reservedValidList1_15 <= PRFValidList_15; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_15 <= _GEN_6580;
        end
      end else begin
        reservedValidList1_15 <= _GEN_6580;
      end
    end else begin
      reservedValidList1_15 <= _GEN_6580;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_16 <= _GEN_6878;
          end else begin
            reservedValidList1_16 <= PRFValidList_16; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_16 <= _GEN_6581;
        end
      end else begin
        reservedValidList1_16 <= _GEN_6581;
      end
    end else begin
      reservedValidList1_16 <= _GEN_6581;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_17 <= _GEN_6879;
          end else begin
            reservedValidList1_17 <= PRFValidList_17; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_17 <= _GEN_6582;
        end
      end else begin
        reservedValidList1_17 <= _GEN_6582;
      end
    end else begin
      reservedValidList1_17 <= _GEN_6582;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_18 <= _GEN_6880;
          end else begin
            reservedValidList1_18 <= PRFValidList_18; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_18 <= _GEN_6583;
        end
      end else begin
        reservedValidList1_18 <= _GEN_6583;
      end
    end else begin
      reservedValidList1_18 <= _GEN_6583;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_19 <= _GEN_6881;
          end else begin
            reservedValidList1_19 <= PRFValidList_19; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_19 <= _GEN_6584;
        end
      end else begin
        reservedValidList1_19 <= _GEN_6584;
      end
    end else begin
      reservedValidList1_19 <= _GEN_6584;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_20 <= _GEN_6882;
          end else begin
            reservedValidList1_20 <= PRFValidList_20; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_20 <= _GEN_6585;
        end
      end else begin
        reservedValidList1_20 <= _GEN_6585;
      end
    end else begin
      reservedValidList1_20 <= _GEN_6585;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_21 <= _GEN_6883;
          end else begin
            reservedValidList1_21 <= PRFValidList_21; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_21 <= _GEN_6586;
        end
      end else begin
        reservedValidList1_21 <= _GEN_6586;
      end
    end else begin
      reservedValidList1_21 <= _GEN_6586;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_22 <= _GEN_6884;
          end else begin
            reservedValidList1_22 <= PRFValidList_22; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_22 <= _GEN_6587;
        end
      end else begin
        reservedValidList1_22 <= _GEN_6587;
      end
    end else begin
      reservedValidList1_22 <= _GEN_6587;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_23 <= _GEN_6885;
          end else begin
            reservedValidList1_23 <= PRFValidList_23; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_23 <= _GEN_6588;
        end
      end else begin
        reservedValidList1_23 <= _GEN_6588;
      end
    end else begin
      reservedValidList1_23 <= _GEN_6588;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_24 <= _GEN_6886;
          end else begin
            reservedValidList1_24 <= PRFValidList_24; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_24 <= _GEN_6589;
        end
      end else begin
        reservedValidList1_24 <= _GEN_6589;
      end
    end else begin
      reservedValidList1_24 <= _GEN_6589;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_25 <= _GEN_6887;
          end else begin
            reservedValidList1_25 <= PRFValidList_25; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_25 <= _GEN_6590;
        end
      end else begin
        reservedValidList1_25 <= _GEN_6590;
      end
    end else begin
      reservedValidList1_25 <= _GEN_6590;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_26 <= _GEN_6888;
          end else begin
            reservedValidList1_26 <= PRFValidList_26; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_26 <= _GEN_6591;
        end
      end else begin
        reservedValidList1_26 <= _GEN_6591;
      end
    end else begin
      reservedValidList1_26 <= _GEN_6591;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_27 <= _GEN_6889;
          end else begin
            reservedValidList1_27 <= PRFValidList_27; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_27 <= _GEN_6592;
        end
      end else begin
        reservedValidList1_27 <= _GEN_6592;
      end
    end else begin
      reservedValidList1_27 <= _GEN_6592;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_28 <= _GEN_6890;
          end else begin
            reservedValidList1_28 <= PRFValidList_28; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_28 <= _GEN_6593;
        end
      end else begin
        reservedValidList1_28 <= _GEN_6593;
      end
    end else begin
      reservedValidList1_28 <= _GEN_6593;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_29 <= _GEN_6891;
          end else begin
            reservedValidList1_29 <= PRFValidList_29; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_29 <= _GEN_6594;
        end
      end else begin
        reservedValidList1_29 <= _GEN_6594;
      end
    end else begin
      reservedValidList1_29 <= _GEN_6594;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_30 <= _GEN_6892;
          end else begin
            reservedValidList1_30 <= PRFValidList_30; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_30 <= _GEN_6595;
        end
      end else begin
        reservedValidList1_30 <= _GEN_6595;
      end
    end else begin
      reservedValidList1_30 <= _GEN_6595;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_31 <= _GEN_6893;
          end else begin
            reservedValidList1_31 <= PRFValidList_31; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_31 <= _GEN_6596;
        end
      end else begin
        reservedValidList1_31 <= _GEN_6596;
      end
    end else begin
      reservedValidList1_31 <= _GEN_6596;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_32 <= _GEN_6894;
          end else begin
            reservedValidList1_32 <= PRFValidList_32; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_32 <= _GEN_6597;
        end
      end else begin
        reservedValidList1_32 <= _GEN_6597;
      end
    end else begin
      reservedValidList1_32 <= _GEN_6597;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_33 <= _GEN_6895;
          end else begin
            reservedValidList1_33 <= PRFValidList_33; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_33 <= _GEN_6598;
        end
      end else begin
        reservedValidList1_33 <= _GEN_6598;
      end
    end else begin
      reservedValidList1_33 <= _GEN_6598;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_34 <= _GEN_6896;
          end else begin
            reservedValidList1_34 <= PRFValidList_34; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_34 <= _GEN_6599;
        end
      end else begin
        reservedValidList1_34 <= _GEN_6599;
      end
    end else begin
      reservedValidList1_34 <= _GEN_6599;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_35 <= _GEN_6897;
          end else begin
            reservedValidList1_35 <= PRFValidList_35; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_35 <= _GEN_6600;
        end
      end else begin
        reservedValidList1_35 <= _GEN_6600;
      end
    end else begin
      reservedValidList1_35 <= _GEN_6600;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_36 <= _GEN_6898;
          end else begin
            reservedValidList1_36 <= PRFValidList_36; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_36 <= _GEN_6601;
        end
      end else begin
        reservedValidList1_36 <= _GEN_6601;
      end
    end else begin
      reservedValidList1_36 <= _GEN_6601;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_37 <= _GEN_6899;
          end else begin
            reservedValidList1_37 <= PRFValidList_37; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_37 <= _GEN_6602;
        end
      end else begin
        reservedValidList1_37 <= _GEN_6602;
      end
    end else begin
      reservedValidList1_37 <= _GEN_6602;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_38 <= _GEN_6900;
          end else begin
            reservedValidList1_38 <= PRFValidList_38; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_38 <= _GEN_6603;
        end
      end else begin
        reservedValidList1_38 <= _GEN_6603;
      end
    end else begin
      reservedValidList1_38 <= _GEN_6603;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_39 <= _GEN_6901;
          end else begin
            reservedValidList1_39 <= PRFValidList_39; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_39 <= _GEN_6604;
        end
      end else begin
        reservedValidList1_39 <= _GEN_6604;
      end
    end else begin
      reservedValidList1_39 <= _GEN_6604;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_40 <= _GEN_6902;
          end else begin
            reservedValidList1_40 <= PRFValidList_40; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_40 <= _GEN_6605;
        end
      end else begin
        reservedValidList1_40 <= _GEN_6605;
      end
    end else begin
      reservedValidList1_40 <= _GEN_6605;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_41 <= _GEN_6903;
          end else begin
            reservedValidList1_41 <= PRFValidList_41; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_41 <= _GEN_6606;
        end
      end else begin
        reservedValidList1_41 <= _GEN_6606;
      end
    end else begin
      reservedValidList1_41 <= _GEN_6606;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_42 <= _GEN_6904;
          end else begin
            reservedValidList1_42 <= PRFValidList_42; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_42 <= _GEN_6607;
        end
      end else begin
        reservedValidList1_42 <= _GEN_6607;
      end
    end else begin
      reservedValidList1_42 <= _GEN_6607;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_43 <= _GEN_6905;
          end else begin
            reservedValidList1_43 <= PRFValidList_43; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_43 <= _GEN_6608;
        end
      end else begin
        reservedValidList1_43 <= _GEN_6608;
      end
    end else begin
      reservedValidList1_43 <= _GEN_6608;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_44 <= _GEN_6906;
          end else begin
            reservedValidList1_44 <= PRFValidList_44; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_44 <= _GEN_6609;
        end
      end else begin
        reservedValidList1_44 <= _GEN_6609;
      end
    end else begin
      reservedValidList1_44 <= _GEN_6609;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_45 <= _GEN_6907;
          end else begin
            reservedValidList1_45 <= PRFValidList_45; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_45 <= _GEN_6610;
        end
      end else begin
        reservedValidList1_45 <= _GEN_6610;
      end
    end else begin
      reservedValidList1_45 <= _GEN_6610;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_46 <= _GEN_6908;
          end else begin
            reservedValidList1_46 <= PRFValidList_46; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_46 <= _GEN_6611;
        end
      end else begin
        reservedValidList1_46 <= _GEN_6611;
      end
    end else begin
      reservedValidList1_46 <= _GEN_6611;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_47 <= _GEN_6909;
          end else begin
            reservedValidList1_47 <= PRFValidList_47; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_47 <= _GEN_6612;
        end
      end else begin
        reservedValidList1_47 <= _GEN_6612;
      end
    end else begin
      reservedValidList1_47 <= _GEN_6612;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_48 <= _GEN_6910;
          end else begin
            reservedValidList1_48 <= PRFValidList_48; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_48 <= _GEN_6613;
        end
      end else begin
        reservedValidList1_48 <= _GEN_6613;
      end
    end else begin
      reservedValidList1_48 <= _GEN_6613;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_49 <= _GEN_6911;
          end else begin
            reservedValidList1_49 <= PRFValidList_49; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_49 <= _GEN_6614;
        end
      end else begin
        reservedValidList1_49 <= _GEN_6614;
      end
    end else begin
      reservedValidList1_49 <= _GEN_6614;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_50 <= _GEN_6912;
          end else begin
            reservedValidList1_50 <= PRFValidList_50; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_50 <= _GEN_6615;
        end
      end else begin
        reservedValidList1_50 <= _GEN_6615;
      end
    end else begin
      reservedValidList1_50 <= _GEN_6615;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_51 <= _GEN_6913;
          end else begin
            reservedValidList1_51 <= PRFValidList_51; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_51 <= _GEN_6616;
        end
      end else begin
        reservedValidList1_51 <= _GEN_6616;
      end
    end else begin
      reservedValidList1_51 <= _GEN_6616;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_52 <= _GEN_6914;
          end else begin
            reservedValidList1_52 <= PRFValidList_52; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_52 <= _GEN_6617;
        end
      end else begin
        reservedValidList1_52 <= _GEN_6617;
      end
    end else begin
      reservedValidList1_52 <= _GEN_6617;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_53 <= _GEN_6915;
          end else begin
            reservedValidList1_53 <= PRFValidList_53; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_53 <= _GEN_6618;
        end
      end else begin
        reservedValidList1_53 <= _GEN_6618;
      end
    end else begin
      reservedValidList1_53 <= _GEN_6618;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_54 <= _GEN_6916;
          end else begin
            reservedValidList1_54 <= PRFValidList_54; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_54 <= _GEN_6619;
        end
      end else begin
        reservedValidList1_54 <= _GEN_6619;
      end
    end else begin
      reservedValidList1_54 <= _GEN_6619;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_55 <= _GEN_6917;
          end else begin
            reservedValidList1_55 <= PRFValidList_55; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_55 <= _GEN_6620;
        end
      end else begin
        reservedValidList1_55 <= _GEN_6620;
      end
    end else begin
      reservedValidList1_55 <= _GEN_6620;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_56 <= _GEN_6918;
          end else begin
            reservedValidList1_56 <= PRFValidList_56; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_56 <= _GEN_6621;
        end
      end else begin
        reservedValidList1_56 <= _GEN_6621;
      end
    end else begin
      reservedValidList1_56 <= _GEN_6621;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_57 <= _GEN_6919;
          end else begin
            reservedValidList1_57 <= PRFValidList_57; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_57 <= _GEN_6622;
        end
      end else begin
        reservedValidList1_57 <= _GEN_6622;
      end
    end else begin
      reservedValidList1_57 <= _GEN_6622;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_58 <= _GEN_6920;
          end else begin
            reservedValidList1_58 <= PRFValidList_58; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_58 <= _GEN_6623;
        end
      end else begin
        reservedValidList1_58 <= _GEN_6623;
      end
    end else begin
      reservedValidList1_58 <= _GEN_6623;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_59 <= _GEN_6921;
          end else begin
            reservedValidList1_59 <= PRFValidList_59; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_59 <= _GEN_6624;
        end
      end else begin
        reservedValidList1_59 <= _GEN_6624;
      end
    end else begin
      reservedValidList1_59 <= _GEN_6624;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_60 <= _GEN_6922;
          end else begin
            reservedValidList1_60 <= PRFValidList_60; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_60 <= _GEN_6625;
        end
      end else begin
        reservedValidList1_60 <= _GEN_6625;
      end
    end else begin
      reservedValidList1_60 <= _GEN_6625;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_61 <= _GEN_6923;
          end else begin
            reservedValidList1_61 <= PRFValidList_61; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_61 <= _GEN_6626;
        end
      end else begin
        reservedValidList1_61 <= _GEN_6626;
      end
    end else begin
      reservedValidList1_61 <= _GEN_6626;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_62 <= _GEN_6924;
          end else begin
            reservedValidList1_62 <= PRFValidList_62; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_62 <= _GEN_6627;
        end
      end else begin
        reservedValidList1_62 <= _GEN_6627;
      end
    end else begin
      reservedValidList1_62 <= _GEN_6627;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 436:44]
            reservedValidList1_63 <= _GEN_6925;
          end else begin
            reservedValidList1_63 <= PRFValidList_63; // @[decode.scala 435:30]
          end
        end else begin
          reservedValidList1_63 <= _GEN_6628;
        end
      end else begin
        reservedValidList1_63 <= _GEN_6628;
      end
    end else begin
      reservedValidList1_63 <= _GEN_6628;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_0 <= _GEN_6629;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_0 <= _GEN_7022;
        end else begin
          reservedValidList2_0 <= _GEN_6629;
        end
      end else begin
        reservedValidList2_0 <= _GEN_6629;
      end
    end else begin
      reservedValidList2_0 <= _GEN_6629;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_1 <= _GEN_6630;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_1 <= _GEN_7023;
        end else begin
          reservedValidList2_1 <= _GEN_6630;
        end
      end else begin
        reservedValidList2_1 <= _GEN_6630;
      end
    end else begin
      reservedValidList2_1 <= _GEN_6630;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_2 <= _GEN_6631;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_2 <= _GEN_7024;
        end else begin
          reservedValidList2_2 <= _GEN_6631;
        end
      end else begin
        reservedValidList2_2 <= _GEN_6631;
      end
    end else begin
      reservedValidList2_2 <= _GEN_6631;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_3 <= _GEN_6632;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_3 <= _GEN_7025;
        end else begin
          reservedValidList2_3 <= _GEN_6632;
        end
      end else begin
        reservedValidList2_3 <= _GEN_6632;
      end
    end else begin
      reservedValidList2_3 <= _GEN_6632;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_4 <= _GEN_6633;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_4 <= _GEN_7026;
        end else begin
          reservedValidList2_4 <= _GEN_6633;
        end
      end else begin
        reservedValidList2_4 <= _GEN_6633;
      end
    end else begin
      reservedValidList2_4 <= _GEN_6633;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_5 <= _GEN_6634;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_5 <= _GEN_7027;
        end else begin
          reservedValidList2_5 <= _GEN_6634;
        end
      end else begin
        reservedValidList2_5 <= _GEN_6634;
      end
    end else begin
      reservedValidList2_5 <= _GEN_6634;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_6 <= _GEN_6635;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_6 <= _GEN_7028;
        end else begin
          reservedValidList2_6 <= _GEN_6635;
        end
      end else begin
        reservedValidList2_6 <= _GEN_6635;
      end
    end else begin
      reservedValidList2_6 <= _GEN_6635;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_7 <= _GEN_6636;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_7 <= _GEN_7029;
        end else begin
          reservedValidList2_7 <= _GEN_6636;
        end
      end else begin
        reservedValidList2_7 <= _GEN_6636;
      end
    end else begin
      reservedValidList2_7 <= _GEN_6636;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_8 <= _GEN_6637;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_8 <= _GEN_7030;
        end else begin
          reservedValidList2_8 <= _GEN_6637;
        end
      end else begin
        reservedValidList2_8 <= _GEN_6637;
      end
    end else begin
      reservedValidList2_8 <= _GEN_6637;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_9 <= _GEN_6638;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_9 <= _GEN_7031;
        end else begin
          reservedValidList2_9 <= _GEN_6638;
        end
      end else begin
        reservedValidList2_9 <= _GEN_6638;
      end
    end else begin
      reservedValidList2_9 <= _GEN_6638;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_10 <= _GEN_6639;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_10 <= _GEN_7032;
        end else begin
          reservedValidList2_10 <= _GEN_6639;
        end
      end else begin
        reservedValidList2_10 <= _GEN_6639;
      end
    end else begin
      reservedValidList2_10 <= _GEN_6639;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_11 <= _GEN_6640;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_11 <= _GEN_7033;
        end else begin
          reservedValidList2_11 <= _GEN_6640;
        end
      end else begin
        reservedValidList2_11 <= _GEN_6640;
      end
    end else begin
      reservedValidList2_11 <= _GEN_6640;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_12 <= _GEN_6641;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_12 <= _GEN_7034;
        end else begin
          reservedValidList2_12 <= _GEN_6641;
        end
      end else begin
        reservedValidList2_12 <= _GEN_6641;
      end
    end else begin
      reservedValidList2_12 <= _GEN_6641;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_13 <= _GEN_6642;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_13 <= _GEN_7035;
        end else begin
          reservedValidList2_13 <= _GEN_6642;
        end
      end else begin
        reservedValidList2_13 <= _GEN_6642;
      end
    end else begin
      reservedValidList2_13 <= _GEN_6642;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_14 <= _GEN_6643;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_14 <= _GEN_7036;
        end else begin
          reservedValidList2_14 <= _GEN_6643;
        end
      end else begin
        reservedValidList2_14 <= _GEN_6643;
      end
    end else begin
      reservedValidList2_14 <= _GEN_6643;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_15 <= _GEN_6644;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_15 <= _GEN_7037;
        end else begin
          reservedValidList2_15 <= _GEN_6644;
        end
      end else begin
        reservedValidList2_15 <= _GEN_6644;
      end
    end else begin
      reservedValidList2_15 <= _GEN_6644;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_16 <= _GEN_6645;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_16 <= _GEN_7038;
        end else begin
          reservedValidList2_16 <= _GEN_6645;
        end
      end else begin
        reservedValidList2_16 <= _GEN_6645;
      end
    end else begin
      reservedValidList2_16 <= _GEN_6645;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_17 <= _GEN_6646;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_17 <= _GEN_7039;
        end else begin
          reservedValidList2_17 <= _GEN_6646;
        end
      end else begin
        reservedValidList2_17 <= _GEN_6646;
      end
    end else begin
      reservedValidList2_17 <= _GEN_6646;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_18 <= _GEN_6647;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_18 <= _GEN_7040;
        end else begin
          reservedValidList2_18 <= _GEN_6647;
        end
      end else begin
        reservedValidList2_18 <= _GEN_6647;
      end
    end else begin
      reservedValidList2_18 <= _GEN_6647;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_19 <= _GEN_6648;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_19 <= _GEN_7041;
        end else begin
          reservedValidList2_19 <= _GEN_6648;
        end
      end else begin
        reservedValidList2_19 <= _GEN_6648;
      end
    end else begin
      reservedValidList2_19 <= _GEN_6648;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_20 <= _GEN_6649;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_20 <= _GEN_7042;
        end else begin
          reservedValidList2_20 <= _GEN_6649;
        end
      end else begin
        reservedValidList2_20 <= _GEN_6649;
      end
    end else begin
      reservedValidList2_20 <= _GEN_6649;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_21 <= _GEN_6650;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_21 <= _GEN_7043;
        end else begin
          reservedValidList2_21 <= _GEN_6650;
        end
      end else begin
        reservedValidList2_21 <= _GEN_6650;
      end
    end else begin
      reservedValidList2_21 <= _GEN_6650;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_22 <= _GEN_6651;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_22 <= _GEN_7044;
        end else begin
          reservedValidList2_22 <= _GEN_6651;
        end
      end else begin
        reservedValidList2_22 <= _GEN_6651;
      end
    end else begin
      reservedValidList2_22 <= _GEN_6651;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_23 <= _GEN_6652;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_23 <= _GEN_7045;
        end else begin
          reservedValidList2_23 <= _GEN_6652;
        end
      end else begin
        reservedValidList2_23 <= _GEN_6652;
      end
    end else begin
      reservedValidList2_23 <= _GEN_6652;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_24 <= _GEN_6653;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_24 <= _GEN_7046;
        end else begin
          reservedValidList2_24 <= _GEN_6653;
        end
      end else begin
        reservedValidList2_24 <= _GEN_6653;
      end
    end else begin
      reservedValidList2_24 <= _GEN_6653;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_25 <= _GEN_6654;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_25 <= _GEN_7047;
        end else begin
          reservedValidList2_25 <= _GEN_6654;
        end
      end else begin
        reservedValidList2_25 <= _GEN_6654;
      end
    end else begin
      reservedValidList2_25 <= _GEN_6654;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_26 <= _GEN_6655;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_26 <= _GEN_7048;
        end else begin
          reservedValidList2_26 <= _GEN_6655;
        end
      end else begin
        reservedValidList2_26 <= _GEN_6655;
      end
    end else begin
      reservedValidList2_26 <= _GEN_6655;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_27 <= _GEN_6656;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_27 <= _GEN_7049;
        end else begin
          reservedValidList2_27 <= _GEN_6656;
        end
      end else begin
        reservedValidList2_27 <= _GEN_6656;
      end
    end else begin
      reservedValidList2_27 <= _GEN_6656;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_28 <= _GEN_6657;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_28 <= _GEN_7050;
        end else begin
          reservedValidList2_28 <= _GEN_6657;
        end
      end else begin
        reservedValidList2_28 <= _GEN_6657;
      end
    end else begin
      reservedValidList2_28 <= _GEN_6657;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_29 <= _GEN_6658;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_29 <= _GEN_7051;
        end else begin
          reservedValidList2_29 <= _GEN_6658;
        end
      end else begin
        reservedValidList2_29 <= _GEN_6658;
      end
    end else begin
      reservedValidList2_29 <= _GEN_6658;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_30 <= _GEN_6659;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_30 <= _GEN_7052;
        end else begin
          reservedValidList2_30 <= _GEN_6659;
        end
      end else begin
        reservedValidList2_30 <= _GEN_6659;
      end
    end else begin
      reservedValidList2_30 <= _GEN_6659;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_31 <= _GEN_6660;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_31 <= _GEN_7053;
        end else begin
          reservedValidList2_31 <= _GEN_6660;
        end
      end else begin
        reservedValidList2_31 <= _GEN_6660;
      end
    end else begin
      reservedValidList2_31 <= _GEN_6660;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_32 <= _GEN_6661;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_32 <= _GEN_7054;
        end else begin
          reservedValidList2_32 <= _GEN_6661;
        end
      end else begin
        reservedValidList2_32 <= _GEN_6661;
      end
    end else begin
      reservedValidList2_32 <= _GEN_6661;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_33 <= _GEN_6662;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_33 <= _GEN_7055;
        end else begin
          reservedValidList2_33 <= _GEN_6662;
        end
      end else begin
        reservedValidList2_33 <= _GEN_6662;
      end
    end else begin
      reservedValidList2_33 <= _GEN_6662;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_34 <= _GEN_6663;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_34 <= _GEN_7056;
        end else begin
          reservedValidList2_34 <= _GEN_6663;
        end
      end else begin
        reservedValidList2_34 <= _GEN_6663;
      end
    end else begin
      reservedValidList2_34 <= _GEN_6663;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_35 <= _GEN_6664;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_35 <= _GEN_7057;
        end else begin
          reservedValidList2_35 <= _GEN_6664;
        end
      end else begin
        reservedValidList2_35 <= _GEN_6664;
      end
    end else begin
      reservedValidList2_35 <= _GEN_6664;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_36 <= _GEN_6665;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_36 <= _GEN_7058;
        end else begin
          reservedValidList2_36 <= _GEN_6665;
        end
      end else begin
        reservedValidList2_36 <= _GEN_6665;
      end
    end else begin
      reservedValidList2_36 <= _GEN_6665;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_37 <= _GEN_6666;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_37 <= _GEN_7059;
        end else begin
          reservedValidList2_37 <= _GEN_6666;
        end
      end else begin
        reservedValidList2_37 <= _GEN_6666;
      end
    end else begin
      reservedValidList2_37 <= _GEN_6666;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_38 <= _GEN_6667;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_38 <= _GEN_7060;
        end else begin
          reservedValidList2_38 <= _GEN_6667;
        end
      end else begin
        reservedValidList2_38 <= _GEN_6667;
      end
    end else begin
      reservedValidList2_38 <= _GEN_6667;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_39 <= _GEN_6668;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_39 <= _GEN_7061;
        end else begin
          reservedValidList2_39 <= _GEN_6668;
        end
      end else begin
        reservedValidList2_39 <= _GEN_6668;
      end
    end else begin
      reservedValidList2_39 <= _GEN_6668;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_40 <= _GEN_6669;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_40 <= _GEN_7062;
        end else begin
          reservedValidList2_40 <= _GEN_6669;
        end
      end else begin
        reservedValidList2_40 <= _GEN_6669;
      end
    end else begin
      reservedValidList2_40 <= _GEN_6669;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_41 <= _GEN_6670;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_41 <= _GEN_7063;
        end else begin
          reservedValidList2_41 <= _GEN_6670;
        end
      end else begin
        reservedValidList2_41 <= _GEN_6670;
      end
    end else begin
      reservedValidList2_41 <= _GEN_6670;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_42 <= _GEN_6671;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_42 <= _GEN_7064;
        end else begin
          reservedValidList2_42 <= _GEN_6671;
        end
      end else begin
        reservedValidList2_42 <= _GEN_6671;
      end
    end else begin
      reservedValidList2_42 <= _GEN_6671;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_43 <= _GEN_6672;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_43 <= _GEN_7065;
        end else begin
          reservedValidList2_43 <= _GEN_6672;
        end
      end else begin
        reservedValidList2_43 <= _GEN_6672;
      end
    end else begin
      reservedValidList2_43 <= _GEN_6672;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_44 <= _GEN_6673;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_44 <= _GEN_7066;
        end else begin
          reservedValidList2_44 <= _GEN_6673;
        end
      end else begin
        reservedValidList2_44 <= _GEN_6673;
      end
    end else begin
      reservedValidList2_44 <= _GEN_6673;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_45 <= _GEN_6674;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_45 <= _GEN_7067;
        end else begin
          reservedValidList2_45 <= _GEN_6674;
        end
      end else begin
        reservedValidList2_45 <= _GEN_6674;
      end
    end else begin
      reservedValidList2_45 <= _GEN_6674;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_46 <= _GEN_6675;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_46 <= _GEN_7068;
        end else begin
          reservedValidList2_46 <= _GEN_6675;
        end
      end else begin
        reservedValidList2_46 <= _GEN_6675;
      end
    end else begin
      reservedValidList2_46 <= _GEN_6675;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_47 <= _GEN_6676;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_47 <= _GEN_7069;
        end else begin
          reservedValidList2_47 <= _GEN_6676;
        end
      end else begin
        reservedValidList2_47 <= _GEN_6676;
      end
    end else begin
      reservedValidList2_47 <= _GEN_6676;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_48 <= _GEN_6677;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_48 <= _GEN_7070;
        end else begin
          reservedValidList2_48 <= _GEN_6677;
        end
      end else begin
        reservedValidList2_48 <= _GEN_6677;
      end
    end else begin
      reservedValidList2_48 <= _GEN_6677;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_49 <= _GEN_6678;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_49 <= _GEN_7071;
        end else begin
          reservedValidList2_49 <= _GEN_6678;
        end
      end else begin
        reservedValidList2_49 <= _GEN_6678;
      end
    end else begin
      reservedValidList2_49 <= _GEN_6678;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_50 <= _GEN_6679;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_50 <= _GEN_7072;
        end else begin
          reservedValidList2_50 <= _GEN_6679;
        end
      end else begin
        reservedValidList2_50 <= _GEN_6679;
      end
    end else begin
      reservedValidList2_50 <= _GEN_6679;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_51 <= _GEN_6680;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_51 <= _GEN_7073;
        end else begin
          reservedValidList2_51 <= _GEN_6680;
        end
      end else begin
        reservedValidList2_51 <= _GEN_6680;
      end
    end else begin
      reservedValidList2_51 <= _GEN_6680;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_52 <= _GEN_6681;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_52 <= _GEN_7074;
        end else begin
          reservedValidList2_52 <= _GEN_6681;
        end
      end else begin
        reservedValidList2_52 <= _GEN_6681;
      end
    end else begin
      reservedValidList2_52 <= _GEN_6681;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_53 <= _GEN_6682;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_53 <= _GEN_7075;
        end else begin
          reservedValidList2_53 <= _GEN_6682;
        end
      end else begin
        reservedValidList2_53 <= _GEN_6682;
      end
    end else begin
      reservedValidList2_53 <= _GEN_6682;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_54 <= _GEN_6683;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_54 <= _GEN_7076;
        end else begin
          reservedValidList2_54 <= _GEN_6683;
        end
      end else begin
        reservedValidList2_54 <= _GEN_6683;
      end
    end else begin
      reservedValidList2_54 <= _GEN_6683;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_55 <= _GEN_6684;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_55 <= _GEN_7077;
        end else begin
          reservedValidList2_55 <= _GEN_6684;
        end
      end else begin
        reservedValidList2_55 <= _GEN_6684;
      end
    end else begin
      reservedValidList2_55 <= _GEN_6684;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_56 <= _GEN_6685;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_56 <= _GEN_7078;
        end else begin
          reservedValidList2_56 <= _GEN_6685;
        end
      end else begin
        reservedValidList2_56 <= _GEN_6685;
      end
    end else begin
      reservedValidList2_56 <= _GEN_6685;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_57 <= _GEN_6686;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_57 <= _GEN_7079;
        end else begin
          reservedValidList2_57 <= _GEN_6686;
        end
      end else begin
        reservedValidList2_57 <= _GEN_6686;
      end
    end else begin
      reservedValidList2_57 <= _GEN_6686;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_58 <= _GEN_6687;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_58 <= _GEN_7080;
        end else begin
          reservedValidList2_58 <= _GEN_6687;
        end
      end else begin
        reservedValidList2_58 <= _GEN_6687;
      end
    end else begin
      reservedValidList2_58 <= _GEN_6687;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_59 <= _GEN_6688;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_59 <= _GEN_7081;
        end else begin
          reservedValidList2_59 <= _GEN_6688;
        end
      end else begin
        reservedValidList2_59 <= _GEN_6688;
      end
    end else begin
      reservedValidList2_59 <= _GEN_6688;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_60 <= _GEN_6689;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_60 <= _GEN_7082;
        end else begin
          reservedValidList2_60 <= _GEN_6689;
        end
      end else begin
        reservedValidList2_60 <= _GEN_6689;
      end
    end else begin
      reservedValidList2_60 <= _GEN_6689;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_61 <= _GEN_6690;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_61 <= _GEN_7083;
        end else begin
          reservedValidList2_61 <= _GEN_6690;
        end
      end else begin
        reservedValidList2_61 <= _GEN_6690;
      end
    end else begin
      reservedValidList2_61 <= _GEN_6690;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_62 <= _GEN_6691;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_62 <= _GEN_7084;
        end else begin
          reservedValidList2_62 <= _GEN_6691;
        end
      end else begin
        reservedValidList2_62 <= _GEN_6691;
      end
    end else begin
      reservedValidList2_62 <= _GEN_6691;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_63 <= _GEN_6692;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList2_63 <= _GEN_7085;
        end else begin
          reservedValidList2_63 <= _GEN_6692;
        end
      end else begin
        reservedValidList2_63 <= _GEN_6692;
      end
    end else begin
      reservedValidList2_63 <= _GEN_6692;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_0 <= _GEN_6693;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_0 <= _GEN_6693;
        end else begin
          reservedValidList3_0 <= _GEN_8302;
        end
      end else begin
        reservedValidList3_0 <= _GEN_6693;
      end
    end else begin
      reservedValidList3_0 <= _GEN_6693;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_1 <= _GEN_6694;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_1 <= _GEN_6694;
        end else begin
          reservedValidList3_1 <= _GEN_8303;
        end
      end else begin
        reservedValidList3_1 <= _GEN_6694;
      end
    end else begin
      reservedValidList3_1 <= _GEN_6694;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_2 <= _GEN_6695;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_2 <= _GEN_6695;
        end else begin
          reservedValidList3_2 <= _GEN_8304;
        end
      end else begin
        reservedValidList3_2 <= _GEN_6695;
      end
    end else begin
      reservedValidList3_2 <= _GEN_6695;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_3 <= _GEN_6696;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_3 <= _GEN_6696;
        end else begin
          reservedValidList3_3 <= _GEN_8305;
        end
      end else begin
        reservedValidList3_3 <= _GEN_6696;
      end
    end else begin
      reservedValidList3_3 <= _GEN_6696;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_4 <= _GEN_6697;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_4 <= _GEN_6697;
        end else begin
          reservedValidList3_4 <= _GEN_8306;
        end
      end else begin
        reservedValidList3_4 <= _GEN_6697;
      end
    end else begin
      reservedValidList3_4 <= _GEN_6697;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_5 <= _GEN_6698;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_5 <= _GEN_6698;
        end else begin
          reservedValidList3_5 <= _GEN_8307;
        end
      end else begin
        reservedValidList3_5 <= _GEN_6698;
      end
    end else begin
      reservedValidList3_5 <= _GEN_6698;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_6 <= _GEN_6699;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_6 <= _GEN_6699;
        end else begin
          reservedValidList3_6 <= _GEN_8308;
        end
      end else begin
        reservedValidList3_6 <= _GEN_6699;
      end
    end else begin
      reservedValidList3_6 <= _GEN_6699;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_7 <= _GEN_6700;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_7 <= _GEN_6700;
        end else begin
          reservedValidList3_7 <= _GEN_8309;
        end
      end else begin
        reservedValidList3_7 <= _GEN_6700;
      end
    end else begin
      reservedValidList3_7 <= _GEN_6700;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_8 <= _GEN_6701;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_8 <= _GEN_6701;
        end else begin
          reservedValidList3_8 <= _GEN_8310;
        end
      end else begin
        reservedValidList3_8 <= _GEN_6701;
      end
    end else begin
      reservedValidList3_8 <= _GEN_6701;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_9 <= _GEN_6702;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_9 <= _GEN_6702;
        end else begin
          reservedValidList3_9 <= _GEN_8311;
        end
      end else begin
        reservedValidList3_9 <= _GEN_6702;
      end
    end else begin
      reservedValidList3_9 <= _GEN_6702;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_10 <= _GEN_6703;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_10 <= _GEN_6703;
        end else begin
          reservedValidList3_10 <= _GEN_8312;
        end
      end else begin
        reservedValidList3_10 <= _GEN_6703;
      end
    end else begin
      reservedValidList3_10 <= _GEN_6703;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_11 <= _GEN_6704;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_11 <= _GEN_6704;
        end else begin
          reservedValidList3_11 <= _GEN_8313;
        end
      end else begin
        reservedValidList3_11 <= _GEN_6704;
      end
    end else begin
      reservedValidList3_11 <= _GEN_6704;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_12 <= _GEN_6705;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_12 <= _GEN_6705;
        end else begin
          reservedValidList3_12 <= _GEN_8314;
        end
      end else begin
        reservedValidList3_12 <= _GEN_6705;
      end
    end else begin
      reservedValidList3_12 <= _GEN_6705;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_13 <= _GEN_6706;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_13 <= _GEN_6706;
        end else begin
          reservedValidList3_13 <= _GEN_8315;
        end
      end else begin
        reservedValidList3_13 <= _GEN_6706;
      end
    end else begin
      reservedValidList3_13 <= _GEN_6706;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_14 <= _GEN_6707;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_14 <= _GEN_6707;
        end else begin
          reservedValidList3_14 <= _GEN_8316;
        end
      end else begin
        reservedValidList3_14 <= _GEN_6707;
      end
    end else begin
      reservedValidList3_14 <= _GEN_6707;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_15 <= _GEN_6708;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_15 <= _GEN_6708;
        end else begin
          reservedValidList3_15 <= _GEN_8317;
        end
      end else begin
        reservedValidList3_15 <= _GEN_6708;
      end
    end else begin
      reservedValidList3_15 <= _GEN_6708;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_16 <= _GEN_6709;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_16 <= _GEN_6709;
        end else begin
          reservedValidList3_16 <= _GEN_8318;
        end
      end else begin
        reservedValidList3_16 <= _GEN_6709;
      end
    end else begin
      reservedValidList3_16 <= _GEN_6709;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_17 <= _GEN_6710;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_17 <= _GEN_6710;
        end else begin
          reservedValidList3_17 <= _GEN_8319;
        end
      end else begin
        reservedValidList3_17 <= _GEN_6710;
      end
    end else begin
      reservedValidList3_17 <= _GEN_6710;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_18 <= _GEN_6711;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_18 <= _GEN_6711;
        end else begin
          reservedValidList3_18 <= _GEN_8320;
        end
      end else begin
        reservedValidList3_18 <= _GEN_6711;
      end
    end else begin
      reservedValidList3_18 <= _GEN_6711;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_19 <= _GEN_6712;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_19 <= _GEN_6712;
        end else begin
          reservedValidList3_19 <= _GEN_8321;
        end
      end else begin
        reservedValidList3_19 <= _GEN_6712;
      end
    end else begin
      reservedValidList3_19 <= _GEN_6712;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_20 <= _GEN_6713;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_20 <= _GEN_6713;
        end else begin
          reservedValidList3_20 <= _GEN_8322;
        end
      end else begin
        reservedValidList3_20 <= _GEN_6713;
      end
    end else begin
      reservedValidList3_20 <= _GEN_6713;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_21 <= _GEN_6714;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_21 <= _GEN_6714;
        end else begin
          reservedValidList3_21 <= _GEN_8323;
        end
      end else begin
        reservedValidList3_21 <= _GEN_6714;
      end
    end else begin
      reservedValidList3_21 <= _GEN_6714;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_22 <= _GEN_6715;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_22 <= _GEN_6715;
        end else begin
          reservedValidList3_22 <= _GEN_8324;
        end
      end else begin
        reservedValidList3_22 <= _GEN_6715;
      end
    end else begin
      reservedValidList3_22 <= _GEN_6715;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_23 <= _GEN_6716;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_23 <= _GEN_6716;
        end else begin
          reservedValidList3_23 <= _GEN_8325;
        end
      end else begin
        reservedValidList3_23 <= _GEN_6716;
      end
    end else begin
      reservedValidList3_23 <= _GEN_6716;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_24 <= _GEN_6717;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_24 <= _GEN_6717;
        end else begin
          reservedValidList3_24 <= _GEN_8326;
        end
      end else begin
        reservedValidList3_24 <= _GEN_6717;
      end
    end else begin
      reservedValidList3_24 <= _GEN_6717;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_25 <= _GEN_6718;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_25 <= _GEN_6718;
        end else begin
          reservedValidList3_25 <= _GEN_8327;
        end
      end else begin
        reservedValidList3_25 <= _GEN_6718;
      end
    end else begin
      reservedValidList3_25 <= _GEN_6718;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_26 <= _GEN_6719;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_26 <= _GEN_6719;
        end else begin
          reservedValidList3_26 <= _GEN_8328;
        end
      end else begin
        reservedValidList3_26 <= _GEN_6719;
      end
    end else begin
      reservedValidList3_26 <= _GEN_6719;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_27 <= _GEN_6720;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_27 <= _GEN_6720;
        end else begin
          reservedValidList3_27 <= _GEN_8329;
        end
      end else begin
        reservedValidList3_27 <= _GEN_6720;
      end
    end else begin
      reservedValidList3_27 <= _GEN_6720;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_28 <= _GEN_6721;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_28 <= _GEN_6721;
        end else begin
          reservedValidList3_28 <= _GEN_8330;
        end
      end else begin
        reservedValidList3_28 <= _GEN_6721;
      end
    end else begin
      reservedValidList3_28 <= _GEN_6721;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_29 <= _GEN_6722;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_29 <= _GEN_6722;
        end else begin
          reservedValidList3_29 <= _GEN_8331;
        end
      end else begin
        reservedValidList3_29 <= _GEN_6722;
      end
    end else begin
      reservedValidList3_29 <= _GEN_6722;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_30 <= _GEN_6723;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_30 <= _GEN_6723;
        end else begin
          reservedValidList3_30 <= _GEN_8332;
        end
      end else begin
        reservedValidList3_30 <= _GEN_6723;
      end
    end else begin
      reservedValidList3_30 <= _GEN_6723;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_31 <= _GEN_6724;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_31 <= _GEN_6724;
        end else begin
          reservedValidList3_31 <= _GEN_8333;
        end
      end else begin
        reservedValidList3_31 <= _GEN_6724;
      end
    end else begin
      reservedValidList3_31 <= _GEN_6724;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_32 <= _GEN_6725;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_32 <= _GEN_6725;
        end else begin
          reservedValidList3_32 <= _GEN_8334;
        end
      end else begin
        reservedValidList3_32 <= _GEN_6725;
      end
    end else begin
      reservedValidList3_32 <= _GEN_6725;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_33 <= _GEN_6726;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_33 <= _GEN_6726;
        end else begin
          reservedValidList3_33 <= _GEN_8335;
        end
      end else begin
        reservedValidList3_33 <= _GEN_6726;
      end
    end else begin
      reservedValidList3_33 <= _GEN_6726;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_34 <= _GEN_6727;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_34 <= _GEN_6727;
        end else begin
          reservedValidList3_34 <= _GEN_8336;
        end
      end else begin
        reservedValidList3_34 <= _GEN_6727;
      end
    end else begin
      reservedValidList3_34 <= _GEN_6727;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_35 <= _GEN_6728;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_35 <= _GEN_6728;
        end else begin
          reservedValidList3_35 <= _GEN_8337;
        end
      end else begin
        reservedValidList3_35 <= _GEN_6728;
      end
    end else begin
      reservedValidList3_35 <= _GEN_6728;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_36 <= _GEN_6729;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_36 <= _GEN_6729;
        end else begin
          reservedValidList3_36 <= _GEN_8338;
        end
      end else begin
        reservedValidList3_36 <= _GEN_6729;
      end
    end else begin
      reservedValidList3_36 <= _GEN_6729;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_37 <= _GEN_6730;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_37 <= _GEN_6730;
        end else begin
          reservedValidList3_37 <= _GEN_8339;
        end
      end else begin
        reservedValidList3_37 <= _GEN_6730;
      end
    end else begin
      reservedValidList3_37 <= _GEN_6730;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_38 <= _GEN_6731;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_38 <= _GEN_6731;
        end else begin
          reservedValidList3_38 <= _GEN_8340;
        end
      end else begin
        reservedValidList3_38 <= _GEN_6731;
      end
    end else begin
      reservedValidList3_38 <= _GEN_6731;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_39 <= _GEN_6732;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_39 <= _GEN_6732;
        end else begin
          reservedValidList3_39 <= _GEN_8341;
        end
      end else begin
        reservedValidList3_39 <= _GEN_6732;
      end
    end else begin
      reservedValidList3_39 <= _GEN_6732;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_40 <= _GEN_6733;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_40 <= _GEN_6733;
        end else begin
          reservedValidList3_40 <= _GEN_8342;
        end
      end else begin
        reservedValidList3_40 <= _GEN_6733;
      end
    end else begin
      reservedValidList3_40 <= _GEN_6733;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_41 <= _GEN_6734;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_41 <= _GEN_6734;
        end else begin
          reservedValidList3_41 <= _GEN_8343;
        end
      end else begin
        reservedValidList3_41 <= _GEN_6734;
      end
    end else begin
      reservedValidList3_41 <= _GEN_6734;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_42 <= _GEN_6735;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_42 <= _GEN_6735;
        end else begin
          reservedValidList3_42 <= _GEN_8344;
        end
      end else begin
        reservedValidList3_42 <= _GEN_6735;
      end
    end else begin
      reservedValidList3_42 <= _GEN_6735;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_43 <= _GEN_6736;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_43 <= _GEN_6736;
        end else begin
          reservedValidList3_43 <= _GEN_8345;
        end
      end else begin
        reservedValidList3_43 <= _GEN_6736;
      end
    end else begin
      reservedValidList3_43 <= _GEN_6736;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_44 <= _GEN_6737;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_44 <= _GEN_6737;
        end else begin
          reservedValidList3_44 <= _GEN_8346;
        end
      end else begin
        reservedValidList3_44 <= _GEN_6737;
      end
    end else begin
      reservedValidList3_44 <= _GEN_6737;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_45 <= _GEN_6738;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_45 <= _GEN_6738;
        end else begin
          reservedValidList3_45 <= _GEN_8347;
        end
      end else begin
        reservedValidList3_45 <= _GEN_6738;
      end
    end else begin
      reservedValidList3_45 <= _GEN_6738;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_46 <= _GEN_6739;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_46 <= _GEN_6739;
        end else begin
          reservedValidList3_46 <= _GEN_8348;
        end
      end else begin
        reservedValidList3_46 <= _GEN_6739;
      end
    end else begin
      reservedValidList3_46 <= _GEN_6739;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_47 <= _GEN_6740;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_47 <= _GEN_6740;
        end else begin
          reservedValidList3_47 <= _GEN_8349;
        end
      end else begin
        reservedValidList3_47 <= _GEN_6740;
      end
    end else begin
      reservedValidList3_47 <= _GEN_6740;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_48 <= _GEN_6741;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_48 <= _GEN_6741;
        end else begin
          reservedValidList3_48 <= _GEN_8350;
        end
      end else begin
        reservedValidList3_48 <= _GEN_6741;
      end
    end else begin
      reservedValidList3_48 <= _GEN_6741;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_49 <= _GEN_6742;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_49 <= _GEN_6742;
        end else begin
          reservedValidList3_49 <= _GEN_8351;
        end
      end else begin
        reservedValidList3_49 <= _GEN_6742;
      end
    end else begin
      reservedValidList3_49 <= _GEN_6742;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_50 <= _GEN_6743;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_50 <= _GEN_6743;
        end else begin
          reservedValidList3_50 <= _GEN_8352;
        end
      end else begin
        reservedValidList3_50 <= _GEN_6743;
      end
    end else begin
      reservedValidList3_50 <= _GEN_6743;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_51 <= _GEN_6744;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_51 <= _GEN_6744;
        end else begin
          reservedValidList3_51 <= _GEN_8353;
        end
      end else begin
        reservedValidList3_51 <= _GEN_6744;
      end
    end else begin
      reservedValidList3_51 <= _GEN_6744;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_52 <= _GEN_6745;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_52 <= _GEN_6745;
        end else begin
          reservedValidList3_52 <= _GEN_8354;
        end
      end else begin
        reservedValidList3_52 <= _GEN_6745;
      end
    end else begin
      reservedValidList3_52 <= _GEN_6745;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_53 <= _GEN_6746;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_53 <= _GEN_6746;
        end else begin
          reservedValidList3_53 <= _GEN_8355;
        end
      end else begin
        reservedValidList3_53 <= _GEN_6746;
      end
    end else begin
      reservedValidList3_53 <= _GEN_6746;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_54 <= _GEN_6747;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_54 <= _GEN_6747;
        end else begin
          reservedValidList3_54 <= _GEN_8356;
        end
      end else begin
        reservedValidList3_54 <= _GEN_6747;
      end
    end else begin
      reservedValidList3_54 <= _GEN_6747;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_55 <= _GEN_6748;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_55 <= _GEN_6748;
        end else begin
          reservedValidList3_55 <= _GEN_8357;
        end
      end else begin
        reservedValidList3_55 <= _GEN_6748;
      end
    end else begin
      reservedValidList3_55 <= _GEN_6748;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_56 <= _GEN_6749;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_56 <= _GEN_6749;
        end else begin
          reservedValidList3_56 <= _GEN_8358;
        end
      end else begin
        reservedValidList3_56 <= _GEN_6749;
      end
    end else begin
      reservedValidList3_56 <= _GEN_6749;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_57 <= _GEN_6750;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_57 <= _GEN_6750;
        end else begin
          reservedValidList3_57 <= _GEN_8359;
        end
      end else begin
        reservedValidList3_57 <= _GEN_6750;
      end
    end else begin
      reservedValidList3_57 <= _GEN_6750;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_58 <= _GEN_6751;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_58 <= _GEN_6751;
        end else begin
          reservedValidList3_58 <= _GEN_8360;
        end
      end else begin
        reservedValidList3_58 <= _GEN_6751;
      end
    end else begin
      reservedValidList3_58 <= _GEN_6751;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_59 <= _GEN_6752;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_59 <= _GEN_6752;
        end else begin
          reservedValidList3_59 <= _GEN_8361;
        end
      end else begin
        reservedValidList3_59 <= _GEN_6752;
      end
    end else begin
      reservedValidList3_59 <= _GEN_6752;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_60 <= _GEN_6753;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_60 <= _GEN_6753;
        end else begin
          reservedValidList3_60 <= _GEN_8362;
        end
      end else begin
        reservedValidList3_60 <= _GEN_6753;
      end
    end else begin
      reservedValidList3_60 <= _GEN_6753;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_61 <= _GEN_6754;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_61 <= _GEN_6754;
        end else begin
          reservedValidList3_61 <= _GEN_8363;
        end
      end else begin
        reservedValidList3_61 <= _GEN_6754;
      end
    end else begin
      reservedValidList3_61 <= _GEN_6754;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_62 <= _GEN_6755;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_62 <= _GEN_6755;
        end else begin
          reservedValidList3_62 <= _GEN_8364;
        end
      end else begin
        reservedValidList3_62 <= _GEN_6755;
      end
    end else begin
      reservedValidList3_62 <= _GEN_6755;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_63 <= _GEN_6756;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 431:29]
          reservedValidList3_63 <= _GEN_6756;
        end else begin
          reservedValidList3_63 <= _GEN_8365;
        end
      end else begin
        reservedValidList3_63 <= _GEN_6756;
      end
    end else begin
      reservedValidList3_63 <= _GEN_6756;
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_0 <= _GEN_8462;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_1 <= _GEN_8463;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_2 <= _GEN_8464;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_3 <= _GEN_8465;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_4 <= _GEN_8466;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_5 <= _GEN_8467;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_6 <= _GEN_8468;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_7 <= _GEN_8469;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_8 <= _GEN_8470;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_9 <= _GEN_8471;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_10 <= _GEN_8472;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_11 <= _GEN_8473;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_12 <= _GEN_8474;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_13 <= _GEN_8475;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_14 <= _GEN_8476;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_15 <= _GEN_8477;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_16 <= _GEN_8478;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_17 <= _GEN_8479;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_18 <= _GEN_8480;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_19 <= _GEN_8481;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_20 <= _GEN_8482;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_21 <= _GEN_8483;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_22 <= _GEN_8484;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_23 <= _GEN_8485;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_24 <= _GEN_8486;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_25 <= _GEN_8487;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_26 <= _GEN_8488;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_27 <= _GEN_8489;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_28 <= _GEN_8490;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_29 <= _GEN_8491;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_30 <= _GEN_8492;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_31 <= _GEN_8493;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_32 <= _GEN_8494;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_33 <= _GEN_8495;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_34 <= _GEN_8496;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_35 <= _GEN_8497;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_36 <= _GEN_8498;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_37 <= _GEN_8499;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_38 <= _GEN_8500;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_39 <= _GEN_8501;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_40 <= _GEN_8502;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_41 <= _GEN_8503;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_42 <= _GEN_8504;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_43 <= _GEN_8505;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_44 <= _GEN_8506;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_45 <= _GEN_8507;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_46 <= _GEN_8508;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_47 <= _GEN_8509;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_48 <= _GEN_8510;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_49 <= _GEN_8511;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_50 <= _GEN_8512;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_51 <= _GEN_8513;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_52 <= _GEN_8514;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_53 <= _GEN_8515;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_54 <= _GEN_8516;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_55 <= _GEN_8517;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_56 <= _GEN_8518;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_57 <= _GEN_8519;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_58 <= _GEN_8520;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_59 <= _GEN_8521;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_60 <= _GEN_8522;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_61 <= _GEN_8523;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_62 <= _GEN_8524;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 419:41]
      if (_T_442 | _T_444 | _T_441) begin // @[decode.scala 420:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 431:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 431:29]
            reservedValidList4_63 <= _GEN_8525;
          end
        end
      end
    end
    if (reset) begin // @[decode.scala 497:28]
      ustatus <= 64'h0; // @[decode.scala 497:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (12'h0 == csrAddrReg) begin // @[decode.scala 573:39]
          ustatus <= csrWriteData; // @[decode.scala 574:37]
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        ustatus <= _GEN_11556;
      end else begin
        ustatus <= _GEN_12852;
      end
    end
    if (reset) begin // @[decode.scala 498:28]
      utvec <= 64'h0; // @[decode.scala 498:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 573:39]
          utvec <= _GEN_11233;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        utvec <= _GEN_11557;
      end else begin
        utvec <= _GEN_12853;
      end
    end
    if (reset) begin // @[decode.scala 499:28]
      uepc <= 64'h0; // @[decode.scala 499:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 573:39]
          uepc <= _GEN_11234;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        uepc <= _GEN_11558;
      end else begin
        uepc <= _GEN_12854;
      end
    end
    if (reset) begin // @[decode.scala 500:28]
      ucause <= 64'h0; // @[decode.scala 500:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 573:39]
          ucause <= _GEN_11235;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        ucause <= _GEN_11559;
      end else begin
        ucause <= _GEN_12855;
      end
    end
    if (reset) begin // @[decode.scala 501:28]
      scounteren <= 64'h0; // @[decode.scala 501:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 573:39]
          scounteren <= _GEN_11236;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        scounteren <= _GEN_11560;
      end else begin
        scounteren <= _GEN_12856;
      end
    end
    if (reset) begin // @[decode.scala 502:28]
      satp <= 64'h0; // @[decode.scala 502:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 573:39]
          satp <= _GEN_11237;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        satp <= _GEN_11561;
      end else begin
        satp <= _GEN_12857;
      end
    end
    if (reset) begin // @[decode.scala 503:28]
      mstatus <= 64'h0; // @[decode.scala 503:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] == 3'h0) begin // @[decode.scala 744:126]
      if (writeBackResult_instruction[31:20] == 12'h302) begin // @[decode.scala 745:60]
        mstatus <= _mstatus_T_9; // @[decode.scala 749:15]
      end else if (~(|writeBackResult_instruction[31:20])) begin // @[decode.scala 750:58]
        mstatus <= _mstatus_T_14; // @[decode.scala 757:15]
      end else begin
        mstatus <= _GEN_12956;
      end
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        mstatus <= _GEN_11262;
      end else begin
        mstatus <= _GEN_12882;
      end
    end else begin
      mstatus <= _mstatus_T_1; // @[decode.scala 522:11]
    end
    misa <= _GEN_16610[63:0]; // @[decode.scala 504:{28,28}]
    if (reset) begin // @[decode.scala 505:28]
      medeleg <= 64'h0; // @[decode.scala 505:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 573:39]
          medeleg <= _GEN_11240;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        medeleg <= _GEN_11564;
      end else begin
        medeleg <= _GEN_12860;
      end
    end
    if (reset) begin // @[decode.scala 506:28]
      mideleg <= 64'h0; // @[decode.scala 506:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 573:39]
          mideleg <= _GEN_11241;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        mideleg <= _GEN_11565;
      end else begin
        mideleg <= _GEN_12861;
      end
    end
    if (reset) begin // @[decode.scala 507:28]
      mie <= 64'h0; // @[decode.scala 507:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 573:39]
          mie <= _GEN_11242;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        mie <= _GEN_11566;
      end else begin
        mie <= _GEN_12862;
      end
    end
    if (reset) begin // @[decode.scala 508:28]
      mtvec <= 64'h0; // @[decode.scala 508:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 573:39]
          mtvec <= _GEN_11243;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        mtvec <= _GEN_11567;
      end else begin
        mtvec <= _GEN_12863;
      end
    end
    if (reset) begin // @[decode.scala 509:28]
      mcounteren <= 64'h0; // @[decode.scala 509:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 573:39]
          mcounteren <= _GEN_11244;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        mcounteren <= _GEN_11568;
      end else begin
        mcounteren <= _GEN_12864;
      end
    end
    if (reset) begin // @[decode.scala 510:28]
      mscratch <= 64'h0; // @[decode.scala 510:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 573:39]
          mscratch <= _GEN_11245;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        mscratch <= _GEN_11569;
      end else begin
        mscratch <= _GEN_12865;
      end
    end
    if (reset) begin // @[decode.scala 511:28]
      mepc <= 64'h0; // @[decode.scala 511:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] == 3'h0) begin // @[decode.scala 744:126]
      if (writeBackResult_instruction[31:20] == 12'h302) begin // @[decode.scala 745:60]
        mepc <= _GEN_12939;
      end else if (~(|writeBackResult_instruction[31:20])) begin // @[decode.scala 750:58]
        mepc <= ecallPC; // @[decode.scala 752:12]
      end else begin
        mepc <= _GEN_12952;
      end
    end else begin
      mepc <= _GEN_12939;
    end
    if (reset) begin // @[decode.scala 512:28]
      mcause <= 64'h0; // @[decode.scala 512:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] == 3'h0) begin // @[decode.scala 744:126]
      if (writeBackResult_instruction[31:20] == 12'h302) begin // @[decode.scala 745:60]
        mcause <= _GEN_12940;
      end else if (~(|writeBackResult_instruction[31:20])) begin // @[decode.scala 750:58]
        mcause <= {{60'd0}, _GEN_12951};
      end else begin
        mcause <= _GEN_12953;
      end
    end else begin
      mcause <= _GEN_12940;
    end
    if (reset) begin // @[decode.scala 513:28]
      mtval <= 64'h0; // @[decode.scala 513:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 573:39]
          mtval <= _GEN_11248;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        mtval <= _GEN_11572;
      end else begin
        mtval <= _GEN_12868;
      end
    end
    if (reset) begin // @[decode.scala 514:28]
      mip <= 64'h0; // @[decode.scala 514:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 573:39]
          mip <= _GEN_11249;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        mip <= _GEN_11573;
      end else begin
        mip <= _GEN_12869;
      end
    end
    if (reset) begin // @[decode.scala 515:28]
      pmpcfg0 <= 64'h0; // @[decode.scala 515:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 573:39]
          pmpcfg0 <= _GEN_11250;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        pmpcfg0 <= _GEN_11574;
      end else begin
        pmpcfg0 <= _GEN_12870;
      end
    end
    if (reset) begin // @[decode.scala 516:28]
      pmpaddr0 <= 64'h0; // @[decode.scala 516:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 573:39]
          pmpaddr0 <= _GEN_11251;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        pmpaddr0 <= _GEN_11575;
      end else begin
        pmpaddr0 <= _GEN_12871;
      end
    end
    if (reset) begin // @[decode.scala 517:28]
      mvendorid <= 64'h0; // @[decode.scala 517:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 573:39]
          mvendorid <= _GEN_11252;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        mvendorid <= _GEN_11576;
      end else begin
        mvendorid <= _GEN_12872;
      end
    end
    if (reset) begin // @[decode.scala 518:28]
      marchid <= 64'h0; // @[decode.scala 518:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 573:39]
          marchid <= _GEN_11253;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        marchid <= _GEN_11577;
      end else begin
        marchid <= _GEN_12873;
      end
    end
    if (reset) begin // @[decode.scala 519:28]
      mimpid <= 64'h0; // @[decode.scala 519:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 573:39]
          mimpid <= _GEN_11254;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        mimpid <= _GEN_11578;
      end else begin
        mimpid <= _GEN_12874;
      end
    end
    if (reset) begin // @[decode.scala 520:28]
      mhartid <= 64'h0; // @[decode.scala 520:28]
    end else if (_T_256 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 568:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 573:39]
          mhartid <= _GEN_11255;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 571:48]
        mhartid <= _GEN_11579;
      end else begin
        mhartid <= _GEN_12875;
      end
    end
    if (reset) begin // @[decode.scala 743:33]
      currentPrivilege <= 64'h2200000000; // @[decode.scala 743:33]
    end else if (_T_256 & writeBackResult_instruction[14:12] == 3'h0) begin // @[decode.scala 744:126]
      if (writeBackResult_instruction[31:20] == 12'h302) begin // @[decode.scala 745:60]
        currentPrivilege <= {{26'd0}, _GEN_12950}; // @[decode.scala 747:24]
      end else if (~(|writeBackResult_instruction[31:20])) begin // @[decode.scala 750:58]
        currentPrivilege <= 64'h2200000000; // @[decode.scala 755:24]
      end else begin
        currentPrivilege <= _GEN_12954;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  inputBuffer_pc = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  inputBuffer_instruction = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  outputBuffer_instruction = _RAND_2[31:0];
  _RAND_3 = {2{`RANDOM}};
  outputBuffer_pc = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  outputBuffer_PRFDest = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  outputBuffer_rs1Addr = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  outputBuffer_rs2Addr = _RAND_6[5:0];
  _RAND_7 = {2{`RANDOM}};
  outputBuffer_immediate = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  branchBuffer_branchPCReady = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  branchBuffer_predictedPCReady = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  branchBuffer_branchPC = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  branchBuffer_predictedPC = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  branchBuffer_branchMask_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  branchBuffer_branchMask_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  branchBuffer_branchMask_2 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  branchBuffer_branchMask_3 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  branchBuffer_branchMask_4 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  branchTracker = _RAND_17[2:0];
  _RAND_18 = {2{`RANDOM}};
  expectedPC = _RAND_18[63:0];
  _RAND_19 = {1{`RANDOM}};
  coherency = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  stateRegInputBuf = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  stateRegOutputBuf = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  stallReg = _RAND_22[0:0];
  _RAND_23 = {2{`RANDOM}};
  ecallPC = _RAND_23[63:0];
  _RAND_24 = {1{`RANDOM}};
  PRFValidList_0 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  PRFValidList_1 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  PRFValidList_2 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  PRFValidList_3 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  PRFValidList_4 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  PRFValidList_5 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  PRFValidList_6 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  PRFValidList_7 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  PRFValidList_8 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  PRFValidList_9 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  PRFValidList_10 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  PRFValidList_11 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  PRFValidList_12 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  PRFValidList_13 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  PRFValidList_14 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  PRFValidList_15 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  PRFValidList_16 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  PRFValidList_17 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  PRFValidList_18 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  PRFValidList_19 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  PRFValidList_20 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  PRFValidList_21 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  PRFValidList_22 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  PRFValidList_23 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  PRFValidList_24 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  PRFValidList_25 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  PRFValidList_26 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  PRFValidList_27 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  PRFValidList_28 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  PRFValidList_29 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  PRFValidList_30 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  PRFValidList_31 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  PRFValidList_32 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  PRFValidList_33 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  PRFValidList_34 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  PRFValidList_35 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  PRFValidList_36 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  PRFValidList_37 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  PRFValidList_38 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  PRFValidList_39 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  PRFValidList_40 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  PRFValidList_41 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  PRFValidList_42 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  PRFValidList_43 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  PRFValidList_44 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  PRFValidList_45 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  PRFValidList_46 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  PRFValidList_47 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  PRFValidList_48 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  PRFValidList_49 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  PRFValidList_50 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  PRFValidList_51 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  PRFValidList_52 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  PRFValidList_53 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  PRFValidList_54 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  PRFValidList_55 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  PRFValidList_56 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  PRFValidList_57 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  PRFValidList_58 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  PRFValidList_59 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  PRFValidList_60 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  PRFValidList_61 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  PRFValidList_62 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  PRFValidList_63 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  frontEndRegMap_31 = _RAND_88[5:0];
  _RAND_89 = {1{`RANDOM}};
  frontEndRegMap_30 = _RAND_89[5:0];
  _RAND_90 = {1{`RANDOM}};
  frontEndRegMap_29 = _RAND_90[5:0];
  _RAND_91 = {1{`RANDOM}};
  frontEndRegMap_28 = _RAND_91[5:0];
  _RAND_92 = {1{`RANDOM}};
  frontEndRegMap_27 = _RAND_92[5:0];
  _RAND_93 = {1{`RANDOM}};
  frontEndRegMap_26 = _RAND_93[5:0];
  _RAND_94 = {1{`RANDOM}};
  frontEndRegMap_25 = _RAND_94[5:0];
  _RAND_95 = {1{`RANDOM}};
  frontEndRegMap_24 = _RAND_95[5:0];
  _RAND_96 = {1{`RANDOM}};
  frontEndRegMap_23 = _RAND_96[5:0];
  _RAND_97 = {1{`RANDOM}};
  frontEndRegMap_22 = _RAND_97[5:0];
  _RAND_98 = {1{`RANDOM}};
  frontEndRegMap_21 = _RAND_98[5:0];
  _RAND_99 = {1{`RANDOM}};
  frontEndRegMap_20 = _RAND_99[5:0];
  _RAND_100 = {1{`RANDOM}};
  frontEndRegMap_19 = _RAND_100[5:0];
  _RAND_101 = {1{`RANDOM}};
  frontEndRegMap_18 = _RAND_101[5:0];
  _RAND_102 = {1{`RANDOM}};
  frontEndRegMap_17 = _RAND_102[5:0];
  _RAND_103 = {1{`RANDOM}};
  frontEndRegMap_16 = _RAND_103[5:0];
  _RAND_104 = {1{`RANDOM}};
  frontEndRegMap_15 = _RAND_104[5:0];
  _RAND_105 = {1{`RANDOM}};
  frontEndRegMap_14 = _RAND_105[5:0];
  _RAND_106 = {1{`RANDOM}};
  frontEndRegMap_13 = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  frontEndRegMap_12 = _RAND_107[5:0];
  _RAND_108 = {1{`RANDOM}};
  frontEndRegMap_11 = _RAND_108[5:0];
  _RAND_109 = {1{`RANDOM}};
  frontEndRegMap_10 = _RAND_109[5:0];
  _RAND_110 = {1{`RANDOM}};
  frontEndRegMap_9 = _RAND_110[5:0];
  _RAND_111 = {1{`RANDOM}};
  frontEndRegMap_8 = _RAND_111[5:0];
  _RAND_112 = {1{`RANDOM}};
  frontEndRegMap_7 = _RAND_112[5:0];
  _RAND_113 = {1{`RANDOM}};
  frontEndRegMap_6 = _RAND_113[5:0];
  _RAND_114 = {1{`RANDOM}};
  frontEndRegMap_5 = _RAND_114[5:0];
  _RAND_115 = {1{`RANDOM}};
  frontEndRegMap_4 = _RAND_115[5:0];
  _RAND_116 = {1{`RANDOM}};
  frontEndRegMap_3 = _RAND_116[5:0];
  _RAND_117 = {1{`RANDOM}};
  frontEndRegMap_2 = _RAND_117[5:0];
  _RAND_118 = {1{`RANDOM}};
  frontEndRegMap_1 = _RAND_118[5:0];
  _RAND_119 = {1{`RANDOM}};
  frontEndRegMap_0 = _RAND_119[5:0];
  _RAND_120 = {1{`RANDOM}};
  PRFFreeList_0 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  PRFFreeList_1 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  PRFFreeList_2 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  PRFFreeList_3 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  PRFFreeList_4 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  PRFFreeList_5 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  PRFFreeList_6 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  PRFFreeList_7 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  PRFFreeList_8 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  PRFFreeList_9 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  PRFFreeList_10 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  PRFFreeList_11 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  PRFFreeList_12 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  PRFFreeList_13 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  PRFFreeList_14 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  PRFFreeList_15 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  PRFFreeList_16 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  PRFFreeList_17 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  PRFFreeList_18 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  PRFFreeList_19 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  PRFFreeList_20 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  PRFFreeList_21 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  PRFFreeList_22 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  PRFFreeList_23 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  PRFFreeList_24 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  PRFFreeList_25 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  PRFFreeList_26 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  PRFFreeList_27 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  PRFFreeList_28 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  PRFFreeList_29 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  PRFFreeList_30 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  PRFFreeList_31 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  PRFFreeList_32 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  PRFFreeList_33 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  PRFFreeList_34 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  PRFFreeList_35 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  PRFFreeList_36 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  PRFFreeList_37 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  PRFFreeList_38 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  PRFFreeList_39 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  PRFFreeList_40 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  PRFFreeList_41 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  PRFFreeList_42 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  PRFFreeList_43 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  PRFFreeList_44 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  PRFFreeList_45 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  PRFFreeList_46 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  PRFFreeList_47 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  PRFFreeList_48 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  PRFFreeList_49 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  PRFFreeList_50 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  PRFFreeList_51 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  PRFFreeList_52 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  PRFFreeList_53 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  PRFFreeList_54 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  PRFFreeList_55 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  PRFFreeList_56 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  PRFFreeList_57 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  PRFFreeList_58 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  PRFFreeList_59 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  PRFFreeList_60 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  PRFFreeList_61 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  PRFFreeList_62 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  branchPCMask = _RAND_183[4:0];
  _RAND_184 = {1{`RANDOM}};
  branchReg = _RAND_184[0:0];
  _RAND_185 = {2{`RANDOM}};
  csrReadDataReg = _RAND_185[63:0];
  _RAND_186 = {1{`RANDOM}};
  csrAddrReg = _RAND_186[11:0];
  _RAND_187 = {2{`RANDOM}};
  csrImmReg = _RAND_187[63:0];
  _RAND_188 = {1{`RANDOM}};
  architecturalRegMap_0 = _RAND_188[5:0];
  _RAND_189 = {1{`RANDOM}};
  architecturalRegMap_1 = _RAND_189[5:0];
  _RAND_190 = {1{`RANDOM}};
  architecturalRegMap_2 = _RAND_190[5:0];
  _RAND_191 = {1{`RANDOM}};
  architecturalRegMap_3 = _RAND_191[5:0];
  _RAND_192 = {1{`RANDOM}};
  architecturalRegMap_4 = _RAND_192[5:0];
  _RAND_193 = {1{`RANDOM}};
  architecturalRegMap_5 = _RAND_193[5:0];
  _RAND_194 = {1{`RANDOM}};
  architecturalRegMap_6 = _RAND_194[5:0];
  _RAND_195 = {1{`RANDOM}};
  architecturalRegMap_7 = _RAND_195[5:0];
  _RAND_196 = {1{`RANDOM}};
  architecturalRegMap_8 = _RAND_196[5:0];
  _RAND_197 = {1{`RANDOM}};
  architecturalRegMap_9 = _RAND_197[5:0];
  _RAND_198 = {1{`RANDOM}};
  architecturalRegMap_10 = _RAND_198[5:0];
  _RAND_199 = {1{`RANDOM}};
  architecturalRegMap_11 = _RAND_199[5:0];
  _RAND_200 = {1{`RANDOM}};
  architecturalRegMap_12 = _RAND_200[5:0];
  _RAND_201 = {1{`RANDOM}};
  architecturalRegMap_13 = _RAND_201[5:0];
  _RAND_202 = {1{`RANDOM}};
  architecturalRegMap_14 = _RAND_202[5:0];
  _RAND_203 = {1{`RANDOM}};
  architecturalRegMap_15 = _RAND_203[5:0];
  _RAND_204 = {1{`RANDOM}};
  architecturalRegMap_16 = _RAND_204[5:0];
  _RAND_205 = {1{`RANDOM}};
  architecturalRegMap_17 = _RAND_205[5:0];
  _RAND_206 = {1{`RANDOM}};
  architecturalRegMap_18 = _RAND_206[5:0];
  _RAND_207 = {1{`RANDOM}};
  architecturalRegMap_19 = _RAND_207[5:0];
  _RAND_208 = {1{`RANDOM}};
  architecturalRegMap_20 = _RAND_208[5:0];
  _RAND_209 = {1{`RANDOM}};
  architecturalRegMap_21 = _RAND_209[5:0];
  _RAND_210 = {1{`RANDOM}};
  architecturalRegMap_22 = _RAND_210[5:0];
  _RAND_211 = {1{`RANDOM}};
  architecturalRegMap_23 = _RAND_211[5:0];
  _RAND_212 = {1{`RANDOM}};
  architecturalRegMap_24 = _RAND_212[5:0];
  _RAND_213 = {1{`RANDOM}};
  architecturalRegMap_25 = _RAND_213[5:0];
  _RAND_214 = {1{`RANDOM}};
  architecturalRegMap_26 = _RAND_214[5:0];
  _RAND_215 = {1{`RANDOM}};
  architecturalRegMap_27 = _RAND_215[5:0];
  _RAND_216 = {1{`RANDOM}};
  architecturalRegMap_28 = _RAND_216[5:0];
  _RAND_217 = {1{`RANDOM}};
  architecturalRegMap_29 = _RAND_217[5:0];
  _RAND_218 = {1{`RANDOM}};
  architecturalRegMap_30 = _RAND_218[5:0];
  _RAND_219 = {1{`RANDOM}};
  architecturalRegMap_31 = _RAND_219[5:0];
  _RAND_220 = {1{`RANDOM}};
  reservedRegMap1_0 = _RAND_220[5:0];
  _RAND_221 = {1{`RANDOM}};
  reservedRegMap1_1 = _RAND_221[5:0];
  _RAND_222 = {1{`RANDOM}};
  reservedRegMap1_2 = _RAND_222[5:0];
  _RAND_223 = {1{`RANDOM}};
  reservedRegMap1_3 = _RAND_223[5:0];
  _RAND_224 = {1{`RANDOM}};
  reservedRegMap1_4 = _RAND_224[5:0];
  _RAND_225 = {1{`RANDOM}};
  reservedRegMap1_5 = _RAND_225[5:0];
  _RAND_226 = {1{`RANDOM}};
  reservedRegMap1_6 = _RAND_226[5:0];
  _RAND_227 = {1{`RANDOM}};
  reservedRegMap1_7 = _RAND_227[5:0];
  _RAND_228 = {1{`RANDOM}};
  reservedRegMap1_8 = _RAND_228[5:0];
  _RAND_229 = {1{`RANDOM}};
  reservedRegMap1_9 = _RAND_229[5:0];
  _RAND_230 = {1{`RANDOM}};
  reservedRegMap1_10 = _RAND_230[5:0];
  _RAND_231 = {1{`RANDOM}};
  reservedRegMap1_11 = _RAND_231[5:0];
  _RAND_232 = {1{`RANDOM}};
  reservedRegMap1_12 = _RAND_232[5:0];
  _RAND_233 = {1{`RANDOM}};
  reservedRegMap1_13 = _RAND_233[5:0];
  _RAND_234 = {1{`RANDOM}};
  reservedRegMap1_14 = _RAND_234[5:0];
  _RAND_235 = {1{`RANDOM}};
  reservedRegMap1_15 = _RAND_235[5:0];
  _RAND_236 = {1{`RANDOM}};
  reservedRegMap1_16 = _RAND_236[5:0];
  _RAND_237 = {1{`RANDOM}};
  reservedRegMap1_17 = _RAND_237[5:0];
  _RAND_238 = {1{`RANDOM}};
  reservedRegMap1_18 = _RAND_238[5:0];
  _RAND_239 = {1{`RANDOM}};
  reservedRegMap1_19 = _RAND_239[5:0];
  _RAND_240 = {1{`RANDOM}};
  reservedRegMap1_20 = _RAND_240[5:0];
  _RAND_241 = {1{`RANDOM}};
  reservedRegMap1_21 = _RAND_241[5:0];
  _RAND_242 = {1{`RANDOM}};
  reservedRegMap1_22 = _RAND_242[5:0];
  _RAND_243 = {1{`RANDOM}};
  reservedRegMap1_23 = _RAND_243[5:0];
  _RAND_244 = {1{`RANDOM}};
  reservedRegMap1_24 = _RAND_244[5:0];
  _RAND_245 = {1{`RANDOM}};
  reservedRegMap1_25 = _RAND_245[5:0];
  _RAND_246 = {1{`RANDOM}};
  reservedRegMap1_26 = _RAND_246[5:0];
  _RAND_247 = {1{`RANDOM}};
  reservedRegMap1_27 = _RAND_247[5:0];
  _RAND_248 = {1{`RANDOM}};
  reservedRegMap1_28 = _RAND_248[5:0];
  _RAND_249 = {1{`RANDOM}};
  reservedRegMap1_29 = _RAND_249[5:0];
  _RAND_250 = {1{`RANDOM}};
  reservedRegMap1_30 = _RAND_250[5:0];
  _RAND_251 = {1{`RANDOM}};
  reservedRegMap1_31 = _RAND_251[5:0];
  _RAND_252 = {1{`RANDOM}};
  reservedRegMap2_0 = _RAND_252[5:0];
  _RAND_253 = {1{`RANDOM}};
  reservedRegMap2_1 = _RAND_253[5:0];
  _RAND_254 = {1{`RANDOM}};
  reservedRegMap2_2 = _RAND_254[5:0];
  _RAND_255 = {1{`RANDOM}};
  reservedRegMap2_3 = _RAND_255[5:0];
  _RAND_256 = {1{`RANDOM}};
  reservedRegMap2_4 = _RAND_256[5:0];
  _RAND_257 = {1{`RANDOM}};
  reservedRegMap2_5 = _RAND_257[5:0];
  _RAND_258 = {1{`RANDOM}};
  reservedRegMap2_6 = _RAND_258[5:0];
  _RAND_259 = {1{`RANDOM}};
  reservedRegMap2_7 = _RAND_259[5:0];
  _RAND_260 = {1{`RANDOM}};
  reservedRegMap2_8 = _RAND_260[5:0];
  _RAND_261 = {1{`RANDOM}};
  reservedRegMap2_9 = _RAND_261[5:0];
  _RAND_262 = {1{`RANDOM}};
  reservedRegMap2_10 = _RAND_262[5:0];
  _RAND_263 = {1{`RANDOM}};
  reservedRegMap2_11 = _RAND_263[5:0];
  _RAND_264 = {1{`RANDOM}};
  reservedRegMap2_12 = _RAND_264[5:0];
  _RAND_265 = {1{`RANDOM}};
  reservedRegMap2_13 = _RAND_265[5:0];
  _RAND_266 = {1{`RANDOM}};
  reservedRegMap2_14 = _RAND_266[5:0];
  _RAND_267 = {1{`RANDOM}};
  reservedRegMap2_15 = _RAND_267[5:0];
  _RAND_268 = {1{`RANDOM}};
  reservedRegMap2_16 = _RAND_268[5:0];
  _RAND_269 = {1{`RANDOM}};
  reservedRegMap2_17 = _RAND_269[5:0];
  _RAND_270 = {1{`RANDOM}};
  reservedRegMap2_18 = _RAND_270[5:0];
  _RAND_271 = {1{`RANDOM}};
  reservedRegMap2_19 = _RAND_271[5:0];
  _RAND_272 = {1{`RANDOM}};
  reservedRegMap2_20 = _RAND_272[5:0];
  _RAND_273 = {1{`RANDOM}};
  reservedRegMap2_21 = _RAND_273[5:0];
  _RAND_274 = {1{`RANDOM}};
  reservedRegMap2_22 = _RAND_274[5:0];
  _RAND_275 = {1{`RANDOM}};
  reservedRegMap2_23 = _RAND_275[5:0];
  _RAND_276 = {1{`RANDOM}};
  reservedRegMap2_24 = _RAND_276[5:0];
  _RAND_277 = {1{`RANDOM}};
  reservedRegMap2_25 = _RAND_277[5:0];
  _RAND_278 = {1{`RANDOM}};
  reservedRegMap2_26 = _RAND_278[5:0];
  _RAND_279 = {1{`RANDOM}};
  reservedRegMap2_27 = _RAND_279[5:0];
  _RAND_280 = {1{`RANDOM}};
  reservedRegMap2_28 = _RAND_280[5:0];
  _RAND_281 = {1{`RANDOM}};
  reservedRegMap2_29 = _RAND_281[5:0];
  _RAND_282 = {1{`RANDOM}};
  reservedRegMap2_30 = _RAND_282[5:0];
  _RAND_283 = {1{`RANDOM}};
  reservedRegMap2_31 = _RAND_283[5:0];
  _RAND_284 = {1{`RANDOM}};
  reservedRegMap3_0 = _RAND_284[5:0];
  _RAND_285 = {1{`RANDOM}};
  reservedRegMap3_1 = _RAND_285[5:0];
  _RAND_286 = {1{`RANDOM}};
  reservedRegMap3_2 = _RAND_286[5:0];
  _RAND_287 = {1{`RANDOM}};
  reservedRegMap3_3 = _RAND_287[5:0];
  _RAND_288 = {1{`RANDOM}};
  reservedRegMap3_4 = _RAND_288[5:0];
  _RAND_289 = {1{`RANDOM}};
  reservedRegMap3_5 = _RAND_289[5:0];
  _RAND_290 = {1{`RANDOM}};
  reservedRegMap3_6 = _RAND_290[5:0];
  _RAND_291 = {1{`RANDOM}};
  reservedRegMap3_7 = _RAND_291[5:0];
  _RAND_292 = {1{`RANDOM}};
  reservedRegMap3_8 = _RAND_292[5:0];
  _RAND_293 = {1{`RANDOM}};
  reservedRegMap3_9 = _RAND_293[5:0];
  _RAND_294 = {1{`RANDOM}};
  reservedRegMap3_10 = _RAND_294[5:0];
  _RAND_295 = {1{`RANDOM}};
  reservedRegMap3_11 = _RAND_295[5:0];
  _RAND_296 = {1{`RANDOM}};
  reservedRegMap3_12 = _RAND_296[5:0];
  _RAND_297 = {1{`RANDOM}};
  reservedRegMap3_13 = _RAND_297[5:0];
  _RAND_298 = {1{`RANDOM}};
  reservedRegMap3_14 = _RAND_298[5:0];
  _RAND_299 = {1{`RANDOM}};
  reservedRegMap3_15 = _RAND_299[5:0];
  _RAND_300 = {1{`RANDOM}};
  reservedRegMap3_16 = _RAND_300[5:0];
  _RAND_301 = {1{`RANDOM}};
  reservedRegMap3_17 = _RAND_301[5:0];
  _RAND_302 = {1{`RANDOM}};
  reservedRegMap3_18 = _RAND_302[5:0];
  _RAND_303 = {1{`RANDOM}};
  reservedRegMap3_19 = _RAND_303[5:0];
  _RAND_304 = {1{`RANDOM}};
  reservedRegMap3_20 = _RAND_304[5:0];
  _RAND_305 = {1{`RANDOM}};
  reservedRegMap3_21 = _RAND_305[5:0];
  _RAND_306 = {1{`RANDOM}};
  reservedRegMap3_22 = _RAND_306[5:0];
  _RAND_307 = {1{`RANDOM}};
  reservedRegMap3_23 = _RAND_307[5:0];
  _RAND_308 = {1{`RANDOM}};
  reservedRegMap3_24 = _RAND_308[5:0];
  _RAND_309 = {1{`RANDOM}};
  reservedRegMap3_25 = _RAND_309[5:0];
  _RAND_310 = {1{`RANDOM}};
  reservedRegMap3_26 = _RAND_310[5:0];
  _RAND_311 = {1{`RANDOM}};
  reservedRegMap3_27 = _RAND_311[5:0];
  _RAND_312 = {1{`RANDOM}};
  reservedRegMap3_28 = _RAND_312[5:0];
  _RAND_313 = {1{`RANDOM}};
  reservedRegMap3_29 = _RAND_313[5:0];
  _RAND_314 = {1{`RANDOM}};
  reservedRegMap3_30 = _RAND_314[5:0];
  _RAND_315 = {1{`RANDOM}};
  reservedRegMap3_31 = _RAND_315[5:0];
  _RAND_316 = {1{`RANDOM}};
  reservedRegMap4_0 = _RAND_316[5:0];
  _RAND_317 = {1{`RANDOM}};
  reservedRegMap4_1 = _RAND_317[5:0];
  _RAND_318 = {1{`RANDOM}};
  reservedRegMap4_2 = _RAND_318[5:0];
  _RAND_319 = {1{`RANDOM}};
  reservedRegMap4_3 = _RAND_319[5:0];
  _RAND_320 = {1{`RANDOM}};
  reservedRegMap4_4 = _RAND_320[5:0];
  _RAND_321 = {1{`RANDOM}};
  reservedRegMap4_5 = _RAND_321[5:0];
  _RAND_322 = {1{`RANDOM}};
  reservedRegMap4_6 = _RAND_322[5:0];
  _RAND_323 = {1{`RANDOM}};
  reservedRegMap4_7 = _RAND_323[5:0];
  _RAND_324 = {1{`RANDOM}};
  reservedRegMap4_8 = _RAND_324[5:0];
  _RAND_325 = {1{`RANDOM}};
  reservedRegMap4_9 = _RAND_325[5:0];
  _RAND_326 = {1{`RANDOM}};
  reservedRegMap4_10 = _RAND_326[5:0];
  _RAND_327 = {1{`RANDOM}};
  reservedRegMap4_11 = _RAND_327[5:0];
  _RAND_328 = {1{`RANDOM}};
  reservedRegMap4_12 = _RAND_328[5:0];
  _RAND_329 = {1{`RANDOM}};
  reservedRegMap4_13 = _RAND_329[5:0];
  _RAND_330 = {1{`RANDOM}};
  reservedRegMap4_14 = _RAND_330[5:0];
  _RAND_331 = {1{`RANDOM}};
  reservedRegMap4_15 = _RAND_331[5:0];
  _RAND_332 = {1{`RANDOM}};
  reservedRegMap4_16 = _RAND_332[5:0];
  _RAND_333 = {1{`RANDOM}};
  reservedRegMap4_17 = _RAND_333[5:0];
  _RAND_334 = {1{`RANDOM}};
  reservedRegMap4_18 = _RAND_334[5:0];
  _RAND_335 = {1{`RANDOM}};
  reservedRegMap4_19 = _RAND_335[5:0];
  _RAND_336 = {1{`RANDOM}};
  reservedRegMap4_20 = _RAND_336[5:0];
  _RAND_337 = {1{`RANDOM}};
  reservedRegMap4_21 = _RAND_337[5:0];
  _RAND_338 = {1{`RANDOM}};
  reservedRegMap4_22 = _RAND_338[5:0];
  _RAND_339 = {1{`RANDOM}};
  reservedRegMap4_23 = _RAND_339[5:0];
  _RAND_340 = {1{`RANDOM}};
  reservedRegMap4_24 = _RAND_340[5:0];
  _RAND_341 = {1{`RANDOM}};
  reservedRegMap4_25 = _RAND_341[5:0];
  _RAND_342 = {1{`RANDOM}};
  reservedRegMap4_26 = _RAND_342[5:0];
  _RAND_343 = {1{`RANDOM}};
  reservedRegMap4_27 = _RAND_343[5:0];
  _RAND_344 = {1{`RANDOM}};
  reservedRegMap4_28 = _RAND_344[5:0];
  _RAND_345 = {1{`RANDOM}};
  reservedRegMap4_29 = _RAND_345[5:0];
  _RAND_346 = {1{`RANDOM}};
  reservedRegMap4_30 = _RAND_346[5:0];
  _RAND_347 = {1{`RANDOM}};
  reservedRegMap4_31 = _RAND_347[5:0];
  _RAND_348 = {1{`RANDOM}};
  reservedFreeList1_0 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  reservedFreeList1_1 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  reservedFreeList1_2 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  reservedFreeList1_3 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  reservedFreeList1_4 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  reservedFreeList1_5 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  reservedFreeList1_6 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  reservedFreeList1_7 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  reservedFreeList1_8 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  reservedFreeList1_9 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  reservedFreeList1_10 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  reservedFreeList1_11 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  reservedFreeList1_12 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  reservedFreeList1_13 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  reservedFreeList1_14 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  reservedFreeList1_15 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  reservedFreeList1_16 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  reservedFreeList1_17 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  reservedFreeList1_18 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  reservedFreeList1_19 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  reservedFreeList1_20 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  reservedFreeList1_21 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  reservedFreeList1_22 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  reservedFreeList1_23 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  reservedFreeList1_24 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  reservedFreeList1_25 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  reservedFreeList1_26 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  reservedFreeList1_27 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  reservedFreeList1_28 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  reservedFreeList1_29 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  reservedFreeList1_30 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  reservedFreeList1_31 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  reservedFreeList1_32 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  reservedFreeList1_33 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  reservedFreeList1_34 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  reservedFreeList1_35 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  reservedFreeList1_36 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  reservedFreeList1_37 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  reservedFreeList1_38 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  reservedFreeList1_39 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  reservedFreeList1_40 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  reservedFreeList1_41 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  reservedFreeList1_42 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  reservedFreeList1_43 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  reservedFreeList1_44 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  reservedFreeList1_45 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  reservedFreeList1_46 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  reservedFreeList1_47 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  reservedFreeList1_48 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  reservedFreeList1_49 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  reservedFreeList1_50 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  reservedFreeList1_51 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  reservedFreeList1_52 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  reservedFreeList1_53 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  reservedFreeList1_54 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  reservedFreeList1_55 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  reservedFreeList1_56 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  reservedFreeList1_57 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  reservedFreeList1_58 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  reservedFreeList1_59 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  reservedFreeList1_60 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  reservedFreeList1_61 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  reservedFreeList1_62 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  reservedFreeList2_0 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  reservedFreeList2_1 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  reservedFreeList2_2 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  reservedFreeList2_3 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  reservedFreeList2_4 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  reservedFreeList2_5 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  reservedFreeList2_6 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  reservedFreeList2_7 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  reservedFreeList2_8 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  reservedFreeList2_9 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  reservedFreeList2_10 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  reservedFreeList2_11 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  reservedFreeList2_12 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  reservedFreeList2_13 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  reservedFreeList2_14 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  reservedFreeList2_15 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  reservedFreeList2_16 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  reservedFreeList2_17 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  reservedFreeList2_18 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  reservedFreeList2_19 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  reservedFreeList2_20 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  reservedFreeList2_21 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  reservedFreeList2_22 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  reservedFreeList2_23 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  reservedFreeList2_24 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  reservedFreeList2_25 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  reservedFreeList2_26 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  reservedFreeList2_27 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  reservedFreeList2_28 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  reservedFreeList2_29 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  reservedFreeList2_30 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  reservedFreeList2_31 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  reservedFreeList2_32 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  reservedFreeList2_33 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  reservedFreeList2_34 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  reservedFreeList2_35 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  reservedFreeList2_36 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  reservedFreeList2_37 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  reservedFreeList2_38 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  reservedFreeList2_39 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  reservedFreeList2_40 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  reservedFreeList2_41 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  reservedFreeList2_42 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  reservedFreeList2_43 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  reservedFreeList2_44 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  reservedFreeList2_45 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  reservedFreeList2_46 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  reservedFreeList2_47 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  reservedFreeList2_48 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  reservedFreeList2_49 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  reservedFreeList2_50 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  reservedFreeList2_51 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  reservedFreeList2_52 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  reservedFreeList2_53 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  reservedFreeList2_54 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  reservedFreeList2_55 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  reservedFreeList2_56 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  reservedFreeList2_57 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  reservedFreeList2_58 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  reservedFreeList2_59 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  reservedFreeList2_60 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  reservedFreeList2_61 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  reservedFreeList2_62 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  reservedFreeList3_0 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  reservedFreeList3_1 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  reservedFreeList3_2 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  reservedFreeList3_3 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  reservedFreeList3_4 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  reservedFreeList3_5 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  reservedFreeList3_6 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  reservedFreeList3_7 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  reservedFreeList3_8 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  reservedFreeList3_9 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  reservedFreeList3_10 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  reservedFreeList3_11 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  reservedFreeList3_12 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  reservedFreeList3_13 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  reservedFreeList3_14 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  reservedFreeList3_15 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  reservedFreeList3_16 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  reservedFreeList3_17 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  reservedFreeList3_18 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  reservedFreeList3_19 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  reservedFreeList3_20 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  reservedFreeList3_21 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  reservedFreeList3_22 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  reservedFreeList3_23 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  reservedFreeList3_24 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  reservedFreeList3_25 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  reservedFreeList3_26 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  reservedFreeList3_27 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  reservedFreeList3_28 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  reservedFreeList3_29 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  reservedFreeList3_30 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  reservedFreeList3_31 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  reservedFreeList3_32 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  reservedFreeList3_33 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  reservedFreeList3_34 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  reservedFreeList3_35 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  reservedFreeList3_36 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  reservedFreeList3_37 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  reservedFreeList3_38 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  reservedFreeList3_39 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  reservedFreeList3_40 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  reservedFreeList3_41 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  reservedFreeList3_42 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  reservedFreeList3_43 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  reservedFreeList3_44 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  reservedFreeList3_45 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  reservedFreeList3_46 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  reservedFreeList3_47 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  reservedFreeList3_48 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  reservedFreeList3_49 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  reservedFreeList3_50 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  reservedFreeList3_51 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  reservedFreeList3_52 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  reservedFreeList3_53 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  reservedFreeList3_54 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  reservedFreeList3_55 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  reservedFreeList3_56 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  reservedFreeList3_57 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  reservedFreeList3_58 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  reservedFreeList3_59 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  reservedFreeList3_60 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  reservedFreeList3_61 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  reservedFreeList3_62 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  reservedFreeList4_0 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  reservedFreeList4_1 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  reservedFreeList4_2 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  reservedFreeList4_3 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  reservedFreeList4_4 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  reservedFreeList4_5 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  reservedFreeList4_6 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  reservedFreeList4_7 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  reservedFreeList4_8 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  reservedFreeList4_9 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  reservedFreeList4_10 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  reservedFreeList4_11 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  reservedFreeList4_12 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  reservedFreeList4_13 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  reservedFreeList4_14 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  reservedFreeList4_15 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  reservedFreeList4_16 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  reservedFreeList4_17 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  reservedFreeList4_18 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  reservedFreeList4_19 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  reservedFreeList4_20 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  reservedFreeList4_21 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  reservedFreeList4_22 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  reservedFreeList4_23 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  reservedFreeList4_24 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  reservedFreeList4_25 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  reservedFreeList4_26 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  reservedFreeList4_27 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  reservedFreeList4_28 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  reservedFreeList4_29 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  reservedFreeList4_30 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  reservedFreeList4_31 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  reservedFreeList4_32 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  reservedFreeList4_33 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  reservedFreeList4_34 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  reservedFreeList4_35 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  reservedFreeList4_36 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  reservedFreeList4_37 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  reservedFreeList4_38 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  reservedFreeList4_39 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  reservedFreeList4_40 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  reservedFreeList4_41 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  reservedFreeList4_42 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  reservedFreeList4_43 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  reservedFreeList4_44 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  reservedFreeList4_45 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  reservedFreeList4_46 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  reservedFreeList4_47 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  reservedFreeList4_48 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  reservedFreeList4_49 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  reservedFreeList4_50 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  reservedFreeList4_51 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  reservedFreeList4_52 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  reservedFreeList4_53 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  reservedFreeList4_54 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  reservedFreeList4_55 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  reservedFreeList4_56 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  reservedFreeList4_57 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  reservedFreeList4_58 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  reservedFreeList4_59 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  reservedFreeList4_60 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  reservedFreeList4_61 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  reservedFreeList4_62 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  reservedValidList1_0 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  reservedValidList1_1 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  reservedValidList1_2 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  reservedValidList1_3 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  reservedValidList1_4 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  reservedValidList1_5 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  reservedValidList1_6 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  reservedValidList1_7 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  reservedValidList1_8 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  reservedValidList1_9 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  reservedValidList1_10 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  reservedValidList1_11 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  reservedValidList1_12 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  reservedValidList1_13 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  reservedValidList1_14 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  reservedValidList1_15 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  reservedValidList1_16 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  reservedValidList1_17 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  reservedValidList1_18 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  reservedValidList1_19 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  reservedValidList1_20 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  reservedValidList1_21 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  reservedValidList1_22 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  reservedValidList1_23 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  reservedValidList1_24 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  reservedValidList1_25 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  reservedValidList1_26 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  reservedValidList1_27 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  reservedValidList1_28 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  reservedValidList1_29 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  reservedValidList1_30 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  reservedValidList1_31 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  reservedValidList1_32 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  reservedValidList1_33 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  reservedValidList1_34 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  reservedValidList1_35 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  reservedValidList1_36 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  reservedValidList1_37 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  reservedValidList1_38 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  reservedValidList1_39 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  reservedValidList1_40 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  reservedValidList1_41 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  reservedValidList1_42 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  reservedValidList1_43 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  reservedValidList1_44 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  reservedValidList1_45 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  reservedValidList1_46 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  reservedValidList1_47 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  reservedValidList1_48 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  reservedValidList1_49 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  reservedValidList1_50 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  reservedValidList1_51 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  reservedValidList1_52 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  reservedValidList1_53 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  reservedValidList1_54 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  reservedValidList1_55 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  reservedValidList1_56 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  reservedValidList1_57 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  reservedValidList1_58 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  reservedValidList1_59 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  reservedValidList1_60 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  reservedValidList1_61 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  reservedValidList1_62 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  reservedValidList1_63 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  reservedValidList2_0 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  reservedValidList2_1 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  reservedValidList2_2 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  reservedValidList2_3 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  reservedValidList2_4 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  reservedValidList2_5 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  reservedValidList2_6 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  reservedValidList2_7 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  reservedValidList2_8 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  reservedValidList2_9 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  reservedValidList2_10 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  reservedValidList2_11 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  reservedValidList2_12 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  reservedValidList2_13 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  reservedValidList2_14 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  reservedValidList2_15 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  reservedValidList2_16 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  reservedValidList2_17 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  reservedValidList2_18 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  reservedValidList2_19 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  reservedValidList2_20 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  reservedValidList2_21 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  reservedValidList2_22 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  reservedValidList2_23 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  reservedValidList2_24 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  reservedValidList2_25 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  reservedValidList2_26 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  reservedValidList2_27 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  reservedValidList2_28 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  reservedValidList2_29 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  reservedValidList2_30 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  reservedValidList2_31 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  reservedValidList2_32 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  reservedValidList2_33 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  reservedValidList2_34 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  reservedValidList2_35 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  reservedValidList2_36 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  reservedValidList2_37 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  reservedValidList2_38 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  reservedValidList2_39 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  reservedValidList2_40 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  reservedValidList2_41 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  reservedValidList2_42 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  reservedValidList2_43 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  reservedValidList2_44 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  reservedValidList2_45 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  reservedValidList2_46 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  reservedValidList2_47 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  reservedValidList2_48 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  reservedValidList2_49 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  reservedValidList2_50 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  reservedValidList2_51 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  reservedValidList2_52 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  reservedValidList2_53 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  reservedValidList2_54 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  reservedValidList2_55 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  reservedValidList2_56 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  reservedValidList2_57 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  reservedValidList2_58 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  reservedValidList2_59 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  reservedValidList2_60 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  reservedValidList2_61 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  reservedValidList2_62 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  reservedValidList2_63 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  reservedValidList3_0 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  reservedValidList3_1 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  reservedValidList3_2 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  reservedValidList3_3 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  reservedValidList3_4 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  reservedValidList3_5 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  reservedValidList3_6 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  reservedValidList3_7 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  reservedValidList3_8 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  reservedValidList3_9 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  reservedValidList3_10 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  reservedValidList3_11 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  reservedValidList3_12 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  reservedValidList3_13 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  reservedValidList3_14 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  reservedValidList3_15 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  reservedValidList3_16 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  reservedValidList3_17 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  reservedValidList3_18 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  reservedValidList3_19 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  reservedValidList3_20 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  reservedValidList3_21 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  reservedValidList3_22 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  reservedValidList3_23 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  reservedValidList3_24 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  reservedValidList3_25 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  reservedValidList3_26 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  reservedValidList3_27 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  reservedValidList3_28 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  reservedValidList3_29 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  reservedValidList3_30 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  reservedValidList3_31 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  reservedValidList3_32 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  reservedValidList3_33 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  reservedValidList3_34 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  reservedValidList3_35 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  reservedValidList3_36 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  reservedValidList3_37 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  reservedValidList3_38 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  reservedValidList3_39 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  reservedValidList3_40 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  reservedValidList3_41 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  reservedValidList3_42 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  reservedValidList3_43 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  reservedValidList3_44 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  reservedValidList3_45 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  reservedValidList3_46 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  reservedValidList3_47 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  reservedValidList3_48 = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  reservedValidList3_49 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  reservedValidList3_50 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  reservedValidList3_51 = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  reservedValidList3_52 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  reservedValidList3_53 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  reservedValidList3_54 = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  reservedValidList3_55 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  reservedValidList3_56 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  reservedValidList3_57 = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  reservedValidList3_58 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  reservedValidList3_59 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  reservedValidList3_60 = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  reservedValidList3_61 = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  reservedValidList3_62 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  reservedValidList3_63 = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  reservedValidList4_0 = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  reservedValidList4_1 = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  reservedValidList4_2 = _RAND_794[0:0];
  _RAND_795 = {1{`RANDOM}};
  reservedValidList4_3 = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  reservedValidList4_4 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  reservedValidList4_5 = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  reservedValidList4_6 = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  reservedValidList4_7 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  reservedValidList4_8 = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  reservedValidList4_9 = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  reservedValidList4_10 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  reservedValidList4_11 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  reservedValidList4_12 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  reservedValidList4_13 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  reservedValidList4_14 = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  reservedValidList4_15 = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  reservedValidList4_16 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  reservedValidList4_17 = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  reservedValidList4_18 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  reservedValidList4_19 = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  reservedValidList4_20 = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  reservedValidList4_21 = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  reservedValidList4_22 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  reservedValidList4_23 = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  reservedValidList4_24 = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  reservedValidList4_25 = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  reservedValidList4_26 = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  reservedValidList4_27 = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  reservedValidList4_28 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  reservedValidList4_29 = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  reservedValidList4_30 = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  reservedValidList4_31 = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  reservedValidList4_32 = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  reservedValidList4_33 = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  reservedValidList4_34 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  reservedValidList4_35 = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  reservedValidList4_36 = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  reservedValidList4_37 = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  reservedValidList4_38 = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  reservedValidList4_39 = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  reservedValidList4_40 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  reservedValidList4_41 = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  reservedValidList4_42 = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  reservedValidList4_43 = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  reservedValidList4_44 = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  reservedValidList4_45 = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  reservedValidList4_46 = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  reservedValidList4_47 = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  reservedValidList4_48 = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  reservedValidList4_49 = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  reservedValidList4_50 = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  reservedValidList4_51 = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  reservedValidList4_52 = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  reservedValidList4_53 = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  reservedValidList4_54 = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  reservedValidList4_55 = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  reservedValidList4_56 = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  reservedValidList4_57 = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  reservedValidList4_58 = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  reservedValidList4_59 = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  reservedValidList4_60 = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  reservedValidList4_61 = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  reservedValidList4_62 = _RAND_854[0:0];
  _RAND_855 = {1{`RANDOM}};
  reservedValidList4_63 = _RAND_855[0:0];
  _RAND_856 = {2{`RANDOM}};
  ustatus = _RAND_856[63:0];
  _RAND_857 = {2{`RANDOM}};
  utvec = _RAND_857[63:0];
  _RAND_858 = {2{`RANDOM}};
  uepc = _RAND_858[63:0];
  _RAND_859 = {2{`RANDOM}};
  ucause = _RAND_859[63:0];
  _RAND_860 = {2{`RANDOM}};
  scounteren = _RAND_860[63:0];
  _RAND_861 = {2{`RANDOM}};
  satp = _RAND_861[63:0];
  _RAND_862 = {2{`RANDOM}};
  mstatus = _RAND_862[63:0];
  _RAND_863 = {2{`RANDOM}};
  misa = _RAND_863[63:0];
  _RAND_864 = {2{`RANDOM}};
  medeleg = _RAND_864[63:0];
  _RAND_865 = {2{`RANDOM}};
  mideleg = _RAND_865[63:0];
  _RAND_866 = {2{`RANDOM}};
  mie = _RAND_866[63:0];
  _RAND_867 = {2{`RANDOM}};
  mtvec = _RAND_867[63:0];
  _RAND_868 = {2{`RANDOM}};
  mcounteren = _RAND_868[63:0];
  _RAND_869 = {2{`RANDOM}};
  mscratch = _RAND_869[63:0];
  _RAND_870 = {2{`RANDOM}};
  mepc = _RAND_870[63:0];
  _RAND_871 = {2{`RANDOM}};
  mcause = _RAND_871[63:0];
  _RAND_872 = {2{`RANDOM}};
  mtval = _RAND_872[63:0];
  _RAND_873 = {2{`RANDOM}};
  mip = _RAND_873[63:0];
  _RAND_874 = {2{`RANDOM}};
  pmpcfg0 = _RAND_874[63:0];
  _RAND_875 = {2{`RANDOM}};
  pmpaddr0 = _RAND_875[63:0];
  _RAND_876 = {2{`RANDOM}};
  mvendorid = _RAND_876[63:0];
  _RAND_877 = {2{`RANDOM}};
  marchid = _RAND_877[63:0];
  _RAND_878 = {2{`RANDOM}};
  mimpid = _RAND_878[63:0];
  _RAND_879 = {2{`RANDOM}};
  mhartid = _RAND_879[63:0];
  _RAND_880 = {2{`RANDOM}};
  currentPrivilege = _RAND_880[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module storeDataIssue_Anon(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [10:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [10:0] io_deq_bits,
  input  [3:0]  modifyVal,
  input         modify,
  output [3:0]  allocatedAddr
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [10:0] memReg [0:15]; // @[storeDataIssue.scala 31:19]
  wire  memReg_io_deq_bits_MPORT_en; // @[storeDataIssue.scala 31:19]
  wire [3:0] memReg_io_deq_bits_MPORT_addr; // @[storeDataIssue.scala 31:19]
  wire [10:0] memReg_io_deq_bits_MPORT_data; // @[storeDataIssue.scala 31:19]
  wire [10:0] memReg_MPORT_data; // @[storeDataIssue.scala 31:19]
  wire [3:0] memReg_MPORT_addr; // @[storeDataIssue.scala 31:19]
  wire  memReg_MPORT_mask; // @[storeDataIssue.scala 31:19]
  wire  memReg_MPORT_en; // @[storeDataIssue.scala 31:19]
  wire [10:0] memReg_MPORT_1_data; // @[storeDataIssue.scala 31:19]
  wire [3:0] memReg_MPORT_1_addr; // @[storeDataIssue.scala 31:19]
  wire  memReg_MPORT_1_mask; // @[storeDataIssue.scala 31:19]
  wire  memReg_MPORT_1_en; // @[storeDataIssue.scala 31:19]
  reg [3:0] readPtr; // @[storeDataIssue.scala 25:24]
  wire [3:0] _nextRead_T_2 = readPtr + 4'h1; // @[storeDataIssue.scala 26:62]
  wire [3:0] nextRead = readPtr == 4'hf ? 4'h0 : _nextRead_T_2; // @[storeDataIssue.scala 26:21]
  reg [3:0] writePtr; // @[storeDataIssue.scala 27:25]
  wire [3:0] _nextWrite_T_2 = writePtr + 4'h1; // @[storeDataIssue.scala 28:65]
  wire [3:0] nextWrite = writePtr == 4'hf ? 4'h0 : _nextWrite_T_2; // @[storeDataIssue.scala 28:22]
  reg  emptyReg; // @[storeDataIssue.scala 34:25]
  reg  fullReg; // @[storeDataIssue.scala 35:24]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[storeDataIssue.scala 64:21]
  wire  _T_3 = io_deq_ready & io_deq_valid & io_enq_valid; // @[storeDataIssue.scala 64:37]
  wire  _T_4 = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready; // @[storeDataIssue.scala 64:53]
  wire  _T_5 = io_enq_valid & io_enq_ready; // @[storeDataIssue.scala 70:27]
  wire  _GEN_110 = io_enq_valid & io_enq_ready ? 1'h0 : _T_2; // @[storeDataIssue.scala 70:44]
  wire  incrRead = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready | _GEN_110; // @[storeDataIssue.scala 64:70 69:14]
  wire  incrWrite = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready | _T_5; // @[storeDataIssue.scala 64:70 68:15]
  wire  _GEN_3 = modify & ~emptyReg ? modifyVal == readPtr : emptyReg; // @[storeDataIssue.scala 53:29 58:14 34:25]
  wire  _GEN_69 = _T_2 ? nextRead == writePtr : _GEN_3; // @[storeDataIssue.scala 76:44 78:14]
  wire  _GEN_108 = io_enq_valid & io_enq_ready ? 1'h0 : _GEN_69; // @[storeDataIssue.scala 70:44 73:14]
  wire  _GEN_139 = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready ? _GEN_3 : _GEN_108; // @[storeDataIssue.scala 64:70]
  assign memReg_io_deq_bits_MPORT_en = 1'h1;
  assign memReg_io_deq_bits_MPORT_addr = readPtr;
  assign memReg_io_deq_bits_MPORT_data = memReg[memReg_io_deq_bits_MPORT_addr]; // @[storeDataIssue.scala 31:19]
  assign memReg_MPORT_data = io_enq_bits;
  assign memReg_MPORT_addr = writePtr;
  assign memReg_MPORT_mask = 1'h1;
  assign memReg_MPORT_en = _T_3 & io_enq_ready;
  assign memReg_MPORT_1_data = io_enq_bits;
  assign memReg_MPORT_1_addr = writePtr;
  assign memReg_MPORT_1_mask = 1'h1;
  assign memReg_MPORT_1_en = _T_4 ? 1'h0 : _T_5;
  assign io_enq_ready = (~fullReg | io_deq_valid & io_deq_ready) & ~modify; // @[storeDataIssue.scala 84:62]
  assign io_deq_valid = ~emptyReg; // @[storeDataIssue.scala 85:19]
  assign io_deq_bits = memReg_io_deq_bits_MPORT_data; // @[storeDataIssue.scala 83:15]
  assign allocatedAddr = writePtr; // @[storeDataIssue.scala 92:17]
  always @(posedge clock) begin
    if (memReg_MPORT_en & memReg_MPORT_mask) begin
      memReg[memReg_MPORT_addr] <= memReg_MPORT_data; // @[storeDataIssue.scala 31:19]
    end
    if (memReg_MPORT_1_en & memReg_MPORT_1_mask) begin
      memReg[memReg_MPORT_1_addr] <= memReg_MPORT_1_data; // @[storeDataIssue.scala 31:19]
    end
    if (reset) begin // @[storeDataIssue.scala 25:24]
      readPtr <= 4'h0; // @[storeDataIssue.scala 25:24]
    end else if (incrRead) begin // @[storeDataIssue.scala 48:19]
      if (readPtr == 4'hf) begin // @[storeDataIssue.scala 26:21]
        readPtr <= 4'h0;
      end else begin
        readPtr <= _nextRead_T_2;
      end
    end
    if (reset) begin // @[storeDataIssue.scala 27:25]
      writePtr <= 4'h0; // @[storeDataIssue.scala 27:25]
    end else if (modify & ~emptyReg) begin // @[storeDataIssue.scala 53:29]
      writePtr <= modifyVal; // @[storeDataIssue.scala 56:14]
    end else if (incrWrite) begin // @[storeDataIssue.scala 59:24]
      if (writePtr == 4'hf) begin // @[storeDataIssue.scala 28:22]
        writePtr <= 4'h0;
      end else begin
        writePtr <= _nextWrite_T_2;
      end
    end
    emptyReg <= reset | _GEN_139; // @[storeDataIssue.scala 34:{25,25}]
    if (reset) begin // @[storeDataIssue.scala 35:24]
      fullReg <= 1'h0; // @[storeDataIssue.scala 35:24]
    end else if (!(io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready)) begin // @[storeDataIssue.scala 64:70]
      if (io_enq_valid & io_enq_ready) begin // @[storeDataIssue.scala 70:44]
        fullReg <= nextWrite == readPtr; // @[storeDataIssue.scala 74:13]
      end else if (_T_2) begin // @[storeDataIssue.scala 76:44]
        fullReg <= 1'h0; // @[storeDataIssue.scala 77:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    memReg[initvar] = _RAND_0[10:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  readPtr = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  writePtr = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  emptyReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  fullReg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module storeDataIssue(
  input        clock,
  input        reset,
  input        fromROB_readyNow,
  input        fromBranch_passOrFail,
  input  [3:0] fromBranch_robAddr,
  input        fromBranch_valid,
  output       fromDecode_ready,
  input        fromDecode_valid,
  input  [5:0] fromDecode_rs2Addr,
  input  [4:0] fromDecode_branchMask,
  output       toPRF_valid,
  output [5:0] toPRF_rs2Addr,
  input        robMapUpdate_valid,
  input  [3:0] robMapUpdate_robAddr
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  wire  sdiFifo_clock; // @[storeDataIssue.scala 146:27]
  wire  sdiFifo_reset; // @[storeDataIssue.scala 146:27]
  wire  sdiFifo_io_enq_ready; // @[storeDataIssue.scala 146:27]
  wire  sdiFifo_io_enq_valid; // @[storeDataIssue.scala 146:27]
  wire [10:0] sdiFifo_io_enq_bits; // @[storeDataIssue.scala 146:27]
  wire  sdiFifo_io_deq_ready; // @[storeDataIssue.scala 146:27]
  wire  sdiFifo_io_deq_valid; // @[storeDataIssue.scala 146:27]
  wire [10:0] sdiFifo_io_deq_bits; // @[storeDataIssue.scala 146:27]
  wire [3:0] sdiFifo_modifyVal; // @[storeDataIssue.scala 146:27]
  wire  sdiFifo_modify; // @[storeDataIssue.scala 146:27]
  wire [3:0] sdiFifo_allocatedAddr; // @[storeDataIssue.scala 146:27]
  reg [3:0] map [0:15]; // @[storeDataIssue.scala 152:16]
  wire  map_sdiFifo_modifyVal_MPORT_en; // @[storeDataIssue.scala 152:16]
  wire [3:0] map_sdiFifo_modifyVal_MPORT_addr; // @[storeDataIssue.scala 152:16]
  wire [3:0] map_sdiFifo_modifyVal_MPORT_data; // @[storeDataIssue.scala 152:16]
  wire [3:0] map_MPORT_data; // @[storeDataIssue.scala 152:16]
  wire [3:0] map_MPORT_addr; // @[storeDataIssue.scala 152:16]
  wire  map_MPORT_mask; // @[storeDataIssue.scala 152:16]
  wire  map_MPORT_en; // @[storeDataIssue.scala 152:16]
  storeDataIssue_Anon sdiFifo ( // @[storeDataIssue.scala 146:27]
    .clock(sdiFifo_clock),
    .reset(sdiFifo_reset),
    .io_enq_ready(sdiFifo_io_enq_ready),
    .io_enq_valid(sdiFifo_io_enq_valid),
    .io_enq_bits(sdiFifo_io_enq_bits),
    .io_deq_ready(sdiFifo_io_deq_ready),
    .io_deq_valid(sdiFifo_io_deq_valid),
    .io_deq_bits(sdiFifo_io_deq_bits),
    .modifyVal(sdiFifo_modifyVal),
    .modify(sdiFifo_modify),
    .allocatedAddr(sdiFifo_allocatedAddr)
  );
  assign map_sdiFifo_modifyVal_MPORT_en = 1'h1;
  assign map_sdiFifo_modifyVal_MPORT_addr = fromBranch_robAddr;
  assign map_sdiFifo_modifyVal_MPORT_data = map[map_sdiFifo_modifyVal_MPORT_addr]; // @[storeDataIssue.scala 152:16]
  assign map_MPORT_data = sdiFifo_allocatedAddr;
  assign map_MPORT_addr = robMapUpdate_robAddr;
  assign map_MPORT_mask = 1'h1;
  assign map_MPORT_en = robMapUpdate_valid;
  assign fromDecode_ready = sdiFifo_io_enq_ready; // @[storeDataIssue.scala 167:29]
  assign toPRF_valid = sdiFifo_io_deq_valid; // @[storeDataIssue.scala 179:21]
  assign toPRF_rs2Addr = sdiFifo_io_deq_bits[5:0]; // @[storeDataIssue.scala 176:43]
  assign sdiFifo_clock = clock;
  assign sdiFifo_reset = reset;
  assign sdiFifo_io_enq_valid = fromDecode_valid; // @[storeDataIssue.scala 166:29]
  assign sdiFifo_io_enq_bits = {fromDecode_branchMask,fromDecode_rs2Addr}; // @[Cat.scala 33:92]
  assign sdiFifo_io_deq_ready = fromROB_readyNow; // @[storeDataIssue.scala 172:29]
  assign sdiFifo_modifyVal = map_sdiFifo_modifyVal_MPORT_data; // @[storeDataIssue.scala 169:21]
  assign sdiFifo_modify = fromBranch_valid & ~fromBranch_passOrFail; // @[storeDataIssue.scala 170:41]
  always @(posedge clock) begin
    if (map_MPORT_en & map_MPORT_mask) begin
      map[map_MPORT_addr] <= map_MPORT_data; // @[storeDataIssue.scala 152:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    map[initvar] = _RAND_0[3:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module rob_Anon(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [101:0] io_enq_bits,
  input          io_deq_ready,
  output         io_deq_valid,
  output [101:0] io_deq_bits,
  input          modify,
  input  [3:0]   modifyVal
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [101:0] memReg [0:15]; // @[Fifo.scala 86:19]
  wire  memReg_io_deq_bits_MPORT_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_io_deq_bits_MPORT_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_io_deq_bits_MPORT_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_2_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_2_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_2_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_3_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_3_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_3_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_4_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_4_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_4_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_5_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_5_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_5_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_6_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_6_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_6_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_7_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_7_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_7_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_8_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_8_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_8_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_9_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_9_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_9_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_10_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_10_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_10_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_11_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_11_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_11_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_12_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_12_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_12_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_13_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_13_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_13_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_14_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_14_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_14_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_15_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_15_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_15_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_16_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_16_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_16_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_17_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_17_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_17_data; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_data; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_addr; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_mask; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_en; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_1_data; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_1_addr; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_1_mask; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_1_en; // @[Fifo.scala 86:19]
  reg [3:0] readPtr; // @[Fifo.scala 75:25]
  wire [3:0] _nextRead_T_2 = readPtr + 4'h1; // @[Fifo.scala 76:61]
  wire [3:0] nextRead = readPtr == 4'hf ? 4'h0 : _nextRead_T_2; // @[Fifo.scala 76:21]
  wire  _T = io_deq_ready & io_deq_valid; // @[Fifo.scala 105:21]
  wire  _T_1 = io_deq_ready & io_deq_valid & io_enq_valid; // @[Fifo.scala 105:37]
  wire  _T_2 = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready; // @[Fifo.scala 105:53]
  wire  _T_3 = io_enq_valid & io_enq_ready; // @[Fifo.scala 109:27]
  wire  _GEN_14 = io_enq_valid & io_enq_ready ? 1'h0 : _T; // @[Fifo.scala 109:44]
  wire  incrRead = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready | _GEN_14; // @[Fifo.scala 105:70 108:14]
  reg [3:0] writePtr; // @[Fifo.scala 81:25]
  wire [3:0] _nextWrite_T_2 = writePtr + 4'h1; // @[Fifo.scala 82:65]
  wire [3:0] nextWrite = writePtr == 4'hf ? 4'h0 : _nextWrite_T_2; // @[Fifo.scala 82:22]
  reg  fullReg; // @[Fifo.scala 84:24]
  reg  emptyReg; // @[Fifo.scala 89:25]
  wire [3:0] _nextval_T_2 = modifyVal + 4'h1; // @[Fifo.scala 91:65]
  wire [3:0] nextval = modifyVal == 4'hf ? 4'h0 : _nextval_T_2; // @[Fifo.scala 91:20]
  wire  incrWrite = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready | _T_3; // @[Fifo.scala 105:70 107:15]
  wire  _GEN_3 = modify ? nextval == readPtr : fullReg; // @[Fifo.scala 93:16 96:13 84:24]
  wire  _GEN_5 = _T ? nextRead == writePtr : emptyReg; // @[Fifo.scala 114:44 116:14 89:25]
  wire  _GEN_12 = io_enq_valid & io_enq_ready ? 1'h0 : _GEN_5; // @[Fifo.scala 109:44 111:14]
  wire  _GEN_27 = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready ? emptyReg : _GEN_12; // @[Fifo.scala 105:70 89:25]
  wire  _io_enq_ready_T_3 = ~modify; // @[Fifo.scala 121:64]
  assign memReg_io_deq_bits_MPORT_en = 1'h1;
  assign memReg_io_deq_bits_MPORT_addr = readPtr;
  assign memReg_io_deq_bits_MPORT_data = memReg[memReg_io_deq_bits_MPORT_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_2_en = 1'h1;
  assign memReg_MPORT_2_addr = 4'h0;
  assign memReg_MPORT_2_data = memReg[memReg_MPORT_2_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_3_en = 1'h1;
  assign memReg_MPORT_3_addr = 4'h1;
  assign memReg_MPORT_3_data = memReg[memReg_MPORT_3_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_4_en = 1'h1;
  assign memReg_MPORT_4_addr = 4'h2;
  assign memReg_MPORT_4_data = memReg[memReg_MPORT_4_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_5_en = 1'h1;
  assign memReg_MPORT_5_addr = 4'h3;
  assign memReg_MPORT_5_data = memReg[memReg_MPORT_5_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_6_en = 1'h1;
  assign memReg_MPORT_6_addr = 4'h4;
  assign memReg_MPORT_6_data = memReg[memReg_MPORT_6_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_7_en = 1'h1;
  assign memReg_MPORT_7_addr = 4'h5;
  assign memReg_MPORT_7_data = memReg[memReg_MPORT_7_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_8_en = 1'h1;
  assign memReg_MPORT_8_addr = 4'h6;
  assign memReg_MPORT_8_data = memReg[memReg_MPORT_8_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_9_en = 1'h1;
  assign memReg_MPORT_9_addr = 4'h7;
  assign memReg_MPORT_9_data = memReg[memReg_MPORT_9_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_10_en = 1'h1;
  assign memReg_MPORT_10_addr = 4'h8;
  assign memReg_MPORT_10_data = memReg[memReg_MPORT_10_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_11_en = 1'h1;
  assign memReg_MPORT_11_addr = 4'h9;
  assign memReg_MPORT_11_data = memReg[memReg_MPORT_11_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_12_en = 1'h1;
  assign memReg_MPORT_12_addr = 4'ha;
  assign memReg_MPORT_12_data = memReg[memReg_MPORT_12_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_13_en = 1'h1;
  assign memReg_MPORT_13_addr = 4'hb;
  assign memReg_MPORT_13_data = memReg[memReg_MPORT_13_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_14_en = 1'h1;
  assign memReg_MPORT_14_addr = 4'hc;
  assign memReg_MPORT_14_data = memReg[memReg_MPORT_14_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_15_en = 1'h1;
  assign memReg_MPORT_15_addr = 4'hd;
  assign memReg_MPORT_15_data = memReg[memReg_MPORT_15_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_16_en = 1'h1;
  assign memReg_MPORT_16_addr = 4'he;
  assign memReg_MPORT_16_data = memReg[memReg_MPORT_16_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_17_en = 1'h1;
  assign memReg_MPORT_17_addr = 4'hf;
  assign memReg_MPORT_17_data = memReg[memReg_MPORT_17_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_data = io_enq_bits;
  assign memReg_MPORT_addr = writePtr;
  assign memReg_MPORT_mask = 1'h1;
  assign memReg_MPORT_en = _T_1 & io_enq_ready;
  assign memReg_MPORT_1_data = io_enq_bits;
  assign memReg_MPORT_1_addr = writePtr;
  assign memReg_MPORT_1_mask = 1'h1;
  assign memReg_MPORT_1_en = _T_2 ? 1'h0 : _T_3;
  assign io_enq_ready = (~fullReg | io_deq_valid & io_deq_ready) & ~modify; // @[Fifo.scala 121:62]
  assign io_deq_valid = ~emptyReg & _io_enq_ready_T_3; // @[Fifo.scala 122:29]
  assign io_deq_bits = memReg_io_deq_bits_MPORT_data; // @[Fifo.scala 120:15]
  always @(posedge clock) begin
    if (memReg_MPORT_en & memReg_MPORT_mask) begin
      memReg[memReg_MPORT_addr] <= memReg_MPORT_data; // @[Fifo.scala 86:19]
    end
    if (memReg_MPORT_1_en & memReg_MPORT_1_mask) begin
      memReg[memReg_MPORT_1_addr] <= memReg_MPORT_1_data; // @[Fifo.scala 86:19]
    end
    if (reset) begin // @[Fifo.scala 75:25]
      readPtr <= 4'h0; // @[Fifo.scala 75:25]
    end else if (incrRead) begin // @[Fifo.scala 77:19]
      if (readPtr == 4'hf) begin // @[Fifo.scala 76:21]
        readPtr <= 4'h0;
      end else begin
        readPtr <= _nextRead_T_2;
      end
    end
    if (reset) begin // @[Fifo.scala 81:25]
      writePtr <= 4'h0; // @[Fifo.scala 81:25]
    end else if (modify) begin // @[Fifo.scala 93:16]
      if (modifyVal == 4'hf) begin // @[Fifo.scala 91:20]
        writePtr <= 4'h0;
      end else begin
        writePtr <= _nextval_T_2;
      end
    end else if (incrWrite) begin // @[Fifo.scala 98:24]
      if (writePtr == 4'hf) begin // @[Fifo.scala 82:22]
        writePtr <= 4'h0;
      end else begin
        writePtr <= _nextWrite_T_2;
      end
    end
    if (reset) begin // @[Fifo.scala 84:24]
      fullReg <= 1'h0; // @[Fifo.scala 84:24]
    end else if (io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready) begin // @[Fifo.scala 105:70]
      fullReg <= _GEN_3;
    end else if (io_enq_valid & io_enq_ready) begin // @[Fifo.scala 109:44]
      fullReg <= nextWrite == readPtr; // @[Fifo.scala 112:13]
    end else if (_T) begin // @[Fifo.scala 114:44]
      fullReg <= 1'h0; // @[Fifo.scala 115:13]
    end else begin
      fullReg <= _GEN_3;
    end
    emptyReg <= reset | _GEN_27; // @[Fifo.scala 89:{25,25}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    memReg[initvar] = _RAND_0[101:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  readPtr = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  writePtr = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  fullReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  emptyReg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module rob_Anon_1(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [129:0] io_enq_bits,
  input          io_deq_ready,
  output         io_deq_valid,
  output [129:0] io_deq_bits,
  input          modify,
  input  [3:0]   modifyVal,
  input          writeports_0_valid,
  input  [129:0] writeports_0_data,
  input  [3:0]   writeports_0_addr,
  input          writeports_1_valid,
  input  [3:0]   writeports_1_addr,
  input          writeports_2_valid,
  input  [3:0]   writeports_2_addr,
  input          writeports_3_valid,
  input  [3:0]   writeports_3_addr,
  input          writeports_4_valid,
  input  [3:0]   writeports_4_addr,
  output [3:0]   allocatedAddr,
  output [3:0]   robAddrRelease
);
`ifdef RANDOMIZE_MEM_INIT
  reg [159:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [129:0] memReg [0:15]; // @[Fifo.scala 86:19]
  wire  memReg_io_deq_bits_MPORT_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_io_deq_bits_MPORT_addr; // @[Fifo.scala 86:19]
  wire [129:0] memReg_io_deq_bits_MPORT_data; // @[Fifo.scala 86:19]
  wire [129:0] memReg_MPORT_data; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_addr; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_mask; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_en; // @[Fifo.scala 86:19]
  wire [129:0] memReg_MPORT_1_data; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_1_addr; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_1_mask; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_1_en; // @[Fifo.scala 86:19]
  wire [129:0] memReg_MPORT_2_data; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_2_addr; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_2_mask; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_2_en; // @[Fifo.scala 86:19]
  wire [129:0] memReg_MPORT_3_data; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_3_addr; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_3_mask; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_3_en; // @[Fifo.scala 86:19]
  wire [129:0] memReg_MPORT_4_data; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_4_addr; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_4_mask; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_4_en; // @[Fifo.scala 86:19]
  wire [129:0] memReg_MPORT_5_data; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_5_addr; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_5_mask; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_5_en; // @[Fifo.scala 86:19]
  wire [129:0] memReg_MPORT_6_data; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_6_addr; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_6_mask; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_6_en; // @[Fifo.scala 86:19]
  reg [3:0] readPtr; // @[Fifo.scala 75:25]
  wire [3:0] _nextRead_T_2 = readPtr + 4'h1; // @[Fifo.scala 76:61]
  wire [3:0] nextRead = readPtr == 4'hf ? 4'h0 : _nextRead_T_2; // @[Fifo.scala 76:21]
  wire  _T = io_deq_ready & io_deq_valid; // @[Fifo.scala 105:21]
  wire  _T_1 = io_deq_ready & io_deq_valid & io_enq_valid; // @[Fifo.scala 105:37]
  wire  _T_2 = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready; // @[Fifo.scala 105:53]
  wire  _T_3 = io_enq_valid & io_enq_ready; // @[Fifo.scala 109:27]
  wire  _GEN_14 = io_enq_valid & io_enq_ready ? 1'h0 : _T; // @[Fifo.scala 109:44]
  wire  incrRead = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready | _GEN_14; // @[Fifo.scala 105:70 108:14]
  reg [3:0] writePtr; // @[Fifo.scala 81:25]
  wire [3:0] _nextWrite_T_2 = writePtr + 4'h1; // @[Fifo.scala 82:65]
  wire [3:0] nextWrite = writePtr == 4'hf ? 4'h0 : _nextWrite_T_2; // @[Fifo.scala 82:22]
  reg  fullReg; // @[Fifo.scala 84:24]
  reg  emptyReg; // @[Fifo.scala 89:25]
  wire [3:0] _nextval_T_2 = modifyVal + 4'h1; // @[Fifo.scala 91:65]
  wire [3:0] nextval = modifyVal == 4'hf ? 4'h0 : _nextval_T_2; // @[Fifo.scala 91:20]
  wire  incrWrite = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready | _T_3; // @[Fifo.scala 105:70 107:15]
  wire  _GEN_3 = modify ? nextval == readPtr : fullReg; // @[Fifo.scala 93:16 96:13 84:24]
  wire  _GEN_5 = _T ? nextRead == writePtr : emptyReg; // @[Fifo.scala 114:44 116:14 89:25]
  wire  _GEN_12 = io_enq_valid & io_enq_ready ? 1'h0 : _GEN_5; // @[Fifo.scala 109:44 111:14]
  wire  _GEN_27 = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready ? emptyReg : _GEN_12; // @[Fifo.scala 105:70 89:25]
  wire  _io_enq_ready_T_3 = ~modify; // @[Fifo.scala 121:64]
  assign memReg_io_deq_bits_MPORT_en = 1'h1;
  assign memReg_io_deq_bits_MPORT_addr = readPtr;
  assign memReg_io_deq_bits_MPORT_data = memReg[memReg_io_deq_bits_MPORT_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_data = io_enq_bits;
  assign memReg_MPORT_addr = writePtr;
  assign memReg_MPORT_mask = 1'h1;
  assign memReg_MPORT_en = _T_1 & io_enq_ready;
  assign memReg_MPORT_1_data = io_enq_bits;
  assign memReg_MPORT_1_addr = writePtr;
  assign memReg_MPORT_1_mask = 1'h1;
  assign memReg_MPORT_1_en = _T_2 ? 1'h0 : _T_3;
  assign memReg_MPORT_2_data = writeports_0_data;
  assign memReg_MPORT_2_addr = writeports_0_addr;
  assign memReg_MPORT_2_mask = 1'h1;
  assign memReg_MPORT_2_en = writeports_0_valid;
  assign memReg_MPORT_3_data = 130'h1;
  assign memReg_MPORT_3_addr = writeports_1_addr;
  assign memReg_MPORT_3_mask = 1'h1;
  assign memReg_MPORT_3_en = writeports_1_valid;
  assign memReg_MPORT_4_data = 130'h1;
  assign memReg_MPORT_4_addr = writeports_2_addr;
  assign memReg_MPORT_4_mask = 1'h1;
  assign memReg_MPORT_4_en = writeports_2_valid;
  assign memReg_MPORT_5_data = 130'h1;
  assign memReg_MPORT_5_addr = writeports_3_addr;
  assign memReg_MPORT_5_mask = 1'h1;
  assign memReg_MPORT_5_en = writeports_3_valid;
  assign memReg_MPORT_6_data = 130'h1;
  assign memReg_MPORT_6_addr = writeports_4_addr;
  assign memReg_MPORT_6_mask = 1'h1;
  assign memReg_MPORT_6_en = writeports_4_valid;
  assign io_enq_ready = (~fullReg | io_deq_valid & io_deq_ready) & ~modify; // @[Fifo.scala 121:62]
  assign io_deq_valid = ~emptyReg & _io_enq_ready_T_3; // @[Fifo.scala 122:29]
  assign io_deq_bits = memReg_io_deq_bits_MPORT_data; // @[Fifo.scala 120:15]
  assign allocatedAddr = writePtr; // @[Fifo.scala 145:17]
  assign robAddrRelease = readPtr; // @[rob.scala 63:20]
  always @(posedge clock) begin
    if (memReg_MPORT_en & memReg_MPORT_mask) begin
      memReg[memReg_MPORT_addr] <= memReg_MPORT_data; // @[Fifo.scala 86:19]
    end
    if (memReg_MPORT_1_en & memReg_MPORT_1_mask) begin
      memReg[memReg_MPORT_1_addr] <= memReg_MPORT_1_data; // @[Fifo.scala 86:19]
    end
    if (memReg_MPORT_2_en & memReg_MPORT_2_mask) begin
      memReg[memReg_MPORT_2_addr] <= memReg_MPORT_2_data; // @[Fifo.scala 86:19]
    end
    if (memReg_MPORT_3_en & memReg_MPORT_3_mask) begin
      memReg[memReg_MPORT_3_addr] <= memReg_MPORT_3_data; // @[Fifo.scala 86:19]
    end
    if (memReg_MPORT_4_en & memReg_MPORT_4_mask) begin
      memReg[memReg_MPORT_4_addr] <= memReg_MPORT_4_data; // @[Fifo.scala 86:19]
    end
    if (memReg_MPORT_5_en & memReg_MPORT_5_mask) begin
      memReg[memReg_MPORT_5_addr] <= memReg_MPORT_5_data; // @[Fifo.scala 86:19]
    end
    if (memReg_MPORT_6_en & memReg_MPORT_6_mask) begin
      memReg[memReg_MPORT_6_addr] <= memReg_MPORT_6_data; // @[Fifo.scala 86:19]
    end
    if (reset) begin // @[Fifo.scala 75:25]
      readPtr <= 4'h0; // @[Fifo.scala 75:25]
    end else if (incrRead) begin // @[Fifo.scala 77:19]
      if (readPtr == 4'hf) begin // @[Fifo.scala 76:21]
        readPtr <= 4'h0;
      end else begin
        readPtr <= _nextRead_T_2;
      end
    end
    if (reset) begin // @[Fifo.scala 81:25]
      writePtr <= 4'h0; // @[Fifo.scala 81:25]
    end else if (modify) begin // @[Fifo.scala 93:16]
      if (modifyVal == 4'hf) begin // @[Fifo.scala 91:20]
        writePtr <= 4'h0;
      end else begin
        writePtr <= _nextval_T_2;
      end
    end else if (incrWrite) begin // @[Fifo.scala 98:24]
      if (writePtr == 4'hf) begin // @[Fifo.scala 82:22]
        writePtr <= 4'h0;
      end else begin
        writePtr <= _nextWrite_T_2;
      end
    end
    if (reset) begin // @[Fifo.scala 84:24]
      fullReg <= 1'h0; // @[Fifo.scala 84:24]
    end else if (io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready) begin // @[Fifo.scala 105:70]
      fullReg <= _GEN_3;
    end else if (io_enq_valid & io_enq_ready) begin // @[Fifo.scala 109:44]
      fullReg <= nextWrite == readPtr; // @[Fifo.scala 112:13]
    end else if (_T) begin // @[Fifo.scala 114:44]
      fullReg <= 1'h0; // @[Fifo.scala 115:13]
    end else begin
      fullReg <= _GEN_3;
    end
    emptyReg <= reset | _GEN_27; // @[Fifo.scala 89:{25,25}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {5{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    memReg[initvar] = _RAND_0[129:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  readPtr = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  writePtr = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  fullReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  emptyReg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module rob(
  input         clock,
  input         reset,
  output        allocate_ready,
  input         allocate_fired,
  input  [63:0] allocate_pc,
  input  [31:0] allocate_instruction,
  input  [5:0]  allocate_prfDest,
  output [3:0]  allocate_robAddr,
  input         allocate_isReady,
  output        commit_ready,
  input         commit_fired,
  output [5:0]  commit_prfDest,
  output [63:0] commit_pc,
  output [31:0] commit_instruction,
  output        commit_exceptionOccurred,
  output [63:0] commit_mtval,
  output        commit_isStore,
  output        commit_is_fence,
  output [3:0]  commit_robAddr,
  input         branch_valid,
  input         branch_pass,
  input  [3:0]  branch_robAddr,
  input  [3:0]  execPorts_0_robAddr,
  input  [63:0] execPorts_0_mtval,
  input         execPorts_0_valid,
  input  [3:0]  execPorts_1_robAddr,
  input         execPorts_1_valid,
  input  [3:0]  execPorts_2_robAddr,
  input         execPorts_2_valid,
  input  [3:0]  execPorts_3_robAddr,
  input         execPorts_3_valid
);
  wire  fifo_clock; // @[rob.scala 24:20]
  wire  fifo_reset; // @[rob.scala 24:20]
  wire  fifo_io_enq_ready; // @[rob.scala 24:20]
  wire  fifo_io_enq_valid; // @[rob.scala 24:20]
  wire [101:0] fifo_io_enq_bits; // @[rob.scala 24:20]
  wire  fifo_io_deq_ready; // @[rob.scala 24:20]
  wire  fifo_io_deq_valid; // @[rob.scala 24:20]
  wire [101:0] fifo_io_deq_bits; // @[rob.scala 24:20]
  wire  fifo_modify; // @[rob.scala 24:20]
  wire [3:0] fifo_modifyVal; // @[rob.scala 24:20]
  wire  results_clock; // @[rob.scala 61:23]
  wire  results_reset; // @[rob.scala 61:23]
  wire  results_io_enq_ready; // @[rob.scala 61:23]
  wire  results_io_enq_valid; // @[rob.scala 61:23]
  wire [129:0] results_io_enq_bits; // @[rob.scala 61:23]
  wire  results_io_deq_ready; // @[rob.scala 61:23]
  wire  results_io_deq_valid; // @[rob.scala 61:23]
  wire [129:0] results_io_deq_bits; // @[rob.scala 61:23]
  wire  results_modify; // @[rob.scala 61:23]
  wire [3:0] results_modifyVal; // @[rob.scala 61:23]
  wire  results_writeports_0_valid; // @[rob.scala 61:23]
  wire [129:0] results_writeports_0_data; // @[rob.scala 61:23]
  wire [3:0] results_writeports_0_addr; // @[rob.scala 61:23]
  wire  results_writeports_1_valid; // @[rob.scala 61:23]
  wire [3:0] results_writeports_1_addr; // @[rob.scala 61:23]
  wire  results_writeports_2_valid; // @[rob.scala 61:23]
  wire [3:0] results_writeports_2_addr; // @[rob.scala 61:23]
  wire  results_writeports_3_valid; // @[rob.scala 61:23]
  wire [3:0] results_writeports_3_addr; // @[rob.scala 61:23]
  wire  results_writeports_4_valid; // @[rob.scala 61:23]
  wire [3:0] results_writeports_4_addr; // @[rob.scala 61:23]
  wire [3:0] results_allocatedAddr; // @[rob.scala 61:23]
  wire [3:0] results_robAddrRelease; // @[rob.scala 61:23]
  wire [37:0] _fifo_data_T = {allocate_instruction,allocate_prfDest}; // @[Cat.scala 33:92]
  wire  is_fence = commit_instruction[6:0] == 7'hf; // @[rob.scala 81:42]
  wire  _fifo_modify_T = ~branch_pass; // @[rob.scala 105:33]
  wire [128:0] _writeval_T_1 = {execPorts_0_mtval,65'h1}; // @[Cat.scala 33:92]
  rob_Anon fifo ( // @[rob.scala 24:20]
    .clock(fifo_clock),
    .reset(fifo_reset),
    .io_enq_ready(fifo_io_enq_ready),
    .io_enq_valid(fifo_io_enq_valid),
    .io_enq_bits(fifo_io_enq_bits),
    .io_deq_ready(fifo_io_deq_ready),
    .io_deq_valid(fifo_io_deq_valid),
    .io_deq_bits(fifo_io_deq_bits),
    .modify(fifo_modify),
    .modifyVal(fifo_modifyVal)
  );
  rob_Anon_1 results ( // @[rob.scala 61:23]
    .clock(results_clock),
    .reset(results_reset),
    .io_enq_ready(results_io_enq_ready),
    .io_enq_valid(results_io_enq_valid),
    .io_enq_bits(results_io_enq_bits),
    .io_deq_ready(results_io_deq_ready),
    .io_deq_valid(results_io_deq_valid),
    .io_deq_bits(results_io_deq_bits),
    .modify(results_modify),
    .modifyVal(results_modifyVal),
    .writeports_0_valid(results_writeports_0_valid),
    .writeports_0_data(results_writeports_0_data),
    .writeports_0_addr(results_writeports_0_addr),
    .writeports_1_valid(results_writeports_1_valid),
    .writeports_1_addr(results_writeports_1_addr),
    .writeports_2_valid(results_writeports_2_valid),
    .writeports_2_addr(results_writeports_2_addr),
    .writeports_3_valid(results_writeports_3_valid),
    .writeports_3_addr(results_writeports_3_addr),
    .writeports_4_valid(results_writeports_4_valid),
    .writeports_4_addr(results_writeports_4_addr),
    .allocatedAddr(results_allocatedAddr),
    .robAddrRelease(results_robAddrRelease)
  );
  assign allocate_ready = commit_ready & ~commit_fired ? 1'h0 : fifo_io_enq_ready & results_io_enq_ready; // @[rob.scala 142:{39,56} 67:18]
  assign allocate_robAddr = results_allocatedAddr; // @[rob.scala 72:20]
  assign commit_ready = (results_io_deq_bits[0] | is_fence | commit_isStore) & fifo_io_deq_valid & results_io_deq_valid; // @[rob.scala 84:92]
  assign commit_prfDest = fifo_io_deq_bits[5:0]; // @[rob.scala 88:37]
  assign commit_pc = fifo_io_deq_bits[101:38]; // @[rob.scala 90:32]
  assign commit_instruction = fifo_io_deq_bits[37:6]; // @[rob.scala 89:41]
  assign commit_exceptionOccurred = results_io_deq_bits[129]; // @[rob.scala 87:50]
  assign commit_mtval = results_io_deq_bits[128:65]; // @[rob.scala 86:38]
  assign commit_isStore = fifo_io_deq_bits[12:6] == 7'h23; // @[rob.scala 102:44]
  assign commit_is_fence = commit_instruction[6:0] == 7'hf; // @[rob.scala 81:42]
  assign commit_robAddr = results_robAddrRelease; // @[rob.scala 92:18]
  assign fifo_clock = clock;
  assign fifo_reset = commit_exceptionOccurred & commit_fired | reset; // @[rob.scala 123:49 124:19]
  assign fifo_io_enq_valid = allocate_fired; // @[rob.scala 73:23 74:23 77:23]
  assign fifo_io_enq_bits = {allocate_pc,_fifo_data_T}; // @[Cat.scala 33:92]
  assign fifo_io_deq_ready = commit_fired; // @[rob.scala 94:22 95:23 98:23]
  assign fifo_modify = branch_valid & ~branch_pass; // @[rob.scala 105:31]
  assign fifo_modifyVal = branch_robAddr; // @[rob.scala 106:18]
  assign results_clock = clock;
  assign results_reset = commit_exceptionOccurred & commit_fired | reset; // @[rob.scala 123:49 124:19]
  assign results_io_enq_valid = allocate_fired; // @[rob.scala 73:23 74:23 77:23]
  assign results_io_enq_bits = {129'h0,allocate_isReady}; // @[Cat.scala 33:92]
  assign results_io_deq_ready = commit_fired; // @[rob.scala 94:22 95:23 98:23]
  assign results_modify = branch_valid & _fifo_modify_T; // @[rob.scala 107:34]
  assign results_modifyVal = branch_robAddr; // @[rob.scala 108:21]
  assign results_writeports_0_valid = execPorts_0_valid; // @[rob.scala 117:33]
  assign results_writeports_0_data = {1'h0,_writeval_T_1}; // @[Cat.scala 33:92]
  assign results_writeports_0_addr = execPorts_0_robAddr; // @[rob.scala 119:32]
  assign results_writeports_1_valid = execPorts_1_valid; // @[rob.scala 117:33]
  assign results_writeports_1_addr = execPorts_1_robAddr; // @[rob.scala 119:32]
  assign results_writeports_2_valid = execPorts_2_valid; // @[rob.scala 117:33]
  assign results_writeports_2_addr = execPorts_2_robAddr; // @[rob.scala 119:32]
  assign results_writeports_3_valid = execPorts_3_valid; // @[rob.scala 117:33]
  assign results_writeports_3_addr = execPorts_3_robAddr; // @[rob.scala 119:32]
  assign results_writeports_4_valid = branch_valid; // @[rob.scala 109:43]
  assign results_writeports_4_addr = branch_robAddr; // @[rob.scala 110:42]
endmodule
module scheduler(
  input         clock,
  input         reset,
  output        allocate_ready,
  input         allocate_fired,
  input  [31:0] allocate_instruction,
  input  [4:0]  allocate_branchMask,
  input         allocate_rs1_ready,
  input  [5:0]  allocate_rs1_prfAddr,
  input         allocate_rs2_ready,
  input  [5:0]  allocate_rs2_prfAddr,
  input  [5:0]  allocate_prfDest,
  input  [3:0]  allocate_robAddr,
  output        release_ready,
  input         release_fired,
  output [31:0] release_instruction,
  output [4:0]  release_branchMask,
  output [5:0]  release_rs1prfAddr,
  output [5:0]  release_rs2prfAddr,
  output [5:0]  release_prfDest,
  output [3:0]  release_robAddr,
  input         wakeUpExt_0_valid,
  input  [5:0]  wakeUpExt_0_prfAddr,
  input         wakeUpExt_1_valid,
  input  [5:0]  wakeUpExt_1_prfAddr,
  input         branchOps_valid,
  input  [4:0]  branchOps_branchMask,
  input         branchOps_passed,
  input         memoryReady,
  input         multuplyAndDivideReady,
  output        instrRetired_valid,
  output [5:0]  instrRetired_prfAddr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
`endif // RANDOMIZE_REG_INIT
  reg  queue_0_opcodeMeta_isBranch; // @[scheduler.scala 26:22]
  reg  queue_0_opcodeMeta_isMemAccess; // @[scheduler.scala 26:22]
  reg  queue_0_opcodeMeta_isM; // @[scheduler.scala 26:22]
  reg  queue_0_valid; // @[scheduler.scala 26:22]
  reg [31:0] queue_0_instruction; // @[scheduler.scala 26:22]
  reg [4:0] queue_0_branchMask; // @[scheduler.scala 26:22]
  reg  queue_0_rs1_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_0_rs1_prfAddr; // @[scheduler.scala 26:22]
  reg  queue_0_rs2_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_0_rs2_prfAddr; // @[scheduler.scala 26:22]
  reg [5:0] queue_0_prfDest; // @[scheduler.scala 26:22]
  reg [3:0] queue_0_robAddr; // @[scheduler.scala 26:22]
  reg  queue_1_opcodeMeta_isBranch; // @[scheduler.scala 26:22]
  reg  queue_1_opcodeMeta_isMemAccess; // @[scheduler.scala 26:22]
  reg  queue_1_opcodeMeta_isM; // @[scheduler.scala 26:22]
  reg  queue_1_valid; // @[scheduler.scala 26:22]
  reg [31:0] queue_1_instruction; // @[scheduler.scala 26:22]
  reg [4:0] queue_1_branchMask; // @[scheduler.scala 26:22]
  reg  queue_1_rs1_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_1_rs1_prfAddr; // @[scheduler.scala 26:22]
  reg  queue_1_rs2_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_1_rs2_prfAddr; // @[scheduler.scala 26:22]
  reg [5:0] queue_1_prfDest; // @[scheduler.scala 26:22]
  reg [3:0] queue_1_robAddr; // @[scheduler.scala 26:22]
  reg  queue_2_opcodeMeta_isBranch; // @[scheduler.scala 26:22]
  reg  queue_2_opcodeMeta_isMemAccess; // @[scheduler.scala 26:22]
  reg  queue_2_opcodeMeta_isM; // @[scheduler.scala 26:22]
  reg  queue_2_valid; // @[scheduler.scala 26:22]
  reg [31:0] queue_2_instruction; // @[scheduler.scala 26:22]
  reg [4:0] queue_2_branchMask; // @[scheduler.scala 26:22]
  reg  queue_2_rs1_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_2_rs1_prfAddr; // @[scheduler.scala 26:22]
  reg  queue_2_rs2_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_2_rs2_prfAddr; // @[scheduler.scala 26:22]
  reg [5:0] queue_2_prfDest; // @[scheduler.scala 26:22]
  reg [3:0] queue_2_robAddr; // @[scheduler.scala 26:22]
  reg  queue_3_opcodeMeta_isBranch; // @[scheduler.scala 26:22]
  reg  queue_3_opcodeMeta_isMemAccess; // @[scheduler.scala 26:22]
  reg  queue_3_opcodeMeta_isM; // @[scheduler.scala 26:22]
  reg  queue_3_valid; // @[scheduler.scala 26:22]
  reg [31:0] queue_3_instruction; // @[scheduler.scala 26:22]
  reg [4:0] queue_3_branchMask; // @[scheduler.scala 26:22]
  reg  queue_3_rs1_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_3_rs1_prfAddr; // @[scheduler.scala 26:22]
  reg  queue_3_rs2_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_3_rs2_prfAddr; // @[scheduler.scala 26:22]
  reg [5:0] queue_3_prfDest; // @[scheduler.scala 26:22]
  reg [3:0] queue_3_robAddr; // @[scheduler.scala 26:22]
  reg  queue_4_opcodeMeta_isBranch; // @[scheduler.scala 26:22]
  reg  queue_4_opcodeMeta_isMemAccess; // @[scheduler.scala 26:22]
  reg  queue_4_opcodeMeta_isM; // @[scheduler.scala 26:22]
  reg  queue_4_valid; // @[scheduler.scala 26:22]
  reg [31:0] queue_4_instruction; // @[scheduler.scala 26:22]
  reg [4:0] queue_4_branchMask; // @[scheduler.scala 26:22]
  reg  queue_4_rs1_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_4_rs1_prfAddr; // @[scheduler.scala 26:22]
  reg  queue_4_rs2_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_4_rs2_prfAddr; // @[scheduler.scala 26:22]
  reg [5:0] queue_4_prfDest; // @[scheduler.scala 26:22]
  reg [3:0] queue_4_robAddr; // @[scheduler.scala 26:22]
  reg  queue_5_opcodeMeta_isBranch; // @[scheduler.scala 26:22]
  reg  queue_5_opcodeMeta_isMemAccess; // @[scheduler.scala 26:22]
  reg  queue_5_opcodeMeta_isM; // @[scheduler.scala 26:22]
  reg  queue_5_valid; // @[scheduler.scala 26:22]
  reg [31:0] queue_5_instruction; // @[scheduler.scala 26:22]
  reg [4:0] queue_5_branchMask; // @[scheduler.scala 26:22]
  reg  queue_5_rs1_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_5_rs1_prfAddr; // @[scheduler.scala 26:22]
  reg  queue_5_rs2_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_5_rs2_prfAddr; // @[scheduler.scala 26:22]
  reg [5:0] queue_5_prfDest; // @[scheduler.scala 26:22]
  reg [3:0] queue_5_robAddr; // @[scheduler.scala 26:22]
  reg  queue_6_opcodeMeta_isBranch; // @[scheduler.scala 26:22]
  reg  queue_6_opcodeMeta_isMemAccess; // @[scheduler.scala 26:22]
  reg  queue_6_opcodeMeta_isM; // @[scheduler.scala 26:22]
  reg  queue_6_valid; // @[scheduler.scala 26:22]
  reg [31:0] queue_6_instruction; // @[scheduler.scala 26:22]
  reg [4:0] queue_6_branchMask; // @[scheduler.scala 26:22]
  reg  queue_6_rs1_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_6_rs1_prfAddr; // @[scheduler.scala 26:22]
  reg  queue_6_rs2_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_6_rs2_prfAddr; // @[scheduler.scala 26:22]
  reg [5:0] queue_6_prfDest; // @[scheduler.scala 26:22]
  reg [3:0] queue_6_robAddr; // @[scheduler.scala 26:22]
  reg  queue_7_opcodeMeta_isBranch; // @[scheduler.scala 26:22]
  reg  queue_7_opcodeMeta_isMemAccess; // @[scheduler.scala 26:22]
  reg  queue_7_opcodeMeta_isM; // @[scheduler.scala 26:22]
  reg  queue_7_valid; // @[scheduler.scala 26:22]
  reg [31:0] queue_7_instruction; // @[scheduler.scala 26:22]
  reg [4:0] queue_7_branchMask; // @[scheduler.scala 26:22]
  reg  queue_7_rs1_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_7_rs1_prfAddr; // @[scheduler.scala 26:22]
  reg  queue_7_rs2_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_7_rs2_prfAddr; // @[scheduler.scala 26:22]
  reg [5:0] queue_7_prfDest; // @[scheduler.scala 26:22]
  reg [3:0] queue_7_robAddr; // @[scheduler.scala 26:22]
  wire  _readyVector_T_1 = queue_0_valid & queue_0_rs1_ready & queue_0_rs2_ready; // @[scheduler.scala 51:42]
  wire  _readyVector_T_7 = ~queue_0_opcodeMeta_isMemAccess | memoryReady; // @[scheduler.scala 53:39]
  wire  _readyVector_T_8 = _readyVector_T_1 & _readyVector_T_7; // @[scheduler.scala 52:151]
  wire  _readyVector_T_10 = ~queue_0_opcodeMeta_isM | multuplyAndDivideReady; // @[scheduler.scala 54:31]
  wire  _readyVector_T_11 = _readyVector_T_8 & _readyVector_T_10; // @[scheduler.scala 53:174]
  wire  _readyVector_T_17 = ~queue_1_opcodeMeta_isBranch | ~(queue_0_valid & queue_0_opcodeMeta_isBranch); // @[scheduler.scala 52:36]
  wire  _readyVector_T_18 = queue_1_valid & queue_1_rs1_ready & queue_1_rs2_ready & _readyVector_T_17; // @[scheduler.scala 51:64]
  wire  _readyVector_T_23 = ~queue_1_opcodeMeta_isMemAccess | ~(queue_0_valid & queue_0_opcodeMeta_isMemAccess) &
    memoryReady; // @[scheduler.scala 53:39]
  wire  _readyVector_T_24 = _readyVector_T_18 & _readyVector_T_23; // @[scheduler.scala 52:151]
  wire  _readyVector_T_26 = ~queue_1_opcodeMeta_isM | multuplyAndDivideReady; // @[scheduler.scala 54:31]
  wire  _readyVector_T_27 = _readyVector_T_24 & _readyVector_T_26; // @[scheduler.scala 53:174]
  wire  _readyVector_T_35 = ~queue_2_opcodeMeta_isBranch | ~(queue_0_valid & queue_0_opcodeMeta_isBranch | queue_1_valid
     & queue_1_opcodeMeta_isBranch); // @[scheduler.scala 52:36]
  wire  _readyVector_T_36 = queue_2_valid & queue_2_rs1_ready & queue_2_rs2_ready & _readyVector_T_35; // @[scheduler.scala 51:64]
  wire  _readyVector_T_43 = ~queue_2_opcodeMeta_isMemAccess | ~(queue_0_valid & queue_0_opcodeMeta_isMemAccess |
    queue_1_valid & queue_1_opcodeMeta_isMemAccess) & memoryReady; // @[scheduler.scala 53:39]
  wire  _readyVector_T_44 = _readyVector_T_36 & _readyVector_T_43; // @[scheduler.scala 52:151]
  wire  _readyVector_T_46 = ~queue_2_opcodeMeta_isM | multuplyAndDivideReady; // @[scheduler.scala 54:31]
  wire  _readyVector_T_47 = _readyVector_T_44 & _readyVector_T_46; // @[scheduler.scala 53:174]
  wire  _readyVector_T_57 = ~queue_3_opcodeMeta_isBranch | ~(queue_0_valid & queue_0_opcodeMeta_isBranch | queue_1_valid
     & queue_1_opcodeMeta_isBranch | queue_2_valid & queue_2_opcodeMeta_isBranch); // @[scheduler.scala 52:36]
  wire  _readyVector_T_58 = queue_3_valid & queue_3_rs1_ready & queue_3_rs2_ready & _readyVector_T_57; // @[scheduler.scala 51:64]
  wire  _readyVector_T_67 = ~queue_3_opcodeMeta_isMemAccess | ~(queue_0_valid & queue_0_opcodeMeta_isMemAccess |
    queue_1_valid & queue_1_opcodeMeta_isMemAccess | queue_2_valid & queue_2_opcodeMeta_isMemAccess) & memoryReady; // @[scheduler.scala 53:39]
  wire  _readyVector_T_68 = _readyVector_T_58 & _readyVector_T_67; // @[scheduler.scala 52:151]
  wire  _readyVector_T_70 = ~queue_3_opcodeMeta_isM | multuplyAndDivideReady; // @[scheduler.scala 54:31]
  wire  _readyVector_T_71 = _readyVector_T_68 & _readyVector_T_70; // @[scheduler.scala 53:174]
  wire  _readyVector_T_83 = ~queue_4_opcodeMeta_isBranch | ~(queue_0_valid & queue_0_opcodeMeta_isBranch | queue_1_valid
     & queue_1_opcodeMeta_isBranch | queue_2_valid & queue_2_opcodeMeta_isBranch | queue_3_valid &
    queue_3_opcodeMeta_isBranch); // @[scheduler.scala 52:36]
  wire  _readyVector_T_84 = queue_4_valid & queue_4_rs1_ready & queue_4_rs2_ready & _readyVector_T_83; // @[scheduler.scala 51:64]
  wire  _readyVector_T_95 = ~queue_4_opcodeMeta_isMemAccess | ~(queue_0_valid & queue_0_opcodeMeta_isMemAccess |
    queue_1_valid & queue_1_opcodeMeta_isMemAccess | queue_2_valid & queue_2_opcodeMeta_isMemAccess | queue_3_valid &
    queue_3_opcodeMeta_isMemAccess) & memoryReady; // @[scheduler.scala 53:39]
  wire  _readyVector_T_96 = _readyVector_T_84 & _readyVector_T_95; // @[scheduler.scala 52:151]
  wire  _readyVector_T_98 = ~queue_4_opcodeMeta_isM | multuplyAndDivideReady; // @[scheduler.scala 54:31]
  wire  _readyVector_T_99 = _readyVector_T_96 & _readyVector_T_98; // @[scheduler.scala 53:174]
  wire  _readyVector_T_113 = ~queue_5_opcodeMeta_isBranch | ~(queue_0_valid & queue_0_opcodeMeta_isBranch |
    queue_1_valid & queue_1_opcodeMeta_isBranch | queue_2_valid & queue_2_opcodeMeta_isBranch | queue_3_valid &
    queue_3_opcodeMeta_isBranch | queue_4_valid & queue_4_opcodeMeta_isBranch); // @[scheduler.scala 52:36]
  wire  _readyVector_T_114 = queue_5_valid & queue_5_rs1_ready & queue_5_rs2_ready & _readyVector_T_113; // @[scheduler.scala 51:64]
  wire  _readyVector_T_127 = ~queue_5_opcodeMeta_isMemAccess | ~(queue_0_valid & queue_0_opcodeMeta_isMemAccess |
    queue_1_valid & queue_1_opcodeMeta_isMemAccess | queue_2_valid & queue_2_opcodeMeta_isMemAccess | queue_3_valid &
    queue_3_opcodeMeta_isMemAccess | queue_4_valid & queue_4_opcodeMeta_isMemAccess) & memoryReady; // @[scheduler.scala 53:39]
  wire  _readyVector_T_128 = _readyVector_T_114 & _readyVector_T_127; // @[scheduler.scala 52:151]
  wire  _readyVector_T_130 = ~queue_5_opcodeMeta_isM | multuplyAndDivideReady; // @[scheduler.scala 54:31]
  wire  _readyVector_T_131 = _readyVector_T_128 & _readyVector_T_130; // @[scheduler.scala 53:174]
  wire  _readyVector_T_147 = ~queue_6_opcodeMeta_isBranch | ~(queue_0_valid & queue_0_opcodeMeta_isBranch |
    queue_1_valid & queue_1_opcodeMeta_isBranch | queue_2_valid & queue_2_opcodeMeta_isBranch | queue_3_valid &
    queue_3_opcodeMeta_isBranch | queue_4_valid & queue_4_opcodeMeta_isBranch | queue_5_valid &
    queue_5_opcodeMeta_isBranch); // @[scheduler.scala 52:36]
  wire  _readyVector_T_148 = queue_6_valid & queue_6_rs1_ready & queue_6_rs2_ready & _readyVector_T_147; // @[scheduler.scala 51:64]
  wire  _readyVector_T_163 = ~queue_6_opcodeMeta_isMemAccess | ~(queue_0_valid & queue_0_opcodeMeta_isMemAccess |
    queue_1_valid & queue_1_opcodeMeta_isMemAccess | queue_2_valid & queue_2_opcodeMeta_isMemAccess | queue_3_valid &
    queue_3_opcodeMeta_isMemAccess | queue_4_valid & queue_4_opcodeMeta_isMemAccess | queue_5_valid &
    queue_5_opcodeMeta_isMemAccess) & memoryReady; // @[scheduler.scala 53:39]
  wire  _readyVector_T_164 = _readyVector_T_148 & _readyVector_T_163; // @[scheduler.scala 52:151]
  wire  _readyVector_T_166 = ~queue_6_opcodeMeta_isM | multuplyAndDivideReady; // @[scheduler.scala 54:31]
  wire  _readyVector_T_167 = _readyVector_T_164 & _readyVector_T_166; // @[scheduler.scala 53:174]
  wire  _readyVector_T_185 = ~queue_7_opcodeMeta_isBranch | ~(queue_0_valid & queue_0_opcodeMeta_isBranch |
    queue_1_valid & queue_1_opcodeMeta_isBranch | queue_2_valid & queue_2_opcodeMeta_isBranch | queue_3_valid &
    queue_3_opcodeMeta_isBranch | queue_4_valid & queue_4_opcodeMeta_isBranch | queue_5_valid &
    queue_5_opcodeMeta_isBranch | queue_6_valid & queue_6_opcodeMeta_isBranch); // @[scheduler.scala 52:36]
  wire  _readyVector_T_186 = queue_7_valid & queue_7_rs1_ready & queue_7_rs2_ready & _readyVector_T_185; // @[scheduler.scala 51:64]
  wire  _readyVector_T_203 = ~queue_7_opcodeMeta_isMemAccess | ~(queue_0_valid & queue_0_opcodeMeta_isMemAccess |
    queue_1_valid & queue_1_opcodeMeta_isMemAccess | queue_2_valid & queue_2_opcodeMeta_isMemAccess | queue_3_valid &
    queue_3_opcodeMeta_isMemAccess | queue_4_valid & queue_4_opcodeMeta_isMemAccess | queue_5_valid &
    queue_5_opcodeMeta_isMemAccess | queue_6_valid & queue_6_opcodeMeta_isMemAccess) & memoryReady; // @[scheduler.scala 53:39]
  wire  _readyVector_T_204 = _readyVector_T_186 & _readyVector_T_203; // @[scheduler.scala 52:151]
  wire  _readyVector_T_206 = ~queue_7_opcodeMeta_isM | multuplyAndDivideReady; // @[scheduler.scala 54:31]
  wire  _readyVector_T_207 = _readyVector_T_204 & _readyVector_T_206; // @[scheduler.scala 53:174]
  wire [7:0] readyVector = {_readyVector_T_207,_readyVector_T_167,_readyVector_T_131,_readyVector_T_99,_readyVector_T_71
    ,_readyVector_T_47,_readyVector_T_27,_readyVector_T_11}; // @[Cat.scala 33:92]
  wire [2:0] _dequeuedIndex_T_16 = readyVector[7] ? 3'h7 : 3'h0; // @[Mux.scala 101:16]
  wire [2:0] _dequeuedIndex_T_17 = readyVector[6] ? 3'h6 : _dequeuedIndex_T_16; // @[Mux.scala 101:16]
  wire [2:0] _dequeuedIndex_T_18 = readyVector[5] ? 3'h5 : _dequeuedIndex_T_17; // @[Mux.scala 101:16]
  wire [2:0] _dequeuedIndex_T_19 = readyVector[4] ? 3'h4 : _dequeuedIndex_T_18; // @[Mux.scala 101:16]
  wire [2:0] _dequeuedIndex_T_20 = readyVector[3] ? 3'h3 : _dequeuedIndex_T_19; // @[Mux.scala 101:16]
  wire [2:0] _dequeuedIndex_T_21 = readyVector[2] ? 3'h2 : _dequeuedIndex_T_20; // @[Mux.scala 101:16]
  wire [2:0] _dequeuedIndex_T_22 = readyVector[1] ? 3'h1 : _dequeuedIndex_T_21; // @[Mux.scala 101:16]
  wire [2:0] dequeuedIndex = readyVector[0] ? 3'h0 : _dequeuedIndex_T_22; // @[Mux.scala 101:16]
  wire  _dequeued_T_14_opcodeMeta_isM = readyVector[6] ? queue_6_opcodeMeta_isM : queue_7_opcodeMeta_isM; // @[Mux.scala 101:16]
  wire  _dequeued_T_14_valid = readyVector[6] ? queue_6_valid : queue_7_valid; // @[Mux.scala 101:16]
  wire [31:0] _dequeued_T_14_instruction = readyVector[6] ? queue_6_instruction : queue_7_instruction; // @[Mux.scala 101:16]
  wire [4:0] _dequeued_T_14_branchMask = readyVector[6] ? queue_6_branchMask : queue_7_branchMask; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_14_rs1_prfAddr = readyVector[6] ? queue_6_rs1_prfAddr : queue_7_rs1_prfAddr; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_14_rs2_prfAddr = readyVector[6] ? queue_6_rs2_prfAddr : queue_7_rs2_prfAddr; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_14_prfDest = readyVector[6] ? queue_6_prfDest : queue_7_prfDest; // @[Mux.scala 101:16]
  wire [3:0] _dequeued_T_14_robAddr = readyVector[6] ? queue_6_robAddr : queue_7_robAddr; // @[Mux.scala 101:16]
  wire  _dequeued_T_15_opcodeMeta_isM = readyVector[5] ? queue_5_opcodeMeta_isM : _dequeued_T_14_opcodeMeta_isM; // @[Mux.scala 101:16]
  wire  _dequeued_T_15_valid = readyVector[5] ? queue_5_valid : _dequeued_T_14_valid; // @[Mux.scala 101:16]
  wire [31:0] _dequeued_T_15_instruction = readyVector[5] ? queue_5_instruction : _dequeued_T_14_instruction; // @[Mux.scala 101:16]
  wire [4:0] _dequeued_T_15_branchMask = readyVector[5] ? queue_5_branchMask : _dequeued_T_14_branchMask; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_15_rs1_prfAddr = readyVector[5] ? queue_5_rs1_prfAddr : _dequeued_T_14_rs1_prfAddr; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_15_rs2_prfAddr = readyVector[5] ? queue_5_rs2_prfAddr : _dequeued_T_14_rs2_prfAddr; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_15_prfDest = readyVector[5] ? queue_5_prfDest : _dequeued_T_14_prfDest; // @[Mux.scala 101:16]
  wire [3:0] _dequeued_T_15_robAddr = readyVector[5] ? queue_5_robAddr : _dequeued_T_14_robAddr; // @[Mux.scala 101:16]
  wire  _dequeued_T_16_opcodeMeta_isM = readyVector[4] ? queue_4_opcodeMeta_isM : _dequeued_T_15_opcodeMeta_isM; // @[Mux.scala 101:16]
  wire  _dequeued_T_16_valid = readyVector[4] ? queue_4_valid : _dequeued_T_15_valid; // @[Mux.scala 101:16]
  wire [31:0] _dequeued_T_16_instruction = readyVector[4] ? queue_4_instruction : _dequeued_T_15_instruction; // @[Mux.scala 101:16]
  wire [4:0] _dequeued_T_16_branchMask = readyVector[4] ? queue_4_branchMask : _dequeued_T_15_branchMask; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_16_rs1_prfAddr = readyVector[4] ? queue_4_rs1_prfAddr : _dequeued_T_15_rs1_prfAddr; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_16_rs2_prfAddr = readyVector[4] ? queue_4_rs2_prfAddr : _dequeued_T_15_rs2_prfAddr; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_16_prfDest = readyVector[4] ? queue_4_prfDest : _dequeued_T_15_prfDest; // @[Mux.scala 101:16]
  wire [3:0] _dequeued_T_16_robAddr = readyVector[4] ? queue_4_robAddr : _dequeued_T_15_robAddr; // @[Mux.scala 101:16]
  wire  _dequeued_T_17_opcodeMeta_isM = readyVector[3] ? queue_3_opcodeMeta_isM : _dequeued_T_16_opcodeMeta_isM; // @[Mux.scala 101:16]
  wire  _dequeued_T_17_valid = readyVector[3] ? queue_3_valid : _dequeued_T_16_valid; // @[Mux.scala 101:16]
  wire [31:0] _dequeued_T_17_instruction = readyVector[3] ? queue_3_instruction : _dequeued_T_16_instruction; // @[Mux.scala 101:16]
  wire [4:0] _dequeued_T_17_branchMask = readyVector[3] ? queue_3_branchMask : _dequeued_T_16_branchMask; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_17_rs1_prfAddr = readyVector[3] ? queue_3_rs1_prfAddr : _dequeued_T_16_rs1_prfAddr; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_17_rs2_prfAddr = readyVector[3] ? queue_3_rs2_prfAddr : _dequeued_T_16_rs2_prfAddr; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_17_prfDest = readyVector[3] ? queue_3_prfDest : _dequeued_T_16_prfDest; // @[Mux.scala 101:16]
  wire [3:0] _dequeued_T_17_robAddr = readyVector[3] ? queue_3_robAddr : _dequeued_T_16_robAddr; // @[Mux.scala 101:16]
  wire  _dequeued_T_18_opcodeMeta_isM = readyVector[2] ? queue_2_opcodeMeta_isM : _dequeued_T_17_opcodeMeta_isM; // @[Mux.scala 101:16]
  wire  _dequeued_T_18_valid = readyVector[2] ? queue_2_valid : _dequeued_T_17_valid; // @[Mux.scala 101:16]
  wire [31:0] _dequeued_T_18_instruction = readyVector[2] ? queue_2_instruction : _dequeued_T_17_instruction; // @[Mux.scala 101:16]
  wire [4:0] _dequeued_T_18_branchMask = readyVector[2] ? queue_2_branchMask : _dequeued_T_17_branchMask; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_18_prfDest = readyVector[2] ? queue_2_prfDest : _dequeued_T_17_prfDest; // @[Mux.scala 101:16]
  wire  _dequeued_T_19_opcodeMeta_isM = readyVector[1] ? queue_1_opcodeMeta_isM : _dequeued_T_18_opcodeMeta_isM; // @[Mux.scala 101:16]
  wire  _dequeued_T_19_valid = readyVector[1] ? queue_1_valid : _dequeued_T_18_valid; // @[Mux.scala 101:16]
  wire [31:0] _dequeued_T_19_instruction = readyVector[1] ? queue_1_instruction : _dequeued_T_18_instruction; // @[Mux.scala 101:16]
  wire [4:0] _dequeued_T_19_branchMask = readyVector[1] ? queue_1_branchMask : _dequeued_T_18_branchMask; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_19_prfDest = readyVector[1] ? queue_1_prfDest : _dequeued_T_18_prfDest; // @[Mux.scala 101:16]
  wire  dequeued_opcodeMeta_isM = readyVector[0] ? queue_0_opcodeMeta_isM : _dequeued_T_19_opcodeMeta_isM; // @[Mux.scala 101:16]
  wire  dequeued_valid = readyVector[0] ? queue_0_valid : _dequeued_T_19_valid; // @[Mux.scala 101:16]
  wire [31:0] dequeued_instruction = readyVector[0] ? queue_0_instruction : _dequeued_T_19_instruction; // @[Mux.scala 101:16]
  wire [4:0] dequeued_branchMask = readyVector[0] ? queue_0_branchMask : _dequeued_T_19_branchMask; // @[Mux.scala 101:16]
  wire [5:0] dequeued_prfDest = readyVector[0] ? queue_0_prfDest : _dequeued_T_19_prfDest; // @[Mux.scala 101:16]
  reg  releasedBuffer_valid; // @[scheduler.scala 59:31]
  reg [31:0] releasedBuffer_instruction; // @[scheduler.scala 59:31]
  reg [4:0] releasedBuffer_branchMask; // @[scheduler.scala 59:31]
  reg [5:0] releasedBuffer_rs1prfAddr; // @[scheduler.scala 59:31]
  reg [5:0] releasedBuffer_rs2prfAddr; // @[scheduler.scala 59:31]
  reg [5:0] releasedBuffer_prfDest; // @[scheduler.scala 59:31]
  reg [3:0] releasedBuffer_robAddr; // @[scheduler.scala 59:31]
  wire  dequeue = ~releasedBuffer_valid | release_fired; // @[scheduler.scala 70:39]
  wire [4:0] _tempQueue_8_opcodeMeta_meta_isM_T_1 = allocate_instruction[6:2] & 5'h1d; // @[scheduler.scala 78:44]
  wire  tempQueue_8_opcodeMeta_meta_isM = 5'hc == _tempQueue_8_opcodeMeta_meta_isM_T_1 & allocate_instruction[25]; // @[scheduler.scala 78:66]
  wire  tempQueue_8_opcodeMeta_meta_isMemAccess = ~allocate_instruction[6] & ~allocate_instruction[4] & ~(5'h3 ==
    allocate_instruction[6:2]); // @[scheduler.scala 79:92]
  wire  tempQueue_8_opcodeMeta_meta_isBranch = allocate_instruction[6:5] == 2'h3; // @[scheduler.scala 80:48]
  wire  tempQueue_8_rs2_ready = allocate_fired & tempQueue_8_opcodeMeta_meta_isMemAccess | allocate_rs2_ready; // @[scheduler.scala 89:116 86:34 89:77]
  wire [4:0] _wakeUpInt_valid_T_1 = dequeued_instruction[6:2] & 5'h15; // @[scheduler.scala 95:49]
  wire  _wakeUpInt_valid_T_6 = |readyVector; // @[scheduler.scala 95:125]
  wire  wakeUpInt_valid = 5'h4 == _wakeUpInt_valid_T_1 & ~dequeued_opcodeMeta_isM & dequeue & |readyVector & |
    dequeued_instruction[11:7]; // @[scheduler.scala 95:129]
  wire  updatedEntries_0_rs1_ready = queue_0_valid & (queue_0_rs1_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_0_rs1_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_0_rs1_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_0_rs1_prfAddr)); // @[scheduler.scala 98:109]
  wire  updatedEntries_1_rs1_ready = queue_1_valid & (queue_1_rs1_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_1_rs1_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_1_rs1_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_1_rs1_prfAddr)); // @[scheduler.scala 98:109]
  wire  updatedEntries_2_rs1_ready = queue_2_valid & (queue_2_rs1_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_2_rs1_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_2_rs1_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_2_rs1_prfAddr)); // @[scheduler.scala 98:109]
  wire  updatedEntries_3_rs1_ready = queue_3_valid & (queue_3_rs1_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_3_rs1_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_3_rs1_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_3_rs1_prfAddr)); // @[scheduler.scala 98:109]
  wire  updatedEntries_4_rs1_ready = queue_4_valid & (queue_4_rs1_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_4_rs1_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_4_rs1_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_4_rs1_prfAddr)); // @[scheduler.scala 98:109]
  wire  updatedEntries_5_rs1_ready = queue_5_valid & (queue_5_rs1_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_5_rs1_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_5_rs1_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_5_rs1_prfAddr)); // @[scheduler.scala 98:109]
  wire  updatedEntries_6_rs1_ready = queue_6_valid & (queue_6_rs1_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_6_rs1_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_6_rs1_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_6_rs1_prfAddr)); // @[scheduler.scala 98:109]
  wire  updatedEntries_7_rs1_ready = queue_7_valid & (queue_7_rs1_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_7_rs1_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_7_rs1_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_7_rs1_prfAddr)); // @[scheduler.scala 98:109]
  wire  updatedEntries_8_rs1_ready = allocate_fired & (allocate_rs1_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    allocate_rs1_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == allocate_rs1_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == allocate_rs1_prfAddr)); // @[scheduler.scala 98:109]
  reg  instrRetired_REG_valid; // @[scheduler.scala 101:26]
  reg [5:0] instrRetired_REG_prfAddr; // @[scheduler.scala 101:26]
  wire  updatedEntries_0_rs2_ready = queue_0_valid & (queue_0_rs2_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_0_rs2_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_0_rs2_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_0_rs2_prfAddr)); // @[scheduler.scala 104:42]
  wire  updatedEntries_1_rs2_ready = queue_1_valid & (queue_1_rs2_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_1_rs2_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_1_rs2_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_1_rs2_prfAddr)); // @[scheduler.scala 104:42]
  wire  updatedEntries_2_rs2_ready = queue_2_valid & (queue_2_rs2_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_2_rs2_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_2_rs2_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_2_rs2_prfAddr)); // @[scheduler.scala 104:42]
  wire  updatedEntries_3_rs2_ready = queue_3_valid & (queue_3_rs2_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_3_rs2_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_3_rs2_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_3_rs2_prfAddr)); // @[scheduler.scala 104:42]
  wire  updatedEntries_4_rs2_ready = queue_4_valid & (queue_4_rs2_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_4_rs2_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_4_rs2_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_4_rs2_prfAddr)); // @[scheduler.scala 104:42]
  wire  updatedEntries_5_rs2_ready = queue_5_valid & (queue_5_rs2_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_5_rs2_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_5_rs2_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_5_rs2_prfAddr)); // @[scheduler.scala 104:42]
  wire  updatedEntries_6_rs2_ready = queue_6_valid & (queue_6_rs2_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_6_rs2_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_6_rs2_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_6_rs2_prfAddr)); // @[scheduler.scala 104:42]
  wire  updatedEntries_7_rs2_ready = queue_7_valid & (queue_7_rs2_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_7_rs2_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_7_rs2_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_7_rs2_prfAddr)); // @[scheduler.scala 104:42]
  wire  updatedEntries_8_rs2_ready = allocate_fired & (tempQueue_8_rs2_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr
     == allocate_rs2_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == allocate_rs2_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == allocate_rs2_prfAddr)); // @[scheduler.scala 104:42]
  wire [4:0] _T_1 = queue_0_branchMask & branchOps_branchMask; // @[scheduler.scala 109:53]
  wire  _T_2 = |_T_1; // @[scheduler.scala 109:77]
  wire [4:0] _updatedEntries_0_branchMask_T = queue_0_branchMask ^ branchOps_branchMask; // @[scheduler.scala 109:127]
  wire  _GEN_2 = branchOps_passed & |_T_1 ? queue_0_valid : queue_0_valid & ~_T_2; // @[scheduler.scala 109:82 110:35 92:81]
  wire  _GEN_4 = branchOps_valid ? _GEN_2 : queue_0_valid; // @[scheduler.scala 108:27 92:81]
  wire [4:0] _T_4 = queue_1_branchMask & branchOps_branchMask; // @[scheduler.scala 109:53]
  wire  _T_5 = |_T_4; // @[scheduler.scala 109:77]
  wire [4:0] _updatedEntries_1_branchMask_T = queue_1_branchMask ^ branchOps_branchMask; // @[scheduler.scala 109:127]
  wire  _GEN_6 = branchOps_passed & |_T_4 ? queue_1_valid : queue_1_valid & ~_T_5; // @[scheduler.scala 109:82 110:35 92:81]
  wire  _GEN_8 = branchOps_valid ? _GEN_6 : queue_1_valid; // @[scheduler.scala 108:27 92:81]
  wire [4:0] _T_7 = queue_2_branchMask & branchOps_branchMask; // @[scheduler.scala 109:53]
  wire  _T_8 = |_T_7; // @[scheduler.scala 109:77]
  wire [4:0] _updatedEntries_2_branchMask_T = queue_2_branchMask ^ branchOps_branchMask; // @[scheduler.scala 109:127]
  wire  _GEN_10 = branchOps_passed & |_T_7 ? queue_2_valid : queue_2_valid & ~_T_8; // @[scheduler.scala 109:82 110:35 92:81]
  wire  _GEN_12 = branchOps_valid ? _GEN_10 : queue_2_valid; // @[scheduler.scala 108:27 92:81]
  wire [4:0] _T_10 = queue_3_branchMask & branchOps_branchMask; // @[scheduler.scala 109:53]
  wire  _T_11 = |_T_10; // @[scheduler.scala 109:77]
  wire [4:0] _updatedEntries_3_branchMask_T = queue_3_branchMask ^ branchOps_branchMask; // @[scheduler.scala 109:127]
  wire  _GEN_14 = branchOps_passed & |_T_10 ? queue_3_valid : queue_3_valid & ~_T_11; // @[scheduler.scala 109:82 110:35 92:81]
  wire  _GEN_16 = branchOps_valid ? _GEN_14 : queue_3_valid; // @[scheduler.scala 108:27 92:81]
  wire [4:0] _T_13 = queue_4_branchMask & branchOps_branchMask; // @[scheduler.scala 109:53]
  wire  _T_14 = |_T_13; // @[scheduler.scala 109:77]
  wire [4:0] _updatedEntries_4_branchMask_T = queue_4_branchMask ^ branchOps_branchMask; // @[scheduler.scala 109:127]
  wire  _GEN_18 = branchOps_passed & |_T_13 ? queue_4_valid : queue_4_valid & ~_T_14; // @[scheduler.scala 109:82 110:35 92:81]
  wire  _GEN_20 = branchOps_valid ? _GEN_18 : queue_4_valid; // @[scheduler.scala 108:27 92:81]
  wire [4:0] _T_16 = queue_5_branchMask & branchOps_branchMask; // @[scheduler.scala 109:53]
  wire  _T_17 = |_T_16; // @[scheduler.scala 109:77]
  wire [4:0] _updatedEntries_5_branchMask_T = queue_5_branchMask ^ branchOps_branchMask; // @[scheduler.scala 109:127]
  wire  _GEN_22 = branchOps_passed & |_T_16 ? queue_5_valid : queue_5_valid & ~_T_17; // @[scheduler.scala 109:82 110:35 92:81]
  wire  _GEN_24 = branchOps_valid ? _GEN_22 : queue_5_valid; // @[scheduler.scala 108:27 92:81]
  wire [4:0] _T_19 = queue_6_branchMask & branchOps_branchMask; // @[scheduler.scala 109:53]
  wire  _T_20 = |_T_19; // @[scheduler.scala 109:77]
  wire [4:0] _updatedEntries_6_branchMask_T = queue_6_branchMask ^ branchOps_branchMask; // @[scheduler.scala 109:127]
  wire  _GEN_26 = branchOps_passed & |_T_19 ? queue_6_valid : queue_6_valid & ~_T_20; // @[scheduler.scala 109:82 110:35 92:81]
  wire  _GEN_28 = branchOps_valid ? _GEN_26 : queue_6_valid; // @[scheduler.scala 108:27 92:81]
  wire [4:0] _T_22 = queue_7_branchMask & branchOps_branchMask; // @[scheduler.scala 109:53]
  wire  _T_23 = |_T_22; // @[scheduler.scala 109:77]
  wire [4:0] _updatedEntries_7_branchMask_T = queue_7_branchMask ^ branchOps_branchMask; // @[scheduler.scala 109:127]
  wire  _GEN_30 = branchOps_passed & |_T_22 ? queue_7_valid : queue_7_valid & ~_T_23; // @[scheduler.scala 109:82 110:35 92:81]
  wire  _GEN_32 = branchOps_valid ? _GEN_30 : queue_7_valid; // @[scheduler.scala 108:27 92:81]
  wire [4:0] _T_25 = allocate_branchMask & branchOps_branchMask; // @[scheduler.scala 109:53]
  wire  _T_26 = |_T_25; // @[scheduler.scala 109:77]
  wire [4:0] _updatedEntries_8_branchMask_T = allocate_branchMask ^ branchOps_branchMask; // @[scheduler.scala 109:127]
  wire  _T_29 = dequeue & _wakeUpInt_valid_T_6; // @[scheduler.scala 114:16]
  wire  _newQueue_T_69 = queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid
     & queue_6_valid & queue_7_valid; // @[scheduler.scala 116:110]
  wire [4:0] _releasedBuffer_branchMask_T = branchOps_branchMask & dequeued_branchMask; // @[scheduler.scala 137:79]
  wire [4:0] _releasedBuffer_branchMask_T_4 = dequeued_branchMask ^ branchOps_branchMask; // @[scheduler.scala 137:147]
  wire  _releasedBuffer_valid_T = ~branchOps_valid; // @[scheduler.scala 143:48]
  wire [4:0] _releasedBuffer_valid_T_1 = dequeued_branchMask & branchOps_branchMask; // @[scheduler.scala 143:90]
  wire [4:0] _releasedBuffer_branchMask_T_6 = releasedBuffer_branchMask ^ branchOps_branchMask; // @[scheduler.scala 145:60]
  wire [4:0] _releasedBuffer_valid_T_10 = releasedBuffer_branchMask & branchOps_branchMask; // @[scheduler.scala 146:102]
  assign allocate_ready = ~_newQueue_T_69; // @[scheduler.scala 134:21]
  assign release_ready = releasedBuffer_valid; // @[scheduler.scala 133:17]
  assign release_instruction = releasedBuffer_instruction; // @[scheduler.scala 128:23]
  assign release_branchMask = releasedBuffer_branchMask; // @[scheduler.scala 127:22]
  assign release_rs1prfAddr = releasedBuffer_rs1prfAddr; // @[scheduler.scala 131:22]
  assign release_rs2prfAddr = releasedBuffer_rs2prfAddr; // @[scheduler.scala 132:22]
  assign release_prfDest = releasedBuffer_prfDest; // @[scheduler.scala 129:19]
  assign release_robAddr = releasedBuffer_robAddr; // @[scheduler.scala 130:19]
  assign instrRetired_valid = instrRetired_REG_valid; // @[scheduler.scala 101:16]
  assign instrRetired_prfAddr = instrRetired_REG_prfAddr; // @[scheduler.scala 101:16]
  always @(posedge clock) begin
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_opcodeMeta_isBranch <= queue_1_opcodeMeta_isBranch;
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_opcodeMeta_isMemAccess <= queue_1_opcodeMeta_isMemAccess;
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_opcodeMeta_isM <= queue_1_opcodeMeta_isM;
    end
    if (reset) begin // @[scheduler.scala 26:22]
      queue_0_valid <= 1'h0; // @[scheduler.scala 26:22]
    end else if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
        if (3'h1 == dequeuedIndex) begin // @[scheduler.scala 114:106]
          queue_0_valid <= 1'h0; // @[scheduler.scala 114:132]
        end else begin
          queue_0_valid <= _GEN_8;
        end
      end else begin
        queue_0_valid <= _GEN_8;
      end
    end else if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
      if (3'h0 == dequeuedIndex) begin // @[scheduler.scala 114:106]
        queue_0_valid <= 1'h0; // @[scheduler.scala 114:132]
      end else begin
        queue_0_valid <= _GEN_4;
      end
    end else begin
      queue_0_valid <= _GEN_4;
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_instruction <= queue_1_instruction;
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      if (branchOps_valid) begin // @[scheduler.scala 108:27]
        if (branchOps_passed & |_T_4) begin // @[scheduler.scala 109:82]
          queue_0_branchMask <= _updatedEntries_1_branchMask_T; // @[scheduler.scala 109:104]
        end else begin
          queue_0_branchMask <= queue_1_branchMask; // @[scheduler.scala 92:81]
        end
      end else begin
        queue_0_branchMask <= queue_1_branchMask; // @[scheduler.scala 92:81]
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 108:27]
      if (branchOps_passed & |_T_1) begin // @[scheduler.scala 109:82]
        queue_0_branchMask <= _updatedEntries_0_branchMask_T; // @[scheduler.scala 109:104]
      end
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_rs1_ready <= updatedEntries_1_rs1_ready;
    end else begin
      queue_0_rs1_ready <= updatedEntries_0_rs1_ready;
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_rs1_prfAddr <= queue_1_rs1_prfAddr;
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_rs2_ready <= updatedEntries_1_rs2_ready;
    end else begin
      queue_0_rs2_ready <= updatedEntries_0_rs2_ready;
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_rs2_prfAddr <= queue_1_rs2_prfAddr;
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_prfDest <= queue_1_prfDest;
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_robAddr <= queue_1_robAddr;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_opcodeMeta_isBranch <= queue_2_opcodeMeta_isBranch;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_opcodeMeta_isMemAccess <= queue_2_opcodeMeta_isMemAccess;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_opcodeMeta_isM <= queue_2_opcodeMeta_isM;
    end
    if (reset) begin // @[scheduler.scala 26:22]
      queue_1_valid <= 1'h0; // @[scheduler.scala 26:22]
    end else if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
        if (3'h2 == dequeuedIndex) begin // @[scheduler.scala 114:106]
          queue_1_valid <= 1'h0; // @[scheduler.scala 114:132]
        end else begin
          queue_1_valid <= _GEN_12;
        end
      end else begin
        queue_1_valid <= _GEN_12;
      end
    end else if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
      if (3'h1 == dequeuedIndex) begin // @[scheduler.scala 114:106]
        queue_1_valid <= 1'h0; // @[scheduler.scala 114:132]
      end else begin
        queue_1_valid <= _GEN_8;
      end
    end else begin
      queue_1_valid <= _GEN_8;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_instruction <= queue_2_instruction;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      if (branchOps_valid) begin // @[scheduler.scala 108:27]
        if (branchOps_passed & |_T_7) begin // @[scheduler.scala 109:82]
          queue_1_branchMask <= _updatedEntries_2_branchMask_T; // @[scheduler.scala 109:104]
        end else begin
          queue_1_branchMask <= queue_2_branchMask; // @[scheduler.scala 92:81]
        end
      end else begin
        queue_1_branchMask <= queue_2_branchMask; // @[scheduler.scala 92:81]
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 108:27]
      if (branchOps_passed & |_T_4) begin // @[scheduler.scala 109:82]
        queue_1_branchMask <= _updatedEntries_1_branchMask_T; // @[scheduler.scala 109:104]
      end
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_rs1_ready <= updatedEntries_2_rs1_ready;
    end else begin
      queue_1_rs1_ready <= updatedEntries_1_rs1_ready;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_rs1_prfAddr <= queue_2_rs1_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_rs2_ready <= updatedEntries_2_rs2_ready;
    end else begin
      queue_1_rs2_ready <= updatedEntries_1_rs2_ready;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_rs2_prfAddr <= queue_2_rs2_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_prfDest <= queue_2_prfDest;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_robAddr <= queue_2_robAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_opcodeMeta_isBranch <= queue_3_opcodeMeta_isBranch;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_opcodeMeta_isMemAccess <= queue_3_opcodeMeta_isMemAccess;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_opcodeMeta_isM <= queue_3_opcodeMeta_isM;
    end
    if (reset) begin // @[scheduler.scala 26:22]
      queue_2_valid <= 1'h0; // @[scheduler.scala 26:22]
    end else if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
        if (3'h3 == dequeuedIndex) begin // @[scheduler.scala 114:106]
          queue_2_valid <= 1'h0; // @[scheduler.scala 114:132]
        end else begin
          queue_2_valid <= _GEN_16;
        end
      end else begin
        queue_2_valid <= _GEN_16;
      end
    end else if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
      if (3'h2 == dequeuedIndex) begin // @[scheduler.scala 114:106]
        queue_2_valid <= 1'h0; // @[scheduler.scala 114:132]
      end else begin
        queue_2_valid <= _GEN_12;
      end
    end else begin
      queue_2_valid <= _GEN_12;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_instruction <= queue_3_instruction;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      if (branchOps_valid) begin // @[scheduler.scala 108:27]
        if (branchOps_passed & |_T_10) begin // @[scheduler.scala 109:82]
          queue_2_branchMask <= _updatedEntries_3_branchMask_T; // @[scheduler.scala 109:104]
        end else begin
          queue_2_branchMask <= queue_3_branchMask; // @[scheduler.scala 92:81]
        end
      end else begin
        queue_2_branchMask <= queue_3_branchMask; // @[scheduler.scala 92:81]
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 108:27]
      if (branchOps_passed & |_T_7) begin // @[scheduler.scala 109:82]
        queue_2_branchMask <= _updatedEntries_2_branchMask_T; // @[scheduler.scala 109:104]
      end
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_rs1_ready <= updatedEntries_3_rs1_ready;
    end else begin
      queue_2_rs1_ready <= updatedEntries_2_rs1_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_rs1_prfAddr <= queue_3_rs1_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_rs2_ready <= updatedEntries_3_rs2_ready;
    end else begin
      queue_2_rs2_ready <= updatedEntries_2_rs2_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_rs2_prfAddr <= queue_3_rs2_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_prfDest <= queue_3_prfDest;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_robAddr <= queue_3_robAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_opcodeMeta_isBranch <= queue_4_opcodeMeta_isBranch;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_opcodeMeta_isMemAccess <= queue_4_opcodeMeta_isMemAccess;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_opcodeMeta_isM <= queue_4_opcodeMeta_isM;
    end
    if (reset) begin // @[scheduler.scala 26:22]
      queue_3_valid <= 1'h0; // @[scheduler.scala 26:22]
    end else if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
        if (3'h4 == dequeuedIndex) begin // @[scheduler.scala 114:106]
          queue_3_valid <= 1'h0; // @[scheduler.scala 114:132]
        end else begin
          queue_3_valid <= _GEN_20;
        end
      end else begin
        queue_3_valid <= _GEN_20;
      end
    end else if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
      if (3'h3 == dequeuedIndex) begin // @[scheduler.scala 114:106]
        queue_3_valid <= 1'h0; // @[scheduler.scala 114:132]
      end else begin
        queue_3_valid <= _GEN_16;
      end
    end else begin
      queue_3_valid <= _GEN_16;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_instruction <= queue_4_instruction;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      if (branchOps_valid) begin // @[scheduler.scala 108:27]
        if (branchOps_passed & |_T_13) begin // @[scheduler.scala 109:82]
          queue_3_branchMask <= _updatedEntries_4_branchMask_T; // @[scheduler.scala 109:104]
        end else begin
          queue_3_branchMask <= queue_4_branchMask; // @[scheduler.scala 92:81]
        end
      end else begin
        queue_3_branchMask <= queue_4_branchMask; // @[scheduler.scala 92:81]
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 108:27]
      if (branchOps_passed & |_T_10) begin // @[scheduler.scala 109:82]
        queue_3_branchMask <= _updatedEntries_3_branchMask_T; // @[scheduler.scala 109:104]
      end
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_rs1_ready <= updatedEntries_4_rs1_ready;
    end else begin
      queue_3_rs1_ready <= updatedEntries_3_rs1_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_rs1_prfAddr <= queue_4_rs1_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_rs2_ready <= updatedEntries_4_rs2_ready;
    end else begin
      queue_3_rs2_ready <= updatedEntries_3_rs2_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_rs2_prfAddr <= queue_4_rs2_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_prfDest <= queue_4_prfDest;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_robAddr <= queue_4_robAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_opcodeMeta_isBranch <= queue_5_opcodeMeta_isBranch;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_opcodeMeta_isMemAccess <= queue_5_opcodeMeta_isMemAccess;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_opcodeMeta_isM <= queue_5_opcodeMeta_isM;
    end
    if (reset) begin // @[scheduler.scala 26:22]
      queue_4_valid <= 1'h0; // @[scheduler.scala 26:22]
    end else if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |
      readyVector[4:0]) begin // @[scheduler.scala 116:60]
      if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
        if (3'h5 == dequeuedIndex) begin // @[scheduler.scala 114:106]
          queue_4_valid <= 1'h0; // @[scheduler.scala 114:132]
        end else begin
          queue_4_valid <= _GEN_24;
        end
      end else begin
        queue_4_valid <= _GEN_24;
      end
    end else if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
      if (3'h4 == dequeuedIndex) begin // @[scheduler.scala 114:106]
        queue_4_valid <= 1'h0; // @[scheduler.scala 114:132]
      end else begin
        queue_4_valid <= _GEN_20;
      end
    end else begin
      queue_4_valid <= _GEN_20;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_instruction <= queue_5_instruction;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      if (branchOps_valid) begin // @[scheduler.scala 108:27]
        if (branchOps_passed & |_T_16) begin // @[scheduler.scala 109:82]
          queue_4_branchMask <= _updatedEntries_5_branchMask_T; // @[scheduler.scala 109:104]
        end else begin
          queue_4_branchMask <= queue_5_branchMask; // @[scheduler.scala 92:81]
        end
      end else begin
        queue_4_branchMask <= queue_5_branchMask; // @[scheduler.scala 92:81]
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 108:27]
      if (branchOps_passed & |_T_13) begin // @[scheduler.scala 109:82]
        queue_4_branchMask <= _updatedEntries_4_branchMask_T; // @[scheduler.scala 109:104]
      end
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_rs1_ready <= updatedEntries_5_rs1_ready;
    end else begin
      queue_4_rs1_ready <= updatedEntries_4_rs1_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_rs1_prfAddr <= queue_5_rs1_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_rs2_ready <= updatedEntries_5_rs2_ready;
    end else begin
      queue_4_rs2_ready <= updatedEntries_4_rs2_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_rs2_prfAddr <= queue_5_rs2_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_prfDest <= queue_5_prfDest;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_robAddr <= queue_5_robAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_opcodeMeta_isBranch <= queue_6_opcodeMeta_isBranch;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_opcodeMeta_isMemAccess <= queue_6_opcodeMeta_isMemAccess;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_opcodeMeta_isM <= queue_6_opcodeMeta_isM;
    end
    if (reset) begin // @[scheduler.scala 26:22]
      queue_5_valid <= 1'h0; // @[scheduler.scala 26:22]
    end else if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) |
      dequeue & |readyVector[5:0]) begin // @[scheduler.scala 116:60]
      if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
        if (3'h6 == dequeuedIndex) begin // @[scheduler.scala 114:106]
          queue_5_valid <= 1'h0; // @[scheduler.scala 114:132]
        end else begin
          queue_5_valid <= _GEN_28;
        end
      end else begin
        queue_5_valid <= _GEN_28;
      end
    end else if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
      if (3'h5 == dequeuedIndex) begin // @[scheduler.scala 114:106]
        queue_5_valid <= 1'h0; // @[scheduler.scala 114:132]
      end else begin
        queue_5_valid <= _GEN_24;
      end
    end else begin
      queue_5_valid <= _GEN_24;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_instruction <= queue_6_instruction;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      if (branchOps_valid) begin // @[scheduler.scala 108:27]
        if (branchOps_passed & |_T_19) begin // @[scheduler.scala 109:82]
          queue_5_branchMask <= _updatedEntries_6_branchMask_T; // @[scheduler.scala 109:104]
        end else begin
          queue_5_branchMask <= queue_6_branchMask; // @[scheduler.scala 92:81]
        end
      end else begin
        queue_5_branchMask <= queue_6_branchMask; // @[scheduler.scala 92:81]
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 108:27]
      if (branchOps_passed & |_T_16) begin // @[scheduler.scala 109:82]
        queue_5_branchMask <= _updatedEntries_5_branchMask_T; // @[scheduler.scala 109:104]
      end
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_rs1_ready <= updatedEntries_6_rs1_ready;
    end else begin
      queue_5_rs1_ready <= updatedEntries_5_rs1_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_rs1_prfAddr <= queue_6_rs1_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_rs2_ready <= updatedEntries_6_rs2_ready;
    end else begin
      queue_5_rs2_ready <= updatedEntries_5_rs2_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_rs2_prfAddr <= queue_6_rs2_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_prfDest <= queue_6_prfDest;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_robAddr <= queue_6_robAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_opcodeMeta_isBranch <= queue_7_opcodeMeta_isBranch;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_opcodeMeta_isMemAccess <= queue_7_opcodeMeta_isMemAccess;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_opcodeMeta_isM <= queue_7_opcodeMeta_isM;
    end
    if (reset) begin // @[scheduler.scala 26:22]
      queue_6_valid <= 1'h0; // @[scheduler.scala 26:22]
    end else if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid &
      queue_6_valid) | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
        if (3'h7 == dequeuedIndex) begin // @[scheduler.scala 114:106]
          queue_6_valid <= 1'h0; // @[scheduler.scala 114:132]
        end else begin
          queue_6_valid <= _GEN_32;
        end
      end else begin
        queue_6_valid <= _GEN_32;
      end
    end else if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
      if (3'h6 == dequeuedIndex) begin // @[scheduler.scala 114:106]
        queue_6_valid <= 1'h0; // @[scheduler.scala 114:132]
      end else begin
        queue_6_valid <= _GEN_28;
      end
    end else begin
      queue_6_valid <= _GEN_28;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_instruction <= queue_7_instruction;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      if (branchOps_valid) begin // @[scheduler.scala 108:27]
        if (branchOps_passed & |_T_22) begin // @[scheduler.scala 109:82]
          queue_6_branchMask <= _updatedEntries_7_branchMask_T; // @[scheduler.scala 109:104]
        end else begin
          queue_6_branchMask <= queue_7_branchMask; // @[scheduler.scala 92:81]
        end
      end else begin
        queue_6_branchMask <= queue_7_branchMask; // @[scheduler.scala 92:81]
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 108:27]
      if (branchOps_passed & |_T_19) begin // @[scheduler.scala 109:82]
        queue_6_branchMask <= _updatedEntries_6_branchMask_T; // @[scheduler.scala 109:104]
      end
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_rs1_ready <= updatedEntries_7_rs1_ready;
    end else begin
      queue_6_rs1_ready <= updatedEntries_6_rs1_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_rs1_prfAddr <= queue_7_rs1_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_rs2_ready <= updatedEntries_7_rs2_ready;
    end else begin
      queue_6_rs2_ready <= updatedEntries_6_rs2_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_rs2_prfAddr <= queue_7_rs2_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_prfDest <= queue_7_prfDest;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_robAddr <= queue_7_robAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_opcodeMeta_isBranch <= tempQueue_8_opcodeMeta_meta_isBranch;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_opcodeMeta_isMemAccess <= tempQueue_8_opcodeMeta_meta_isMemAccess;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_opcodeMeta_isM <= tempQueue_8_opcodeMeta_meta_isM;
    end
    if (reset) begin // @[scheduler.scala 26:22]
      queue_7_valid <= 1'h0; // @[scheduler.scala 26:22]
    end else if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid &
      queue_6_valid & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      if (branchOps_valid) begin // @[scheduler.scala 108:27]
        if (branchOps_passed & |_T_25) begin // @[scheduler.scala 109:82]
          queue_7_valid <= allocate_fired; // @[scheduler.scala 92:81]
        end else begin
          queue_7_valid <= allocate_fired & ~_T_26; // @[scheduler.scala 110:35]
        end
      end else begin
        queue_7_valid <= allocate_fired; // @[scheduler.scala 92:81]
      end
    end else if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
      if (3'h7 == dequeuedIndex) begin // @[scheduler.scala 114:106]
        queue_7_valid <= 1'h0; // @[scheduler.scala 114:132]
      end else begin
        queue_7_valid <= _GEN_32;
      end
    end else begin
      queue_7_valid <= _GEN_32;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_instruction <= allocate_instruction;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      if (branchOps_valid) begin // @[scheduler.scala 108:27]
        if (branchOps_passed & |_T_25) begin // @[scheduler.scala 109:82]
          queue_7_branchMask <= _updatedEntries_8_branchMask_T; // @[scheduler.scala 109:104]
        end else begin
          queue_7_branchMask <= allocate_branchMask; // @[scheduler.scala 92:81]
        end
      end else begin
        queue_7_branchMask <= allocate_branchMask; // @[scheduler.scala 92:81]
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 108:27]
      if (branchOps_passed & |_T_22) begin // @[scheduler.scala 109:82]
        queue_7_branchMask <= _updatedEntries_7_branchMask_T; // @[scheduler.scala 109:104]
      end
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_rs1_ready <= updatedEntries_8_rs1_ready;
    end else begin
      queue_7_rs1_ready <= updatedEntries_7_rs1_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_rs1_prfAddr <= allocate_rs1_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_rs2_ready <= updatedEntries_8_rs2_ready;
    end else begin
      queue_7_rs2_ready <= updatedEntries_7_rs2_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_rs2_prfAddr <= allocate_rs2_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_prfDest <= allocate_prfDest;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_robAddr <= allocate_robAddr;
    end
    if (reset) begin // @[scheduler.scala 59:31]
      releasedBuffer_valid <= 1'h0; // @[scheduler.scala 59:31]
    end else if (dequeue) begin // @[scheduler.scala 136:17]
      releasedBuffer_valid <= dequeued_valid & (~branchOps_valid | ~(|_releasedBuffer_valid_T_1) | branchOps_passed) &
        _wakeUpInt_valid_T_6; // @[scheduler.scala 143:26]
    end else if (branchOps_valid) begin // @[scheduler.scala 144:31]
      releasedBuffer_valid <= releasedBuffer_valid & (_releasedBuffer_valid_T | ~(|_releasedBuffer_valid_T_10) |
        branchOps_passed); // @[scheduler.scala 146:26]
    end
    if (dequeue) begin // @[scheduler.scala 136:17]
      if (readyVector[0]) begin // @[Mux.scala 101:16]
        releasedBuffer_instruction <= queue_0_instruction;
      end else if (readyVector[1]) begin // @[Mux.scala 101:16]
        releasedBuffer_instruction <= queue_1_instruction;
      end else if (readyVector[2]) begin // @[Mux.scala 101:16]
        releasedBuffer_instruction <= queue_2_instruction;
      end else begin
        releasedBuffer_instruction <= _dequeued_T_17_instruction;
      end
    end
    if (dequeue) begin // @[scheduler.scala 136:17]
      if (branchOps_valid & |_releasedBuffer_branchMask_T & branchOps_passed) begin // @[scheduler.scala 137:37]
        releasedBuffer_branchMask <= _releasedBuffer_branchMask_T_4;
      end else if (readyVector[0]) begin // @[Mux.scala 101:16]
        releasedBuffer_branchMask <= queue_0_branchMask;
      end else if (readyVector[1]) begin // @[Mux.scala 101:16]
        releasedBuffer_branchMask <= queue_1_branchMask;
      end else begin
        releasedBuffer_branchMask <= _dequeued_T_18_branchMask;
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 144:31]
      releasedBuffer_branchMask <= _releasedBuffer_branchMask_T_6; // @[scheduler.scala 145:31]
    end
    if (dequeue) begin // @[scheduler.scala 136:17]
      if (readyVector[0]) begin // @[Mux.scala 101:16]
        releasedBuffer_rs1prfAddr <= queue_0_rs1_prfAddr;
      end else if (readyVector[1]) begin // @[Mux.scala 101:16]
        releasedBuffer_rs1prfAddr <= queue_1_rs1_prfAddr;
      end else if (readyVector[2]) begin // @[Mux.scala 101:16]
        releasedBuffer_rs1prfAddr <= queue_2_rs1_prfAddr;
      end else begin
        releasedBuffer_rs1prfAddr <= _dequeued_T_17_rs1_prfAddr;
      end
    end
    if (dequeue) begin // @[scheduler.scala 136:17]
      if (readyVector[0]) begin // @[Mux.scala 101:16]
        releasedBuffer_rs2prfAddr <= queue_0_rs2_prfAddr;
      end else if (readyVector[1]) begin // @[Mux.scala 101:16]
        releasedBuffer_rs2prfAddr <= queue_1_rs2_prfAddr;
      end else if (readyVector[2]) begin // @[Mux.scala 101:16]
        releasedBuffer_rs2prfAddr <= queue_2_rs2_prfAddr;
      end else begin
        releasedBuffer_rs2prfAddr <= _dequeued_T_17_rs2_prfAddr;
      end
    end
    if (dequeue) begin // @[scheduler.scala 136:17]
      if (readyVector[0]) begin // @[Mux.scala 101:16]
        releasedBuffer_prfDest <= queue_0_prfDest;
      end else if (readyVector[1]) begin // @[Mux.scala 101:16]
        releasedBuffer_prfDest <= queue_1_prfDest;
      end else if (readyVector[2]) begin // @[Mux.scala 101:16]
        releasedBuffer_prfDest <= queue_2_prfDest;
      end else begin
        releasedBuffer_prfDest <= _dequeued_T_17_prfDest;
      end
    end
    if (dequeue) begin // @[scheduler.scala 136:17]
      if (readyVector[0]) begin // @[Mux.scala 101:16]
        releasedBuffer_robAddr <= queue_0_robAddr;
      end else if (readyVector[1]) begin // @[Mux.scala 101:16]
        releasedBuffer_robAddr <= queue_1_robAddr;
      end else if (readyVector[2]) begin // @[Mux.scala 101:16]
        releasedBuffer_robAddr <= queue_2_robAddr;
      end else begin
        releasedBuffer_robAddr <= _dequeued_T_17_robAddr;
      end
    end
    instrRetired_REG_valid <= 5'h4 == _wakeUpInt_valid_T_1 & ~dequeued_opcodeMeta_isM & dequeue & |readyVector & |
      dequeued_instruction[11:7]; // @[scheduler.scala 95:129]
    if (readyVector[0]) begin // @[Mux.scala 101:16]
      instrRetired_REG_prfAddr <= queue_0_prfDest;
    end else if (readyVector[1]) begin // @[Mux.scala 101:16]
      instrRetired_REG_prfAddr <= queue_1_prfDest;
    end else if (readyVector[2]) begin // @[Mux.scala 101:16]
      instrRetired_REG_prfAddr <= queue_2_prfDest;
    end else if (readyVector[3]) begin // @[Mux.scala 101:16]
      instrRetired_REG_prfAddr <= queue_3_prfDest;
    end else begin
      instrRetired_REG_prfAddr <= _dequeued_T_16_prfDest;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  queue_0_opcodeMeta_isBranch = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  queue_0_opcodeMeta_isMemAccess = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  queue_0_opcodeMeta_isM = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  queue_0_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  queue_0_instruction = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  queue_0_branchMask = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  queue_0_rs1_ready = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  queue_0_rs1_prfAddr = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  queue_0_rs2_ready = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  queue_0_rs2_prfAddr = _RAND_9[5:0];
  _RAND_10 = {1{`RANDOM}};
  queue_0_prfDest = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  queue_0_robAddr = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  queue_1_opcodeMeta_isBranch = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  queue_1_opcodeMeta_isMemAccess = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  queue_1_opcodeMeta_isM = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  queue_1_valid = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  queue_1_instruction = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  queue_1_branchMask = _RAND_17[4:0];
  _RAND_18 = {1{`RANDOM}};
  queue_1_rs1_ready = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  queue_1_rs1_prfAddr = _RAND_19[5:0];
  _RAND_20 = {1{`RANDOM}};
  queue_1_rs2_ready = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  queue_1_rs2_prfAddr = _RAND_21[5:0];
  _RAND_22 = {1{`RANDOM}};
  queue_1_prfDest = _RAND_22[5:0];
  _RAND_23 = {1{`RANDOM}};
  queue_1_robAddr = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  queue_2_opcodeMeta_isBranch = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  queue_2_opcodeMeta_isMemAccess = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  queue_2_opcodeMeta_isM = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  queue_2_valid = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  queue_2_instruction = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  queue_2_branchMask = _RAND_29[4:0];
  _RAND_30 = {1{`RANDOM}};
  queue_2_rs1_ready = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  queue_2_rs1_prfAddr = _RAND_31[5:0];
  _RAND_32 = {1{`RANDOM}};
  queue_2_rs2_ready = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  queue_2_rs2_prfAddr = _RAND_33[5:0];
  _RAND_34 = {1{`RANDOM}};
  queue_2_prfDest = _RAND_34[5:0];
  _RAND_35 = {1{`RANDOM}};
  queue_2_robAddr = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  queue_3_opcodeMeta_isBranch = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  queue_3_opcodeMeta_isMemAccess = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  queue_3_opcodeMeta_isM = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  queue_3_valid = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  queue_3_instruction = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  queue_3_branchMask = _RAND_41[4:0];
  _RAND_42 = {1{`RANDOM}};
  queue_3_rs1_ready = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  queue_3_rs1_prfAddr = _RAND_43[5:0];
  _RAND_44 = {1{`RANDOM}};
  queue_3_rs2_ready = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  queue_3_rs2_prfAddr = _RAND_45[5:0];
  _RAND_46 = {1{`RANDOM}};
  queue_3_prfDest = _RAND_46[5:0];
  _RAND_47 = {1{`RANDOM}};
  queue_3_robAddr = _RAND_47[3:0];
  _RAND_48 = {1{`RANDOM}};
  queue_4_opcodeMeta_isBranch = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  queue_4_opcodeMeta_isMemAccess = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  queue_4_opcodeMeta_isM = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  queue_4_valid = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  queue_4_instruction = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  queue_4_branchMask = _RAND_53[4:0];
  _RAND_54 = {1{`RANDOM}};
  queue_4_rs1_ready = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  queue_4_rs1_prfAddr = _RAND_55[5:0];
  _RAND_56 = {1{`RANDOM}};
  queue_4_rs2_ready = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  queue_4_rs2_prfAddr = _RAND_57[5:0];
  _RAND_58 = {1{`RANDOM}};
  queue_4_prfDest = _RAND_58[5:0];
  _RAND_59 = {1{`RANDOM}};
  queue_4_robAddr = _RAND_59[3:0];
  _RAND_60 = {1{`RANDOM}};
  queue_5_opcodeMeta_isBranch = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  queue_5_opcodeMeta_isMemAccess = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  queue_5_opcodeMeta_isM = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  queue_5_valid = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  queue_5_instruction = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  queue_5_branchMask = _RAND_65[4:0];
  _RAND_66 = {1{`RANDOM}};
  queue_5_rs1_ready = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  queue_5_rs1_prfAddr = _RAND_67[5:0];
  _RAND_68 = {1{`RANDOM}};
  queue_5_rs2_ready = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  queue_5_rs2_prfAddr = _RAND_69[5:0];
  _RAND_70 = {1{`RANDOM}};
  queue_5_prfDest = _RAND_70[5:0];
  _RAND_71 = {1{`RANDOM}};
  queue_5_robAddr = _RAND_71[3:0];
  _RAND_72 = {1{`RANDOM}};
  queue_6_opcodeMeta_isBranch = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  queue_6_opcodeMeta_isMemAccess = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  queue_6_opcodeMeta_isM = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  queue_6_valid = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  queue_6_instruction = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  queue_6_branchMask = _RAND_77[4:0];
  _RAND_78 = {1{`RANDOM}};
  queue_6_rs1_ready = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  queue_6_rs1_prfAddr = _RAND_79[5:0];
  _RAND_80 = {1{`RANDOM}};
  queue_6_rs2_ready = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  queue_6_rs2_prfAddr = _RAND_81[5:0];
  _RAND_82 = {1{`RANDOM}};
  queue_6_prfDest = _RAND_82[5:0];
  _RAND_83 = {1{`RANDOM}};
  queue_6_robAddr = _RAND_83[3:0];
  _RAND_84 = {1{`RANDOM}};
  queue_7_opcodeMeta_isBranch = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  queue_7_opcodeMeta_isMemAccess = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  queue_7_opcodeMeta_isM = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  queue_7_valid = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  queue_7_instruction = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  queue_7_branchMask = _RAND_89[4:0];
  _RAND_90 = {1{`RANDOM}};
  queue_7_rs1_ready = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  queue_7_rs1_prfAddr = _RAND_91[5:0];
  _RAND_92 = {1{`RANDOM}};
  queue_7_rs2_ready = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  queue_7_rs2_prfAddr = _RAND_93[5:0];
  _RAND_94 = {1{`RANDOM}};
  queue_7_prfDest = _RAND_94[5:0];
  _RAND_95 = {1{`RANDOM}};
  queue_7_robAddr = _RAND_95[3:0];
  _RAND_96 = {1{`RANDOM}};
  releasedBuffer_valid = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  releasedBuffer_instruction = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  releasedBuffer_branchMask = _RAND_98[4:0];
  _RAND_99 = {1{`RANDOM}};
  releasedBuffer_rs1prfAddr = _RAND_99[5:0];
  _RAND_100 = {1{`RANDOM}};
  releasedBuffer_rs2prfAddr = _RAND_100[5:0];
  _RAND_101 = {1{`RANDOM}};
  releasedBuffer_prfDest = _RAND_101[5:0];
  _RAND_102 = {1{`RANDOM}};
  releasedBuffer_robAddr = _RAND_102[3:0];
  _RAND_103 = {1{`RANDOM}};
  instrRetired_REG_valid = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  instrRetired_REG_prfAddr = _RAND_104[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module fifoWithAddrCheck(
  input         clock,
  input         reset,
  output        write_ready,
  input         write_data_valid,
  input  [31:0] write_data_address,
  input  [31:0] write_data_core_instruction,
  input  [3:0]  write_data_core_robAddr,
  input  [5:0]  write_data_core_prfDest,
  input         write_data_branch_valid,
  input  [4:0]  write_data_branch_mask,
  input         read_ready,
  output        read_data_valid,
  output [31:0] read_data_address,
  output [31:0] read_data_core_instruction,
  output [3:0]  read_data_core_robAddr,
  output [5:0]  read_data_core_prfDest,
  output        read_data_branch_valid,
  output [4:0]  read_data_branch_mask,
  output        isEmpty,
  input         branchOps_valid,
  input  [4:0]  branchOps_branchMask,
  input         branchOps_passed,
  input  [31:0] checkAddress,
  output        matchFound
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
`endif // RANDOMIZE_REG_INIT
  reg  memReg_0_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_0_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_0_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_0_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_0_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_0_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_0_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_1_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_1_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_1_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_1_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_1_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_1_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_1_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_2_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_2_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_2_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_2_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_2_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_2_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_2_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_3_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_3_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_3_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_3_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_3_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_3_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_3_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_4_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_4_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_4_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_4_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_4_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_4_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_4_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_5_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_5_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_5_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_5_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_5_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_5_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_5_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_6_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_6_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_6_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_6_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_6_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_6_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_6_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_7_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_7_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_7_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_7_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_7_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_7_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_7_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_8_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_8_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_8_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_8_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_8_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_8_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_8_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_9_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_9_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_9_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_9_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_9_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_9_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_9_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_10_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_10_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_10_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_10_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_10_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_10_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_10_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_11_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_11_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_11_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_11_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_11_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_11_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_11_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_12_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_12_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_12_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_12_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_12_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_12_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_12_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_13_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_13_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_13_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_13_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_13_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_13_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_13_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_14_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_14_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_14_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_14_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_14_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_14_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_14_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_15_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_15_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_15_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_15_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_15_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_15_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_15_branch_mask; // @[fifo.scala 27:33]
  reg [3:0] readPtr; // @[fifo.scala 33:25]
  wire [3:0] _nextVal_T_2 = readPtr + 4'h1; // @[fifo.scala 34:60]
  wire [3:0] nextRead = readPtr == 4'hf ? 4'h0 : _nextVal_T_2; // @[fifo.scala 34:22]
  wire [1:0] op = {write_data_valid,read_ready}; // @[fifo.scala 46:29]
  reg  emptyReg; // @[fifo.scala 43:25]
  wire  _T_2 = ~emptyReg; // @[fifo.scala 52:12]
  wire  _GEN_21 = 2'h2 == op ? 1'h0 : 2'h3 == op & _T_2; // @[fifo.scala 49:14]
  wire  _GEN_24 = 2'h1 == op ? _T_2 : _GEN_21; // @[fifo.scala 49:14]
  wire  incrRead = 2'h0 == op ? 1'h0 : _GEN_24; // @[fifo.scala 49:14]
  reg [3:0] writePtr; // @[fifo.scala 33:25]
  wire [3:0] _nextVal_T_5 = writePtr + 4'h1; // @[fifo.scala 34:60]
  wire [3:0] nextWrite = writePtr == 4'hf ? 4'h0 : _nextVal_T_5; // @[fifo.scala 34:22]
  reg  fullReg; // @[fifo.scala 44:34]
  wire  _T_4 = ~fullReg; // @[fifo.scala 59:12]
  wire  _GEN_18 = 2'h2 == op ? _T_4 : 2'h3 == op & _T_4; // @[fifo.scala 49:14]
  wire  _GEN_25 = 2'h1 == op ? 1'h0 : _GEN_18; // @[fifo.scala 49:14]
  wire  incrWrite = 2'h0 == op ? 1'h0 : _GEN_25; // @[fifo.scala 49:14]
  wire  _GEN_3 = ~emptyReg ? nextRead == writePtr : emptyReg; // @[fifo.scala 52:23 54:18 43:25]
  wire  _GEN_6 = ~fullReg ? 1'h0 : emptyReg; // @[fifo.scala 59:22 61:18 43:25]
  wire  _GEN_7 = ~fullReg ? nextWrite == readPtr : fullReg; // @[fifo.scala 59:22 62:17 44:34]
  wire  _fullReg_T_2 = emptyReg ? 1'h0 : nextWrite == nextRead; // @[fifo.scala 70:23]
  wire  _GEN_10 = _T_4 ? _fullReg_T_2 : fullReg; // @[fifo.scala 67:22 70:17 44:34]
  wire  _emptyReg_T_2 = fullReg ? 1'h0 : nextRead == nextWrite; // @[fifo.scala 75:24]
  wire  _GEN_11 = _T_2 ? 1'h0 : _GEN_10; // @[fifo.scala 73:23 74:17]
  wire  _GEN_12 = _T_2 ? _emptyReg_T_2 : _GEN_6; // @[fifo.scala 73:23 75:18]
  wire  _GEN_15 = 2'h3 == op ? _GEN_12 : emptyReg; // @[fifo.scala 49:14 43:25]
  wire  _GEN_16 = 2'h3 == op ? _GEN_11 : fullReg; // @[fifo.scala 49:14 44:34]
  wire  _GEN_19 = 2'h2 == op ? _GEN_6 : _GEN_15; // @[fifo.scala 49:14]
  wire  _GEN_23 = 2'h1 == op ? _GEN_3 : _GEN_19; // @[fifo.scala 49:14]
  wire  _GEN_27 = 2'h0 == op ? emptyReg : _GEN_23; // @[fifo.scala 49:14 43:25]
  wire  _GEN_110 = 4'h0 == writePtr ? write_data_branch_valid : memReg_0_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_111 = 4'h1 == writePtr ? write_data_branch_valid : memReg_1_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_112 = 4'h2 == writePtr ? write_data_branch_valid : memReg_2_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_113 = 4'h3 == writePtr ? write_data_branch_valid : memReg_3_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_114 = 4'h4 == writePtr ? write_data_branch_valid : memReg_4_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_115 = 4'h5 == writePtr ? write_data_branch_valid : memReg_5_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_116 = 4'h6 == writePtr ? write_data_branch_valid : memReg_6_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_117 = 4'h7 == writePtr ? write_data_branch_valid : memReg_7_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_118 = 4'h8 == writePtr ? write_data_branch_valid : memReg_8_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_119 = 4'h9 == writePtr ? write_data_branch_valid : memReg_9_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_120 = 4'ha == writePtr ? write_data_branch_valid : memReg_10_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_121 = 4'hb == writePtr ? write_data_branch_valid : memReg_11_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_122 = 4'hc == writePtr ? write_data_branch_valid : memReg_12_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_123 = 4'hd == writePtr ? write_data_branch_valid : memReg_13_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_124 = 4'he == writePtr ? write_data_branch_valid : memReg_14_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_125 = 4'hf == writePtr ? write_data_branch_valid : memReg_15_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_126 = 4'h0 == writePtr ? write_data_branch_mask : memReg_0_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_127 = 4'h1 == writePtr ? write_data_branch_mask : memReg_1_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_128 = 4'h2 == writePtr ? write_data_branch_mask : memReg_2_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_129 = 4'h3 == writePtr ? write_data_branch_mask : memReg_3_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_130 = 4'h4 == writePtr ? write_data_branch_mask : memReg_4_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_131 = 4'h5 == writePtr ? write_data_branch_mask : memReg_5_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_132 = 4'h6 == writePtr ? write_data_branch_mask : memReg_6_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_133 = 4'h7 == writePtr ? write_data_branch_mask : memReg_7_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_134 = 4'h8 == writePtr ? write_data_branch_mask : memReg_8_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_135 = 4'h9 == writePtr ? write_data_branch_mask : memReg_9_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_136 = 4'ha == writePtr ? write_data_branch_mask : memReg_10_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_137 = 4'hb == writePtr ? write_data_branch_mask : memReg_11_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_138 = 4'hc == writePtr ? write_data_branch_mask : memReg_12_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_139 = 4'hd == writePtr ? write_data_branch_mask : memReg_13_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_140 = 4'he == writePtr ? write_data_branch_mask : memReg_14_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_141 = 4'hf == writePtr ? write_data_branch_mask : memReg_15_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_302 = incrWrite ? _GEN_110 : memReg_0_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_303 = incrWrite ? _GEN_111 : memReg_1_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_304 = incrWrite ? _GEN_112 : memReg_2_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_305 = incrWrite ? _GEN_113 : memReg_3_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_306 = incrWrite ? _GEN_114 : memReg_4_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_307 = incrWrite ? _GEN_115 : memReg_5_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_308 = incrWrite ? _GEN_116 : memReg_6_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_309 = incrWrite ? _GEN_117 : memReg_7_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_310 = incrWrite ? _GEN_118 : memReg_8_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_311 = incrWrite ? _GEN_119 : memReg_9_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_312 = incrWrite ? _GEN_120 : memReg_10_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_313 = incrWrite ? _GEN_121 : memReg_11_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_314 = incrWrite ? _GEN_122 : memReg_12_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_315 = incrWrite ? _GEN_123 : memReg_13_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_316 = incrWrite ? _GEN_124 : memReg_14_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_317 = incrWrite ? _GEN_125 : memReg_15_branch_valid; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_318 = incrWrite ? _GEN_126 : memReg_0_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_319 = incrWrite ? _GEN_127 : memReg_1_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_320 = incrWrite ? _GEN_128 : memReg_2_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_321 = incrWrite ? _GEN_129 : memReg_3_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_322 = incrWrite ? _GEN_130 : memReg_4_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_323 = incrWrite ? _GEN_131 : memReg_5_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_324 = incrWrite ? _GEN_132 : memReg_6_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_325 = incrWrite ? _GEN_133 : memReg_7_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_326 = incrWrite ? _GEN_134 : memReg_8_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_327 = incrWrite ? _GEN_135 : memReg_9_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_328 = incrWrite ? _GEN_136 : memReg_10_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_329 = incrWrite ? _GEN_137 : memReg_11_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_330 = incrWrite ? _GEN_138 : memReg_12_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_331 = incrWrite ? _GEN_139 : memReg_13_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_332 = incrWrite ? _GEN_140 : memReg_14_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_333 = incrWrite ? _GEN_141 : memReg_15_branch_mask; // @[fifo.scala 81:17 27:33]
  wire  _GEN_415 = 4'h1 == readPtr ? memReg_1_valid : memReg_0_valid; // @[fifo.scala 86:{13,13}]
  wire  _GEN_416 = 4'h2 == readPtr ? memReg_2_valid : _GEN_415; // @[fifo.scala 86:{13,13}]
  wire  _GEN_417 = 4'h3 == readPtr ? memReg_3_valid : _GEN_416; // @[fifo.scala 86:{13,13}]
  wire  _GEN_418 = 4'h4 == readPtr ? memReg_4_valid : _GEN_417; // @[fifo.scala 86:{13,13}]
  wire  _GEN_419 = 4'h5 == readPtr ? memReg_5_valid : _GEN_418; // @[fifo.scala 86:{13,13}]
  wire  _GEN_420 = 4'h6 == readPtr ? memReg_6_valid : _GEN_419; // @[fifo.scala 86:{13,13}]
  wire  _GEN_421 = 4'h7 == readPtr ? memReg_7_valid : _GEN_420; // @[fifo.scala 86:{13,13}]
  wire  _GEN_422 = 4'h8 == readPtr ? memReg_8_valid : _GEN_421; // @[fifo.scala 86:{13,13}]
  wire  _GEN_423 = 4'h9 == readPtr ? memReg_9_valid : _GEN_422; // @[fifo.scala 86:{13,13}]
  wire  _GEN_424 = 4'ha == readPtr ? memReg_10_valid : _GEN_423; // @[fifo.scala 86:{13,13}]
  wire  _GEN_425 = 4'hb == readPtr ? memReg_11_valid : _GEN_424; // @[fifo.scala 86:{13,13}]
  wire  _GEN_426 = 4'hc == readPtr ? memReg_12_valid : _GEN_425; // @[fifo.scala 86:{13,13}]
  wire  _GEN_427 = 4'hd == readPtr ? memReg_13_valid : _GEN_426; // @[fifo.scala 86:{13,13}]
  wire  _GEN_428 = 4'he == readPtr ? memReg_14_valid : _GEN_427; // @[fifo.scala 86:{13,13}]
  wire  _GEN_429 = 4'hf == readPtr ? memReg_15_valid : _GEN_428; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_431 = 4'h1 == readPtr ? memReg_1_address : memReg_0_address; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_432 = 4'h2 == readPtr ? memReg_2_address : _GEN_431; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_433 = 4'h3 == readPtr ? memReg_3_address : _GEN_432; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_434 = 4'h4 == readPtr ? memReg_4_address : _GEN_433; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_435 = 4'h5 == readPtr ? memReg_5_address : _GEN_434; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_436 = 4'h6 == readPtr ? memReg_6_address : _GEN_435; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_437 = 4'h7 == readPtr ? memReg_7_address : _GEN_436; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_438 = 4'h8 == readPtr ? memReg_8_address : _GEN_437; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_439 = 4'h9 == readPtr ? memReg_9_address : _GEN_438; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_440 = 4'ha == readPtr ? memReg_10_address : _GEN_439; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_441 = 4'hb == readPtr ? memReg_11_address : _GEN_440; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_442 = 4'hc == readPtr ? memReg_12_address : _GEN_441; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_443 = 4'hd == readPtr ? memReg_13_address : _GEN_442; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_444 = 4'he == readPtr ? memReg_14_address : _GEN_443; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_447 = 4'h1 == readPtr ? memReg_1_core_instruction : memReg_0_core_instruction; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_448 = 4'h2 == readPtr ? memReg_2_core_instruction : _GEN_447; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_449 = 4'h3 == readPtr ? memReg_3_core_instruction : _GEN_448; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_450 = 4'h4 == readPtr ? memReg_4_core_instruction : _GEN_449; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_451 = 4'h5 == readPtr ? memReg_5_core_instruction : _GEN_450; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_452 = 4'h6 == readPtr ? memReg_6_core_instruction : _GEN_451; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_453 = 4'h7 == readPtr ? memReg_7_core_instruction : _GEN_452; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_454 = 4'h8 == readPtr ? memReg_8_core_instruction : _GEN_453; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_455 = 4'h9 == readPtr ? memReg_9_core_instruction : _GEN_454; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_456 = 4'ha == readPtr ? memReg_10_core_instruction : _GEN_455; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_457 = 4'hb == readPtr ? memReg_11_core_instruction : _GEN_456; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_458 = 4'hc == readPtr ? memReg_12_core_instruction : _GEN_457; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_459 = 4'hd == readPtr ? memReg_13_core_instruction : _GEN_458; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_460 = 4'he == readPtr ? memReg_14_core_instruction : _GEN_459; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_463 = 4'h1 == readPtr ? memReg_1_core_robAddr : memReg_0_core_robAddr; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_464 = 4'h2 == readPtr ? memReg_2_core_robAddr : _GEN_463; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_465 = 4'h3 == readPtr ? memReg_3_core_robAddr : _GEN_464; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_466 = 4'h4 == readPtr ? memReg_4_core_robAddr : _GEN_465; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_467 = 4'h5 == readPtr ? memReg_5_core_robAddr : _GEN_466; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_468 = 4'h6 == readPtr ? memReg_6_core_robAddr : _GEN_467; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_469 = 4'h7 == readPtr ? memReg_7_core_robAddr : _GEN_468; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_470 = 4'h8 == readPtr ? memReg_8_core_robAddr : _GEN_469; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_471 = 4'h9 == readPtr ? memReg_9_core_robAddr : _GEN_470; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_472 = 4'ha == readPtr ? memReg_10_core_robAddr : _GEN_471; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_473 = 4'hb == readPtr ? memReg_11_core_robAddr : _GEN_472; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_474 = 4'hc == readPtr ? memReg_12_core_robAddr : _GEN_473; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_475 = 4'hd == readPtr ? memReg_13_core_robAddr : _GEN_474; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_476 = 4'he == readPtr ? memReg_14_core_robAddr : _GEN_475; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_479 = 4'h1 == readPtr ? memReg_1_core_prfDest : memReg_0_core_prfDest; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_480 = 4'h2 == readPtr ? memReg_2_core_prfDest : _GEN_479; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_481 = 4'h3 == readPtr ? memReg_3_core_prfDest : _GEN_480; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_482 = 4'h4 == readPtr ? memReg_4_core_prfDest : _GEN_481; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_483 = 4'h5 == readPtr ? memReg_5_core_prfDest : _GEN_482; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_484 = 4'h6 == readPtr ? memReg_6_core_prfDest : _GEN_483; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_485 = 4'h7 == readPtr ? memReg_7_core_prfDest : _GEN_484; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_486 = 4'h8 == readPtr ? memReg_8_core_prfDest : _GEN_485; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_487 = 4'h9 == readPtr ? memReg_9_core_prfDest : _GEN_486; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_488 = 4'ha == readPtr ? memReg_10_core_prfDest : _GEN_487; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_489 = 4'hb == readPtr ? memReg_11_core_prfDest : _GEN_488; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_490 = 4'hc == readPtr ? memReg_12_core_prfDest : _GEN_489; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_491 = 4'hd == readPtr ? memReg_13_core_prfDest : _GEN_490; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_492 = 4'he == readPtr ? memReg_14_core_prfDest : _GEN_491; // @[fifo.scala 86:{13,13}]
  wire  _GEN_495 = 4'h1 == readPtr ? memReg_1_branch_valid : memReg_0_branch_valid; // @[fifo.scala 86:{13,13}]
  wire  _GEN_496 = 4'h2 == readPtr ? memReg_2_branch_valid : _GEN_495; // @[fifo.scala 86:{13,13}]
  wire  _GEN_497 = 4'h3 == readPtr ? memReg_3_branch_valid : _GEN_496; // @[fifo.scala 86:{13,13}]
  wire  _GEN_498 = 4'h4 == readPtr ? memReg_4_branch_valid : _GEN_497; // @[fifo.scala 86:{13,13}]
  wire  _GEN_499 = 4'h5 == readPtr ? memReg_5_branch_valid : _GEN_498; // @[fifo.scala 86:{13,13}]
  wire  _GEN_500 = 4'h6 == readPtr ? memReg_6_branch_valid : _GEN_499; // @[fifo.scala 86:{13,13}]
  wire  _GEN_501 = 4'h7 == readPtr ? memReg_7_branch_valid : _GEN_500; // @[fifo.scala 86:{13,13}]
  wire  _GEN_502 = 4'h8 == readPtr ? memReg_8_branch_valid : _GEN_501; // @[fifo.scala 86:{13,13}]
  wire  _GEN_503 = 4'h9 == readPtr ? memReg_9_branch_valid : _GEN_502; // @[fifo.scala 86:{13,13}]
  wire  _GEN_504 = 4'ha == readPtr ? memReg_10_branch_valid : _GEN_503; // @[fifo.scala 86:{13,13}]
  wire  _GEN_505 = 4'hb == readPtr ? memReg_11_branch_valid : _GEN_504; // @[fifo.scala 86:{13,13}]
  wire  _GEN_506 = 4'hc == readPtr ? memReg_12_branch_valid : _GEN_505; // @[fifo.scala 86:{13,13}]
  wire  _GEN_507 = 4'hd == readPtr ? memReg_13_branch_valid : _GEN_506; // @[fifo.scala 86:{13,13}]
  wire  _GEN_508 = 4'he == readPtr ? memReg_14_branch_valid : _GEN_507; // @[fifo.scala 86:{13,13}]
  wire  _GEN_509 = 4'hf == readPtr ? memReg_15_branch_valid : _GEN_508; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_511 = 4'h1 == readPtr ? memReg_1_branch_mask : memReg_0_branch_mask; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_512 = 4'h2 == readPtr ? memReg_2_branch_mask : _GEN_511; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_513 = 4'h3 == readPtr ? memReg_3_branch_mask : _GEN_512; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_514 = 4'h4 == readPtr ? memReg_4_branch_mask : _GEN_513; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_515 = 4'h5 == readPtr ? memReg_5_branch_mask : _GEN_514; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_516 = 4'h6 == readPtr ? memReg_6_branch_mask : _GEN_515; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_517 = 4'h7 == readPtr ? memReg_7_branch_mask : _GEN_516; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_518 = 4'h8 == readPtr ? memReg_8_branch_mask : _GEN_517; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_519 = 4'h9 == readPtr ? memReg_9_branch_mask : _GEN_518; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_520 = 4'ha == readPtr ? memReg_10_branch_mask : _GEN_519; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_521 = 4'hb == readPtr ? memReg_11_branch_mask : _GEN_520; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_522 = 4'hc == readPtr ? memReg_12_branch_mask : _GEN_521; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_523 = 4'hd == readPtr ? memReg_13_branch_mask : _GEN_522; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_524 = 4'he == readPtr ? memReg_14_branch_mask : _GEN_523; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_525 = 4'hf == readPtr ? memReg_15_branch_mask : _GEN_524; // @[fifo.scala 86:{13,13}]
  wire [4:0] _T_8 = write_data_branch_mask & branchOps_branchMask; // @[utils.scala 62:31]
  wire  _T_9 = |_T_8; // @[utils.scala 62:55]
  wire [4:0] _memReg_branch_mask_T = write_data_branch_mask ^ branchOps_branchMask; // @[utils.scala 63:42]
  wire [4:0] _GEN_606 = 4'h0 == writePtr ? _memReg_branch_mask_T : _GEN_318; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_607 = 4'h1 == writePtr ? _memReg_branch_mask_T : _GEN_319; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_608 = 4'h2 == writePtr ? _memReg_branch_mask_T : _GEN_320; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_609 = 4'h3 == writePtr ? _memReg_branch_mask_T : _GEN_321; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_610 = 4'h4 == writePtr ? _memReg_branch_mask_T : _GEN_322; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_611 = 4'h5 == writePtr ? _memReg_branch_mask_T : _GEN_323; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_612 = 4'h6 == writePtr ? _memReg_branch_mask_T : _GEN_324; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_613 = 4'h7 == writePtr ? _memReg_branch_mask_T : _GEN_325; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_614 = 4'h8 == writePtr ? _memReg_branch_mask_T : _GEN_326; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_615 = 4'h9 == writePtr ? _memReg_branch_mask_T : _GEN_327; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_616 = 4'ha == writePtr ? _memReg_branch_mask_T : _GEN_328; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_617 = 4'hb == writePtr ? _memReg_branch_mask_T : _GEN_329; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_618 = 4'hc == writePtr ? _memReg_branch_mask_T : _GEN_330; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_619 = 4'hd == writePtr ? _memReg_branch_mask_T : _GEN_331; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_620 = 4'he == writePtr ? _memReg_branch_mask_T : _GEN_332; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_621 = 4'hf == writePtr ? _memReg_branch_mask_T : _GEN_333; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_622 = 4'h0 == writePtr ? write_data_branch_mask : _GEN_318; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_623 = 4'h1 == writePtr ? write_data_branch_mask : _GEN_319; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_624 = 4'h2 == writePtr ? write_data_branch_mask : _GEN_320; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_625 = 4'h3 == writePtr ? write_data_branch_mask : _GEN_321; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_626 = 4'h4 == writePtr ? write_data_branch_mask : _GEN_322; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_627 = 4'h5 == writePtr ? write_data_branch_mask : _GEN_323; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_628 = 4'h6 == writePtr ? write_data_branch_mask : _GEN_324; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_629 = 4'h7 == writePtr ? write_data_branch_mask : _GEN_325; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_630 = 4'h8 == writePtr ? write_data_branch_mask : _GEN_326; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_631 = 4'h9 == writePtr ? write_data_branch_mask : _GEN_327; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_632 = 4'ha == writePtr ? write_data_branch_mask : _GEN_328; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_633 = 4'hb == writePtr ? write_data_branch_mask : _GEN_329; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_634 = 4'hc == writePtr ? write_data_branch_mask : _GEN_330; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_635 = 4'hd == writePtr ? write_data_branch_mask : _GEN_331; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_636 = 4'he == writePtr ? write_data_branch_mask : _GEN_332; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_637 = 4'hf == writePtr ? write_data_branch_mask : _GEN_333; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_638 = |_T_8 ? _GEN_606 : _GEN_622; // @[utils.scala 62:60]
  wire [4:0] _GEN_639 = |_T_8 ? _GEN_607 : _GEN_623; // @[utils.scala 62:60]
  wire [4:0] _GEN_640 = |_T_8 ? _GEN_608 : _GEN_624; // @[utils.scala 62:60]
  wire [4:0] _GEN_641 = |_T_8 ? _GEN_609 : _GEN_625; // @[utils.scala 62:60]
  wire [4:0] _GEN_642 = |_T_8 ? _GEN_610 : _GEN_626; // @[utils.scala 62:60]
  wire [4:0] _GEN_643 = |_T_8 ? _GEN_611 : _GEN_627; // @[utils.scala 62:60]
  wire [4:0] _GEN_644 = |_T_8 ? _GEN_612 : _GEN_628; // @[utils.scala 62:60]
  wire [4:0] _GEN_645 = |_T_8 ? _GEN_613 : _GEN_629; // @[utils.scala 62:60]
  wire [4:0] _GEN_646 = |_T_8 ? _GEN_614 : _GEN_630; // @[utils.scala 62:60]
  wire [4:0] _GEN_647 = |_T_8 ? _GEN_615 : _GEN_631; // @[utils.scala 62:60]
  wire [4:0] _GEN_648 = |_T_8 ? _GEN_616 : _GEN_632; // @[utils.scala 62:60]
  wire [4:0] _GEN_649 = |_T_8 ? _GEN_617 : _GEN_633; // @[utils.scala 62:60]
  wire [4:0] _GEN_650 = |_T_8 ? _GEN_618 : _GEN_634; // @[utils.scala 62:60]
  wire [4:0] _GEN_651 = |_T_8 ? _GEN_619 : _GEN_635; // @[utils.scala 62:60]
  wire [4:0] _GEN_652 = |_T_8 ? _GEN_620 : _GEN_636; // @[utils.scala 62:60]
  wire [4:0] _GEN_653 = |_T_8 ? _GEN_621 : _GEN_637; // @[utils.scala 62:60]
  wire  _GEN_654 = 4'h0 == writePtr ? write_data_branch_valid : _GEN_302; // @[utils.scala 67:{22,22}]
  wire  _GEN_655 = 4'h1 == writePtr ? write_data_branch_valid : _GEN_303; // @[utils.scala 67:{22,22}]
  wire  _GEN_656 = 4'h2 == writePtr ? write_data_branch_valid : _GEN_304; // @[utils.scala 67:{22,22}]
  wire  _GEN_657 = 4'h3 == writePtr ? write_data_branch_valid : _GEN_305; // @[utils.scala 67:{22,22}]
  wire  _GEN_658 = 4'h4 == writePtr ? write_data_branch_valid : _GEN_306; // @[utils.scala 67:{22,22}]
  wire  _GEN_659 = 4'h5 == writePtr ? write_data_branch_valid : _GEN_307; // @[utils.scala 67:{22,22}]
  wire  _GEN_660 = 4'h6 == writePtr ? write_data_branch_valid : _GEN_308; // @[utils.scala 67:{22,22}]
  wire  _GEN_661 = 4'h7 == writePtr ? write_data_branch_valid : _GEN_309; // @[utils.scala 67:{22,22}]
  wire  _GEN_662 = 4'h8 == writePtr ? write_data_branch_valid : _GEN_310; // @[utils.scala 67:{22,22}]
  wire  _GEN_663 = 4'h9 == writePtr ? write_data_branch_valid : _GEN_311; // @[utils.scala 67:{22,22}]
  wire  _GEN_664 = 4'ha == writePtr ? write_data_branch_valid : _GEN_312; // @[utils.scala 67:{22,22}]
  wire  _GEN_665 = 4'hb == writePtr ? write_data_branch_valid : _GEN_313; // @[utils.scala 67:{22,22}]
  wire  _GEN_666 = 4'hc == writePtr ? write_data_branch_valid : _GEN_314; // @[utils.scala 67:{22,22}]
  wire  _GEN_667 = 4'hd == writePtr ? write_data_branch_valid : _GEN_315; // @[utils.scala 67:{22,22}]
  wire  _GEN_668 = 4'he == writePtr ? write_data_branch_valid : _GEN_316; // @[utils.scala 67:{22,22}]
  wire  _GEN_669 = 4'hf == writePtr ? write_data_branch_valid : _GEN_317; // @[utils.scala 67:{22,22}]
  wire  _GEN_670 = 4'h0 == writePtr ? 1'h0 : _GEN_302; // @[utils.scala 71:{24,24}]
  wire  _GEN_671 = 4'h1 == writePtr ? 1'h0 : _GEN_303; // @[utils.scala 71:{24,24}]
  wire  _GEN_672 = 4'h2 == writePtr ? 1'h0 : _GEN_304; // @[utils.scala 71:{24,24}]
  wire  _GEN_673 = 4'h3 == writePtr ? 1'h0 : _GEN_305; // @[utils.scala 71:{24,24}]
  wire  _GEN_674 = 4'h4 == writePtr ? 1'h0 : _GEN_306; // @[utils.scala 71:{24,24}]
  wire  _GEN_675 = 4'h5 == writePtr ? 1'h0 : _GEN_307; // @[utils.scala 71:{24,24}]
  wire  _GEN_676 = 4'h6 == writePtr ? 1'h0 : _GEN_308; // @[utils.scala 71:{24,24}]
  wire  _GEN_677 = 4'h7 == writePtr ? 1'h0 : _GEN_309; // @[utils.scala 71:{24,24}]
  wire  _GEN_678 = 4'h8 == writePtr ? 1'h0 : _GEN_310; // @[utils.scala 71:{24,24}]
  wire  _GEN_679 = 4'h9 == writePtr ? 1'h0 : _GEN_311; // @[utils.scala 71:{24,24}]
  wire  _GEN_680 = 4'ha == writePtr ? 1'h0 : _GEN_312; // @[utils.scala 71:{24,24}]
  wire  _GEN_681 = 4'hb == writePtr ? 1'h0 : _GEN_313; // @[utils.scala 71:{24,24}]
  wire  _GEN_682 = 4'hc == writePtr ? 1'h0 : _GEN_314; // @[utils.scala 71:{24,24}]
  wire  _GEN_683 = 4'hd == writePtr ? 1'h0 : _GEN_315; // @[utils.scala 71:{24,24}]
  wire  _GEN_684 = 4'he == writePtr ? 1'h0 : _GEN_316; // @[utils.scala 71:{24,24}]
  wire  _GEN_685 = 4'hf == writePtr ? 1'h0 : _GEN_317; // @[utils.scala 71:{24,24}]
  wire [4:0] _GEN_686 = 4'h0 == writePtr ? 5'h0 : _GEN_318; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_687 = 4'h1 == writePtr ? 5'h0 : _GEN_319; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_688 = 4'h2 == writePtr ? 5'h0 : _GEN_320; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_689 = 4'h3 == writePtr ? 5'h0 : _GEN_321; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_690 = 4'h4 == writePtr ? 5'h0 : _GEN_322; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_691 = 4'h5 == writePtr ? 5'h0 : _GEN_323; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_692 = 4'h6 == writePtr ? 5'h0 : _GEN_324; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_693 = 4'h7 == writePtr ? 5'h0 : _GEN_325; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_694 = 4'h8 == writePtr ? 5'h0 : _GEN_326; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_695 = 4'h9 == writePtr ? 5'h0 : _GEN_327; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_696 = 4'ha == writePtr ? 5'h0 : _GEN_328; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_697 = 4'hb == writePtr ? 5'h0 : _GEN_329; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_698 = 4'hc == writePtr ? 5'h0 : _GEN_330; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_699 = 4'hd == writePtr ? 5'h0 : _GEN_331; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_700 = 4'he == writePtr ? 5'h0 : _GEN_332; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_701 = 4'hf == writePtr ? 5'h0 : _GEN_333; // @[utils.scala 72:{23,23}]
  wire  _GEN_734 = _T_9 ? _GEN_670 : _GEN_654; // @[utils.scala 70:60]
  wire  _GEN_735 = _T_9 ? _GEN_671 : _GEN_655; // @[utils.scala 70:60]
  wire  _GEN_736 = _T_9 ? _GEN_672 : _GEN_656; // @[utils.scala 70:60]
  wire  _GEN_737 = _T_9 ? _GEN_673 : _GEN_657; // @[utils.scala 70:60]
  wire  _GEN_738 = _T_9 ? _GEN_674 : _GEN_658; // @[utils.scala 70:60]
  wire  _GEN_739 = _T_9 ? _GEN_675 : _GEN_659; // @[utils.scala 70:60]
  wire  _GEN_740 = _T_9 ? _GEN_676 : _GEN_660; // @[utils.scala 70:60]
  wire  _GEN_741 = _T_9 ? _GEN_677 : _GEN_661; // @[utils.scala 70:60]
  wire  _GEN_742 = _T_9 ? _GEN_678 : _GEN_662; // @[utils.scala 70:60]
  wire  _GEN_743 = _T_9 ? _GEN_679 : _GEN_663; // @[utils.scala 70:60]
  wire  _GEN_744 = _T_9 ? _GEN_680 : _GEN_664; // @[utils.scala 70:60]
  wire  _GEN_745 = _T_9 ? _GEN_681 : _GEN_665; // @[utils.scala 70:60]
  wire  _GEN_746 = _T_9 ? _GEN_682 : _GEN_666; // @[utils.scala 70:60]
  wire  _GEN_747 = _T_9 ? _GEN_683 : _GEN_667; // @[utils.scala 70:60]
  wire  _GEN_748 = _T_9 ? _GEN_684 : _GEN_668; // @[utils.scala 70:60]
  wire  _GEN_749 = _T_9 ? _GEN_685 : _GEN_669; // @[utils.scala 70:60]
  wire [4:0] _GEN_750 = _T_9 ? _GEN_686 : _GEN_622; // @[utils.scala 70:60]
  wire [4:0] _GEN_751 = _T_9 ? _GEN_687 : _GEN_623; // @[utils.scala 70:60]
  wire [4:0] _GEN_752 = _T_9 ? _GEN_688 : _GEN_624; // @[utils.scala 70:60]
  wire [4:0] _GEN_753 = _T_9 ? _GEN_689 : _GEN_625; // @[utils.scala 70:60]
  wire [4:0] _GEN_754 = _T_9 ? _GEN_690 : _GEN_626; // @[utils.scala 70:60]
  wire [4:0] _GEN_755 = _T_9 ? _GEN_691 : _GEN_627; // @[utils.scala 70:60]
  wire [4:0] _GEN_756 = _T_9 ? _GEN_692 : _GEN_628; // @[utils.scala 70:60]
  wire [4:0] _GEN_757 = _T_9 ? _GEN_693 : _GEN_629; // @[utils.scala 70:60]
  wire [4:0] _GEN_758 = _T_9 ? _GEN_694 : _GEN_630; // @[utils.scala 70:60]
  wire [4:0] _GEN_759 = _T_9 ? _GEN_695 : _GEN_631; // @[utils.scala 70:60]
  wire [4:0] _GEN_760 = _T_9 ? _GEN_696 : _GEN_632; // @[utils.scala 70:60]
  wire [4:0] _GEN_761 = _T_9 ? _GEN_697 : _GEN_633; // @[utils.scala 70:60]
  wire [4:0] _GEN_762 = _T_9 ? _GEN_698 : _GEN_634; // @[utils.scala 70:60]
  wire [4:0] _GEN_763 = _T_9 ? _GEN_699 : _GEN_635; // @[utils.scala 70:60]
  wire [4:0] _GEN_764 = _T_9 ? _GEN_700 : _GEN_636; // @[utils.scala 70:60]
  wire [4:0] _GEN_765 = _T_9 ? _GEN_701 : _GEN_637; // @[utils.scala 70:60]
  wire [4:0] _GEN_766 = branchOps_passed ? _GEN_638 : _GEN_750; // @[utils.scala 60:30]
  wire [4:0] _GEN_767 = branchOps_passed ? _GEN_639 : _GEN_751; // @[utils.scala 60:30]
  wire [4:0] _GEN_768 = branchOps_passed ? _GEN_640 : _GEN_752; // @[utils.scala 60:30]
  wire [4:0] _GEN_769 = branchOps_passed ? _GEN_641 : _GEN_753; // @[utils.scala 60:30]
  wire [4:0] _GEN_770 = branchOps_passed ? _GEN_642 : _GEN_754; // @[utils.scala 60:30]
  wire [4:0] _GEN_771 = branchOps_passed ? _GEN_643 : _GEN_755; // @[utils.scala 60:30]
  wire [4:0] _GEN_772 = branchOps_passed ? _GEN_644 : _GEN_756; // @[utils.scala 60:30]
  wire [4:0] _GEN_773 = branchOps_passed ? _GEN_645 : _GEN_757; // @[utils.scala 60:30]
  wire [4:0] _GEN_774 = branchOps_passed ? _GEN_646 : _GEN_758; // @[utils.scala 60:30]
  wire [4:0] _GEN_775 = branchOps_passed ? _GEN_647 : _GEN_759; // @[utils.scala 60:30]
  wire [4:0] _GEN_776 = branchOps_passed ? _GEN_648 : _GEN_760; // @[utils.scala 60:30]
  wire [4:0] _GEN_777 = branchOps_passed ? _GEN_649 : _GEN_761; // @[utils.scala 60:30]
  wire [4:0] _GEN_778 = branchOps_passed ? _GEN_650 : _GEN_762; // @[utils.scala 60:30]
  wire [4:0] _GEN_779 = branchOps_passed ? _GEN_651 : _GEN_763; // @[utils.scala 60:30]
  wire [4:0] _GEN_780 = branchOps_passed ? _GEN_652 : _GEN_764; // @[utils.scala 60:30]
  wire [4:0] _GEN_781 = branchOps_passed ? _GEN_653 : _GEN_765; // @[utils.scala 60:30]
  wire  _GEN_782 = branchOps_passed ? _GEN_654 : _GEN_734; // @[utils.scala 60:30]
  wire  _GEN_783 = branchOps_passed ? _GEN_655 : _GEN_735; // @[utils.scala 60:30]
  wire  _GEN_784 = branchOps_passed ? _GEN_656 : _GEN_736; // @[utils.scala 60:30]
  wire  _GEN_785 = branchOps_passed ? _GEN_657 : _GEN_737; // @[utils.scala 60:30]
  wire  _GEN_786 = branchOps_passed ? _GEN_658 : _GEN_738; // @[utils.scala 60:30]
  wire  _GEN_787 = branchOps_passed ? _GEN_659 : _GEN_739; // @[utils.scala 60:30]
  wire  _GEN_788 = branchOps_passed ? _GEN_660 : _GEN_740; // @[utils.scala 60:30]
  wire  _GEN_789 = branchOps_passed ? _GEN_661 : _GEN_741; // @[utils.scala 60:30]
  wire  _GEN_790 = branchOps_passed ? _GEN_662 : _GEN_742; // @[utils.scala 60:30]
  wire  _GEN_791 = branchOps_passed ? _GEN_663 : _GEN_743; // @[utils.scala 60:30]
  wire  _GEN_792 = branchOps_passed ? _GEN_664 : _GEN_744; // @[utils.scala 60:30]
  wire  _GEN_793 = branchOps_passed ? _GEN_665 : _GEN_745; // @[utils.scala 60:30]
  wire  _GEN_794 = branchOps_passed ? _GEN_666 : _GEN_746; // @[utils.scala 60:30]
  wire  _GEN_795 = branchOps_passed ? _GEN_667 : _GEN_747; // @[utils.scala 60:30]
  wire  _GEN_796 = branchOps_passed ? _GEN_668 : _GEN_748; // @[utils.scala 60:30]
  wire  _GEN_797 = branchOps_passed ? _GEN_669 : _GEN_749; // @[utils.scala 60:30]
  wire [4:0] _GEN_830 = branchOps_valid ? _GEN_766 : _GEN_622; // @[utils.scala 59:26]
  wire [4:0] _GEN_831 = branchOps_valid ? _GEN_767 : _GEN_623; // @[utils.scala 59:26]
  wire [4:0] _GEN_832 = branchOps_valid ? _GEN_768 : _GEN_624; // @[utils.scala 59:26]
  wire [4:0] _GEN_833 = branchOps_valid ? _GEN_769 : _GEN_625; // @[utils.scala 59:26]
  wire [4:0] _GEN_834 = branchOps_valid ? _GEN_770 : _GEN_626; // @[utils.scala 59:26]
  wire [4:0] _GEN_835 = branchOps_valid ? _GEN_771 : _GEN_627; // @[utils.scala 59:26]
  wire [4:0] _GEN_836 = branchOps_valid ? _GEN_772 : _GEN_628; // @[utils.scala 59:26]
  wire [4:0] _GEN_837 = branchOps_valid ? _GEN_773 : _GEN_629; // @[utils.scala 59:26]
  wire [4:0] _GEN_838 = branchOps_valid ? _GEN_774 : _GEN_630; // @[utils.scala 59:26]
  wire [4:0] _GEN_839 = branchOps_valid ? _GEN_775 : _GEN_631; // @[utils.scala 59:26]
  wire [4:0] _GEN_840 = branchOps_valid ? _GEN_776 : _GEN_632; // @[utils.scala 59:26]
  wire [4:0] _GEN_841 = branchOps_valid ? _GEN_777 : _GEN_633; // @[utils.scala 59:26]
  wire [4:0] _GEN_842 = branchOps_valid ? _GEN_778 : _GEN_634; // @[utils.scala 59:26]
  wire [4:0] _GEN_843 = branchOps_valid ? _GEN_779 : _GEN_635; // @[utils.scala 59:26]
  wire [4:0] _GEN_844 = branchOps_valid ? _GEN_780 : _GEN_636; // @[utils.scala 59:26]
  wire [4:0] _GEN_845 = branchOps_valid ? _GEN_781 : _GEN_637; // @[utils.scala 59:26]
  wire  _GEN_846 = branchOps_valid ? _GEN_782 : _GEN_654; // @[utils.scala 59:26]
  wire  _GEN_847 = branchOps_valid ? _GEN_783 : _GEN_655; // @[utils.scala 59:26]
  wire  _GEN_848 = branchOps_valid ? _GEN_784 : _GEN_656; // @[utils.scala 59:26]
  wire  _GEN_849 = branchOps_valid ? _GEN_785 : _GEN_657; // @[utils.scala 59:26]
  wire  _GEN_850 = branchOps_valid ? _GEN_786 : _GEN_658; // @[utils.scala 59:26]
  wire  _GEN_851 = branchOps_valid ? _GEN_787 : _GEN_659; // @[utils.scala 59:26]
  wire  _GEN_852 = branchOps_valid ? _GEN_788 : _GEN_660; // @[utils.scala 59:26]
  wire  _GEN_853 = branchOps_valid ? _GEN_789 : _GEN_661; // @[utils.scala 59:26]
  wire  _GEN_854 = branchOps_valid ? _GEN_790 : _GEN_662; // @[utils.scala 59:26]
  wire  _GEN_855 = branchOps_valid ? _GEN_791 : _GEN_663; // @[utils.scala 59:26]
  wire  _GEN_856 = branchOps_valid ? _GEN_792 : _GEN_664; // @[utils.scala 59:26]
  wire  _GEN_857 = branchOps_valid ? _GEN_793 : _GEN_665; // @[utils.scala 59:26]
  wire  _GEN_858 = branchOps_valid ? _GEN_794 : _GEN_666; // @[utils.scala 59:26]
  wire  _GEN_859 = branchOps_valid ? _GEN_795 : _GEN_667; // @[utils.scala 59:26]
  wire  _GEN_860 = branchOps_valid ? _GEN_796 : _GEN_668; // @[utils.scala 59:26]
  wire  _GEN_861 = branchOps_valid ? _GEN_797 : _GEN_669; // @[utils.scala 59:26]
  wire [4:0] _GEN_862 = incrWrite ? _GEN_830 : _GEN_318; // @[fifo.scala 97:16]
  wire [4:0] _GEN_863 = incrWrite ? _GEN_831 : _GEN_319; // @[fifo.scala 97:16]
  wire [4:0] _GEN_864 = incrWrite ? _GEN_832 : _GEN_320; // @[fifo.scala 97:16]
  wire [4:0] _GEN_865 = incrWrite ? _GEN_833 : _GEN_321; // @[fifo.scala 97:16]
  wire [4:0] _GEN_866 = incrWrite ? _GEN_834 : _GEN_322; // @[fifo.scala 97:16]
  wire [4:0] _GEN_867 = incrWrite ? _GEN_835 : _GEN_323; // @[fifo.scala 97:16]
  wire [4:0] _GEN_868 = incrWrite ? _GEN_836 : _GEN_324; // @[fifo.scala 97:16]
  wire [4:0] _GEN_869 = incrWrite ? _GEN_837 : _GEN_325; // @[fifo.scala 97:16]
  wire [4:0] _GEN_870 = incrWrite ? _GEN_838 : _GEN_326; // @[fifo.scala 97:16]
  wire [4:0] _GEN_871 = incrWrite ? _GEN_839 : _GEN_327; // @[fifo.scala 97:16]
  wire [4:0] _GEN_872 = incrWrite ? _GEN_840 : _GEN_328; // @[fifo.scala 97:16]
  wire [4:0] _GEN_873 = incrWrite ? _GEN_841 : _GEN_329; // @[fifo.scala 97:16]
  wire [4:0] _GEN_874 = incrWrite ? _GEN_842 : _GEN_330; // @[fifo.scala 97:16]
  wire [4:0] _GEN_875 = incrWrite ? _GEN_843 : _GEN_331; // @[fifo.scala 97:16]
  wire [4:0] _GEN_876 = incrWrite ? _GEN_844 : _GEN_332; // @[fifo.scala 97:16]
  wire [4:0] _GEN_877 = incrWrite ? _GEN_845 : _GEN_333; // @[fifo.scala 97:16]
  wire  _GEN_878 = incrWrite ? _GEN_846 : _GEN_302; // @[fifo.scala 97:16]
  wire  _GEN_879 = incrWrite ? _GEN_847 : _GEN_303; // @[fifo.scala 97:16]
  wire  _GEN_880 = incrWrite ? _GEN_848 : _GEN_304; // @[fifo.scala 97:16]
  wire  _GEN_881 = incrWrite ? _GEN_849 : _GEN_305; // @[fifo.scala 97:16]
  wire  _GEN_882 = incrWrite ? _GEN_850 : _GEN_306; // @[fifo.scala 97:16]
  wire  _GEN_883 = incrWrite ? _GEN_851 : _GEN_307; // @[fifo.scala 97:16]
  wire  _GEN_884 = incrWrite ? _GEN_852 : _GEN_308; // @[fifo.scala 97:16]
  wire  _GEN_885 = incrWrite ? _GEN_853 : _GEN_309; // @[fifo.scala 97:16]
  wire  _GEN_886 = incrWrite ? _GEN_854 : _GEN_310; // @[fifo.scala 97:16]
  wire  _GEN_887 = incrWrite ? _GEN_855 : _GEN_311; // @[fifo.scala 97:16]
  wire  _GEN_888 = incrWrite ? _GEN_856 : _GEN_312; // @[fifo.scala 97:16]
  wire  _GEN_889 = incrWrite ? _GEN_857 : _GEN_313; // @[fifo.scala 97:16]
  wire  _GEN_890 = incrWrite ? _GEN_858 : _GEN_314; // @[fifo.scala 97:16]
  wire  _GEN_891 = incrWrite ? _GEN_859 : _GEN_315; // @[fifo.scala 97:16]
  wire  _GEN_892 = incrWrite ? _GEN_860 : _GEN_316; // @[fifo.scala 97:16]
  wire  _GEN_893 = incrWrite ? _GEN_861 : _GEN_317; // @[fifo.scala 97:16]
  wire [3:0] startPointer = read_ready ? _nextVal_T_2 : readPtr; // @[fifo.scala 102:25]
  wire [3:0] endPointer = writePtr - 4'h1; // @[fifo.scala 103:29]
  wire [4:0] _T_15 = memReg_0_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_16 = |_T_15; // @[fifo.scala 109:63]
  wire [4:0] _memReg_0_branch_mask_T = memReg_0_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _T_22 = memReg_1_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_23 = |_T_22; // @[fifo.scala 109:63]
  wire [4:0] _memReg_1_branch_mask_T = memReg_1_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_900 = |_T_22 ? _memReg_1_branch_mask_T : _GEN_863; // @[fifo.scala 109:68 110:35]
  wire  _GEN_901 = _T_23 ? 1'h0 : _GEN_879; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_29 = memReg_2_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_30 = |_T_29; // @[fifo.scala 109:63]
  wire [4:0] _memReg_2_branch_mask_T = memReg_2_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_906 = |_T_29 ? _memReg_2_branch_mask_T : _GEN_864; // @[fifo.scala 109:68 110:35]
  wire  _GEN_907 = _T_30 ? 1'h0 : _GEN_880; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_36 = memReg_3_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_37 = |_T_36; // @[fifo.scala 109:63]
  wire [4:0] _memReg_3_branch_mask_T = memReg_3_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_912 = |_T_36 ? _memReg_3_branch_mask_T : _GEN_865; // @[fifo.scala 109:68 110:35]
  wire  _GEN_913 = _T_37 ? 1'h0 : _GEN_881; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_43 = memReg_4_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_44 = |_T_43; // @[fifo.scala 109:63]
  wire [4:0] _memReg_4_branch_mask_T = memReg_4_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_918 = |_T_43 ? _memReg_4_branch_mask_T : _GEN_866; // @[fifo.scala 109:68 110:35]
  wire  _GEN_919 = _T_44 ? 1'h0 : _GEN_882; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_50 = memReg_5_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_51 = |_T_50; // @[fifo.scala 109:63]
  wire [4:0] _memReg_5_branch_mask_T = memReg_5_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_924 = |_T_50 ? _memReg_5_branch_mask_T : _GEN_867; // @[fifo.scala 109:68 110:35]
  wire  _GEN_925 = _T_51 ? 1'h0 : _GEN_883; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_57 = memReg_6_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_58 = |_T_57; // @[fifo.scala 109:63]
  wire [4:0] _memReg_6_branch_mask_T = memReg_6_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_930 = |_T_57 ? _memReg_6_branch_mask_T : _GEN_868; // @[fifo.scala 109:68 110:35]
  wire  _GEN_931 = _T_58 ? 1'h0 : _GEN_884; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_64 = memReg_7_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_65 = |_T_64; // @[fifo.scala 109:63]
  wire [4:0] _memReg_7_branch_mask_T = memReg_7_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_936 = |_T_64 ? _memReg_7_branch_mask_T : _GEN_869; // @[fifo.scala 109:68 110:35]
  wire  _GEN_937 = _T_65 ? 1'h0 : _GEN_885; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_71 = memReg_8_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_72 = |_T_71; // @[fifo.scala 109:63]
  wire [4:0] _memReg_8_branch_mask_T = memReg_8_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_942 = |_T_71 ? _memReg_8_branch_mask_T : _GEN_870; // @[fifo.scala 109:68 110:35]
  wire  _GEN_943 = _T_72 ? 1'h0 : _GEN_886; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_78 = memReg_9_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_79 = |_T_78; // @[fifo.scala 109:63]
  wire [4:0] _memReg_9_branch_mask_T = memReg_9_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_948 = |_T_78 ? _memReg_9_branch_mask_T : _GEN_871; // @[fifo.scala 109:68 110:35]
  wire  _GEN_949 = _T_79 ? 1'h0 : _GEN_887; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_85 = memReg_10_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_86 = |_T_85; // @[fifo.scala 109:63]
  wire [4:0] _memReg_10_branch_mask_T = memReg_10_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_954 = |_T_85 ? _memReg_10_branch_mask_T : _GEN_872; // @[fifo.scala 109:68 110:35]
  wire  _GEN_955 = _T_86 ? 1'h0 : _GEN_888; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_92 = memReg_11_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_93 = |_T_92; // @[fifo.scala 109:63]
  wire [4:0] _memReg_11_branch_mask_T = memReg_11_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_960 = |_T_92 ? _memReg_11_branch_mask_T : _GEN_873; // @[fifo.scala 109:68 110:35]
  wire  _GEN_961 = _T_93 ? 1'h0 : _GEN_889; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_99 = memReg_12_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_100 = |_T_99; // @[fifo.scala 109:63]
  wire [4:0] _memReg_12_branch_mask_T = memReg_12_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_966 = |_T_99 ? _memReg_12_branch_mask_T : _GEN_874; // @[fifo.scala 109:68 110:35]
  wire  _GEN_967 = _T_100 ? 1'h0 : _GEN_890; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_106 = memReg_13_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_107 = |_T_106; // @[fifo.scala 109:63]
  wire [4:0] _memReg_13_branch_mask_T = memReg_13_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_972 = |_T_106 ? _memReg_13_branch_mask_T : _GEN_875; // @[fifo.scala 109:68 110:35]
  wire  _GEN_973 = _T_107 ? 1'h0 : _GEN_891; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_113 = memReg_14_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_114 = |_T_113; // @[fifo.scala 109:63]
  wire [4:0] _memReg_14_branch_mask_T = memReg_14_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_978 = |_T_113 ? _memReg_14_branch_mask_T : _GEN_876; // @[fifo.scala 109:68 110:35]
  wire  _GEN_979 = _T_114 ? 1'h0 : _GEN_892; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_120 = memReg_15_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_121 = |_T_120; // @[fifo.scala 109:63]
  wire [4:0] _memReg_15_branch_mask_T = memReg_15_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _T_124 = _GEN_525 & branchOps_branchMask; // @[utils.scala 92:27]
  wire  _T_125 = |_T_124; // @[utils.scala 92:51]
  wire [4:0] _read_data_branch_mask_T = _GEN_525 ^ branchOps_branchMask; // @[utils.scala 93:42]
  wire [4:0] _GEN_1022 = |_T_124 ? _read_data_branch_mask_T : _GEN_525; // @[utils.scala 92:56 93:27 96:27]
  wire [4:0] _GEN_1023 = _T_125 ? 5'h0 : _GEN_525; // @[utils.scala 101:56 102:27 106:27]
  wire  _GEN_1024 = _T_125 ? 1'h0 : _GEN_509; // @[utils.scala 101:56 103:28 107:28]
  wire [4:0] _GEN_1025 = branchOps_passed ? _GEN_1022 : _GEN_1023; // @[utils.scala 90:30]
  wire  _GEN_1026 = branchOps_passed ? _GEN_509 : _GEN_1024; // @[utils.scala 90:30 98:26]
  wire  _matchFound_T_3 = memReg_0_valid & memReg_0_address[31:3] == checkAddress[31:3]; // @[fifo.scala 132:26]
  wire  _matchFound_T_7 = memReg_1_valid & memReg_1_address[31:3] == checkAddress[31:3]; // @[fifo.scala 132:26]
  wire  _matchFound_T_11 = memReg_2_valid & memReg_2_address[31:3] == checkAddress[31:3]; // @[fifo.scala 132:26]
  wire  _matchFound_T_15 = memReg_3_valid & memReg_3_address[31:3] == checkAddress[31:3]; // @[fifo.scala 132:26]
  wire  _matchFound_T_19 = memReg_4_valid & memReg_4_address[31:3] == checkAddress[31:3]; // @[fifo.scala 132:26]
  wire  _matchFound_T_23 = memReg_5_valid & memReg_5_address[31:3] == checkAddress[31:3]; // @[fifo.scala 132:26]
  wire  _matchFound_T_27 = memReg_6_valid & memReg_6_address[31:3] == checkAddress[31:3]; // @[fifo.scala 132:26]
  wire  _matchFound_T_31 = memReg_7_valid & memReg_7_address[31:3] == checkAddress[31:3]; // @[fifo.scala 132:26]
  wire  _matchFound_T_35 = memReg_8_valid & memReg_8_address[31:3] == checkAddress[31:3]; // @[fifo.scala 132:26]
  wire  _matchFound_T_39 = memReg_9_valid & memReg_9_address[31:3] == checkAddress[31:3]; // @[fifo.scala 132:26]
  wire  _matchFound_T_43 = memReg_10_valid & memReg_10_address[31:3] == checkAddress[31:3]; // @[fifo.scala 132:26]
  wire  _matchFound_T_47 = memReg_11_valid & memReg_11_address[31:3] == checkAddress[31:3]; // @[fifo.scala 132:26]
  wire  _matchFound_T_51 = memReg_12_valid & memReg_12_address[31:3] == checkAddress[31:3]; // @[fifo.scala 132:26]
  wire  _matchFound_T_55 = memReg_13_valid & memReg_13_address[31:3] == checkAddress[31:3]; // @[fifo.scala 132:26]
  wire  _matchFound_T_59 = memReg_14_valid & memReg_14_address[31:3] == checkAddress[31:3]; // @[fifo.scala 132:26]
  wire  _matchFound_T_63 = memReg_15_valid & memReg_15_address[31:3] == checkAddress[31:3]; // @[fifo.scala 132:26]
  assign write_ready = ~fullReg; // @[fifo.scala 88:18]
  assign read_data_valid = _T_2 & _GEN_429; // @[fifo.scala 122:32]
  assign read_data_address = 4'hf == readPtr ? memReg_15_address : _GEN_444; // @[fifo.scala 86:{13,13}]
  assign read_data_core_instruction = 4'hf == readPtr ? memReg_15_core_instruction : _GEN_460; // @[fifo.scala 86:{13,13}]
  assign read_data_core_robAddr = 4'hf == readPtr ? memReg_15_core_robAddr : _GEN_476; // @[fifo.scala 86:{13,13}]
  assign read_data_core_prfDest = 4'hf == readPtr ? memReg_15_core_prfDest : _GEN_492; // @[fifo.scala 86:{13,13}]
  assign read_data_branch_valid = branchOps_valid ? _GEN_1026 : _GEN_509; // @[utils.scala 112:24 89:27]
  assign read_data_branch_mask = branchOps_valid ? _GEN_1025 : _GEN_525; // @[utils.scala 111:23 89:27]
  assign isEmpty = emptyReg; // @[fifo.scala 89:11]
  assign matchFound = _matchFound_T_3 | _matchFound_T_7 | _matchFound_T_11 | _matchFound_T_15 | _matchFound_T_19 |
    _matchFound_T_23 | _matchFound_T_27 | _matchFound_T_31 | _matchFound_T_35 | _matchFound_T_39 | _matchFound_T_43 |
    _matchFound_T_47 | _matchFound_T_51 | _matchFound_T_55 | _matchFound_T_59 | _matchFound_T_63; // @[fifo.scala 133:16]
  always @(posedge clock) begin
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (branchOps_passed) begin // @[fifo.scala 108:32]
        memReg_0_branch_valid <= _GEN_878;
      end else if (_T_16) begin // @[fifo.scala 113:68]
        memReg_0_branch_valid <= 1'h0; // @[fifo.scala 114:36]
      end else begin
        memReg_0_branch_valid <= _GEN_878;
      end
    end else begin
      memReg_0_branch_valid <= _GEN_878;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (branchOps_passed) begin // @[fifo.scala 108:32]
        if (|_T_15) begin // @[fifo.scala 109:68]
          memReg_0_branch_mask <= _memReg_0_branch_mask_T; // @[fifo.scala 110:35]
        end else begin
          memReg_0_branch_mask <= _GEN_862;
        end
      end else begin
        memReg_0_branch_mask <= _GEN_862;
      end
    end else begin
      memReg_0_branch_mask <= _GEN_862;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h1 | 4'h1 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_1_branch_valid <= _GEN_879;
        end else begin
          memReg_1_branch_valid <= _GEN_901;
        end
      end else begin
        memReg_1_branch_valid <= _GEN_879;
      end
    end else begin
      memReg_1_branch_valid <= _GEN_879;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h1 | 4'h1 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_1_branch_mask <= _GEN_900;
        end else begin
          memReg_1_branch_mask <= _GEN_863;
        end
      end else begin
        memReg_1_branch_mask <= _GEN_863;
      end
    end else begin
      memReg_1_branch_mask <= _GEN_863;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h2 | 4'h2 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_2_branch_valid <= _GEN_880;
        end else begin
          memReg_2_branch_valid <= _GEN_907;
        end
      end else begin
        memReg_2_branch_valid <= _GEN_880;
      end
    end else begin
      memReg_2_branch_valid <= _GEN_880;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h2 | 4'h2 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_2_branch_mask <= _GEN_906;
        end else begin
          memReg_2_branch_mask <= _GEN_864;
        end
      end else begin
        memReg_2_branch_mask <= _GEN_864;
      end
    end else begin
      memReg_2_branch_mask <= _GEN_864;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h3 | 4'h3 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_3_branch_valid <= _GEN_881;
        end else begin
          memReg_3_branch_valid <= _GEN_913;
        end
      end else begin
        memReg_3_branch_valid <= _GEN_881;
      end
    end else begin
      memReg_3_branch_valid <= _GEN_881;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h3 | 4'h3 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_3_branch_mask <= _GEN_912;
        end else begin
          memReg_3_branch_mask <= _GEN_865;
        end
      end else begin
        memReg_3_branch_mask <= _GEN_865;
      end
    end else begin
      memReg_3_branch_mask <= _GEN_865;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h4 | 4'h4 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_4_branch_valid <= _GEN_882;
        end else begin
          memReg_4_branch_valid <= _GEN_919;
        end
      end else begin
        memReg_4_branch_valid <= _GEN_882;
      end
    end else begin
      memReg_4_branch_valid <= _GEN_882;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h4 | 4'h4 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_4_branch_mask <= _GEN_918;
        end else begin
          memReg_4_branch_mask <= _GEN_866;
        end
      end else begin
        memReg_4_branch_mask <= _GEN_866;
      end
    end else begin
      memReg_4_branch_mask <= _GEN_866;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h5 | 4'h5 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_5_branch_valid <= _GEN_883;
        end else begin
          memReg_5_branch_valid <= _GEN_925;
        end
      end else begin
        memReg_5_branch_valid <= _GEN_883;
      end
    end else begin
      memReg_5_branch_valid <= _GEN_883;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h5 | 4'h5 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_5_branch_mask <= _GEN_924;
        end else begin
          memReg_5_branch_mask <= _GEN_867;
        end
      end else begin
        memReg_5_branch_mask <= _GEN_867;
      end
    end else begin
      memReg_5_branch_mask <= _GEN_867;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h6 | 4'h6 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_6_branch_valid <= _GEN_884;
        end else begin
          memReg_6_branch_valid <= _GEN_931;
        end
      end else begin
        memReg_6_branch_valid <= _GEN_884;
      end
    end else begin
      memReg_6_branch_valid <= _GEN_884;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h6 | 4'h6 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_6_branch_mask <= _GEN_930;
        end else begin
          memReg_6_branch_mask <= _GEN_868;
        end
      end else begin
        memReg_6_branch_mask <= _GEN_868;
      end
    end else begin
      memReg_6_branch_mask <= _GEN_868;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h7 | 4'h7 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_7_branch_valid <= _GEN_885;
        end else begin
          memReg_7_branch_valid <= _GEN_937;
        end
      end else begin
        memReg_7_branch_valid <= _GEN_885;
      end
    end else begin
      memReg_7_branch_valid <= _GEN_885;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h7 | 4'h7 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_7_branch_mask <= _GEN_936;
        end else begin
          memReg_7_branch_mask <= _GEN_869;
        end
      end else begin
        memReg_7_branch_mask <= _GEN_869;
      end
    end else begin
      memReg_7_branch_mask <= _GEN_869;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h8 | 4'h8 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_8_branch_valid <= _GEN_886;
        end else begin
          memReg_8_branch_valid <= _GEN_943;
        end
      end else begin
        memReg_8_branch_valid <= _GEN_886;
      end
    end else begin
      memReg_8_branch_valid <= _GEN_886;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h8 | 4'h8 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_8_branch_mask <= _GEN_942;
        end else begin
          memReg_8_branch_mask <= _GEN_870;
        end
      end else begin
        memReg_8_branch_mask <= _GEN_870;
      end
    end else begin
      memReg_8_branch_mask <= _GEN_870;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h9 | 4'h9 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_9_branch_valid <= _GEN_887;
        end else begin
          memReg_9_branch_valid <= _GEN_949;
        end
      end else begin
        memReg_9_branch_valid <= _GEN_887;
      end
    end else begin
      memReg_9_branch_valid <= _GEN_887;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h9 | 4'h9 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_9_branch_mask <= _GEN_948;
        end else begin
          memReg_9_branch_mask <= _GEN_871;
        end
      end else begin
        memReg_9_branch_mask <= _GEN_871;
      end
    end else begin
      memReg_9_branch_mask <= _GEN_871;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'ha | 4'ha <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_10_branch_valid <= _GEN_888;
        end else begin
          memReg_10_branch_valid <= _GEN_955;
        end
      end else begin
        memReg_10_branch_valid <= _GEN_888;
      end
    end else begin
      memReg_10_branch_valid <= _GEN_888;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'ha | 4'ha <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_10_branch_mask <= _GEN_954;
        end else begin
          memReg_10_branch_mask <= _GEN_872;
        end
      end else begin
        memReg_10_branch_mask <= _GEN_872;
      end
    end else begin
      memReg_10_branch_mask <= _GEN_872;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'hb | 4'hb <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_11_branch_valid <= _GEN_889;
        end else begin
          memReg_11_branch_valid <= _GEN_961;
        end
      end else begin
        memReg_11_branch_valid <= _GEN_889;
      end
    end else begin
      memReg_11_branch_valid <= _GEN_889;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'hb | 4'hb <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_11_branch_mask <= _GEN_960;
        end else begin
          memReg_11_branch_mask <= _GEN_873;
        end
      end else begin
        memReg_11_branch_mask <= _GEN_873;
      end
    end else begin
      memReg_11_branch_mask <= _GEN_873;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'hc | 4'hc <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_12_branch_valid <= _GEN_890;
        end else begin
          memReg_12_branch_valid <= _GEN_967;
        end
      end else begin
        memReg_12_branch_valid <= _GEN_890;
      end
    end else begin
      memReg_12_branch_valid <= _GEN_890;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'hc | 4'hc <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_12_branch_mask <= _GEN_966;
        end else begin
          memReg_12_branch_mask <= _GEN_874;
        end
      end else begin
        memReg_12_branch_mask <= _GEN_874;
      end
    end else begin
      memReg_12_branch_mask <= _GEN_874;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'hd | 4'hd <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_13_branch_valid <= _GEN_891;
        end else begin
          memReg_13_branch_valid <= _GEN_973;
        end
      end else begin
        memReg_13_branch_valid <= _GEN_891;
      end
    end else begin
      memReg_13_branch_valid <= _GEN_891;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'hd | 4'hd <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_13_branch_mask <= _GEN_972;
        end else begin
          memReg_13_branch_mask <= _GEN_875;
        end
      end else begin
        memReg_13_branch_mask <= _GEN_875;
      end
    end else begin
      memReg_13_branch_mask <= _GEN_875;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'he | 4'he <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_14_branch_valid <= _GEN_892;
        end else begin
          memReg_14_branch_valid <= _GEN_979;
        end
      end else begin
        memReg_14_branch_valid <= _GEN_892;
      end
    end else begin
      memReg_14_branch_valid <= _GEN_892;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'he | 4'he <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_14_branch_mask <= _GEN_978;
        end else begin
          memReg_14_branch_mask <= _GEN_876;
        end
      end else begin
        memReg_14_branch_mask <= _GEN_876;
      end
    end else begin
      memReg_14_branch_mask <= _GEN_876;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (branchOps_passed) begin // @[fifo.scala 108:32]
        memReg_15_branch_valid <= _GEN_893;
      end else if (_T_121) begin // @[fifo.scala 113:68]
        memReg_15_branch_valid <= 1'h0; // @[fifo.scala 114:36]
      end else begin
        memReg_15_branch_valid <= _GEN_893;
      end
    end else begin
      memReg_15_branch_valid <= _GEN_893;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (branchOps_passed) begin // @[fifo.scala 108:32]
        if (|_T_120) begin // @[fifo.scala 109:68]
          memReg_15_branch_mask <= _memReg_15_branch_mask_T; // @[fifo.scala 110:35]
        end else begin
          memReg_15_branch_mask <= _GEN_877;
        end
      end else begin
        memReg_15_branch_mask <= _GEN_877;
      end
    end else begin
      memReg_15_branch_mask <= _GEN_877;
    end
    if (reset) begin // @[fifo.scala 33:25]
      readPtr <= 4'h0; // @[fifo.scala 33:25]
    end else if (incrRead) begin // @[fifo.scala 35:15]
      if (readPtr == 4'hf) begin // @[fifo.scala 34:22]
        readPtr <= 4'h0;
      end else begin
        readPtr <= _nextVal_T_2;
      end
    end
    emptyReg <= reset | _GEN_27; // @[fifo.scala 43:{25,25}]
    if (reset) begin // @[fifo.scala 33:25]
      writePtr <= 4'h0; // @[fifo.scala 33:25]
    end else if (incrWrite) begin // @[fifo.scala 35:15]
      if (writePtr == 4'hf) begin // @[fifo.scala 34:22]
        writePtr <= 4'h0;
      end else begin
        writePtr <= _nextVal_T_5;
      end
    end
    if (reset) begin // @[fifo.scala 44:34]
      fullReg <= 1'h0; // @[fifo.scala 44:34]
    end else if (!(2'h0 == op)) begin // @[fifo.scala 49:14]
      if (2'h1 == op) begin // @[fifo.scala 49:14]
        if (~emptyReg) begin // @[fifo.scala 52:23]
          fullReg <= 1'h0; // @[fifo.scala 53:17]
        end
      end else if (2'h2 == op) begin // @[fifo.scala 49:14]
        fullReg <= _GEN_7;
      end else begin
        fullReg <= _GEN_16;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  memReg_0_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  memReg_0_address = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  memReg_0_core_instruction = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  memReg_0_core_robAddr = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  memReg_0_core_prfDest = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  memReg_0_branch_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  memReg_0_branch_mask = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  memReg_1_valid = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  memReg_1_address = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  memReg_1_core_instruction = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  memReg_1_core_robAddr = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  memReg_1_core_prfDest = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  memReg_1_branch_valid = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  memReg_1_branch_mask = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  memReg_2_valid = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  memReg_2_address = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  memReg_2_core_instruction = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  memReg_2_core_robAddr = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  memReg_2_core_prfDest = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  memReg_2_branch_valid = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  memReg_2_branch_mask = _RAND_20[4:0];
  _RAND_21 = {1{`RANDOM}};
  memReg_3_valid = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  memReg_3_address = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  memReg_3_core_instruction = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  memReg_3_core_robAddr = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  memReg_3_core_prfDest = _RAND_25[5:0];
  _RAND_26 = {1{`RANDOM}};
  memReg_3_branch_valid = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  memReg_3_branch_mask = _RAND_27[4:0];
  _RAND_28 = {1{`RANDOM}};
  memReg_4_valid = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  memReg_4_address = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  memReg_4_core_instruction = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  memReg_4_core_robAddr = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  memReg_4_core_prfDest = _RAND_32[5:0];
  _RAND_33 = {1{`RANDOM}};
  memReg_4_branch_valid = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  memReg_4_branch_mask = _RAND_34[4:0];
  _RAND_35 = {1{`RANDOM}};
  memReg_5_valid = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  memReg_5_address = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  memReg_5_core_instruction = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  memReg_5_core_robAddr = _RAND_38[3:0];
  _RAND_39 = {1{`RANDOM}};
  memReg_5_core_prfDest = _RAND_39[5:0];
  _RAND_40 = {1{`RANDOM}};
  memReg_5_branch_valid = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  memReg_5_branch_mask = _RAND_41[4:0];
  _RAND_42 = {1{`RANDOM}};
  memReg_6_valid = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  memReg_6_address = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  memReg_6_core_instruction = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  memReg_6_core_robAddr = _RAND_45[3:0];
  _RAND_46 = {1{`RANDOM}};
  memReg_6_core_prfDest = _RAND_46[5:0];
  _RAND_47 = {1{`RANDOM}};
  memReg_6_branch_valid = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  memReg_6_branch_mask = _RAND_48[4:0];
  _RAND_49 = {1{`RANDOM}};
  memReg_7_valid = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  memReg_7_address = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  memReg_7_core_instruction = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  memReg_7_core_robAddr = _RAND_52[3:0];
  _RAND_53 = {1{`RANDOM}};
  memReg_7_core_prfDest = _RAND_53[5:0];
  _RAND_54 = {1{`RANDOM}};
  memReg_7_branch_valid = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  memReg_7_branch_mask = _RAND_55[4:0];
  _RAND_56 = {1{`RANDOM}};
  memReg_8_valid = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  memReg_8_address = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  memReg_8_core_instruction = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  memReg_8_core_robAddr = _RAND_59[3:0];
  _RAND_60 = {1{`RANDOM}};
  memReg_8_core_prfDest = _RAND_60[5:0];
  _RAND_61 = {1{`RANDOM}};
  memReg_8_branch_valid = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  memReg_8_branch_mask = _RAND_62[4:0];
  _RAND_63 = {1{`RANDOM}};
  memReg_9_valid = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  memReg_9_address = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  memReg_9_core_instruction = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  memReg_9_core_robAddr = _RAND_66[3:0];
  _RAND_67 = {1{`RANDOM}};
  memReg_9_core_prfDest = _RAND_67[5:0];
  _RAND_68 = {1{`RANDOM}};
  memReg_9_branch_valid = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  memReg_9_branch_mask = _RAND_69[4:0];
  _RAND_70 = {1{`RANDOM}};
  memReg_10_valid = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  memReg_10_address = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  memReg_10_core_instruction = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  memReg_10_core_robAddr = _RAND_73[3:0];
  _RAND_74 = {1{`RANDOM}};
  memReg_10_core_prfDest = _RAND_74[5:0];
  _RAND_75 = {1{`RANDOM}};
  memReg_10_branch_valid = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  memReg_10_branch_mask = _RAND_76[4:0];
  _RAND_77 = {1{`RANDOM}};
  memReg_11_valid = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  memReg_11_address = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  memReg_11_core_instruction = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  memReg_11_core_robAddr = _RAND_80[3:0];
  _RAND_81 = {1{`RANDOM}};
  memReg_11_core_prfDest = _RAND_81[5:0];
  _RAND_82 = {1{`RANDOM}};
  memReg_11_branch_valid = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  memReg_11_branch_mask = _RAND_83[4:0];
  _RAND_84 = {1{`RANDOM}};
  memReg_12_valid = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  memReg_12_address = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  memReg_12_core_instruction = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  memReg_12_core_robAddr = _RAND_87[3:0];
  _RAND_88 = {1{`RANDOM}};
  memReg_12_core_prfDest = _RAND_88[5:0];
  _RAND_89 = {1{`RANDOM}};
  memReg_12_branch_valid = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  memReg_12_branch_mask = _RAND_90[4:0];
  _RAND_91 = {1{`RANDOM}};
  memReg_13_valid = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  memReg_13_address = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  memReg_13_core_instruction = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  memReg_13_core_robAddr = _RAND_94[3:0];
  _RAND_95 = {1{`RANDOM}};
  memReg_13_core_prfDest = _RAND_95[5:0];
  _RAND_96 = {1{`RANDOM}};
  memReg_13_branch_valid = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  memReg_13_branch_mask = _RAND_97[4:0];
  _RAND_98 = {1{`RANDOM}};
  memReg_14_valid = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  memReg_14_address = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  memReg_14_core_instruction = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  memReg_14_core_robAddr = _RAND_101[3:0];
  _RAND_102 = {1{`RANDOM}};
  memReg_14_core_prfDest = _RAND_102[5:0];
  _RAND_103 = {1{`RANDOM}};
  memReg_14_branch_valid = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  memReg_14_branch_mask = _RAND_104[4:0];
  _RAND_105 = {1{`RANDOM}};
  memReg_15_valid = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  memReg_15_address = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  memReg_15_core_instruction = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  memReg_15_core_robAddr = _RAND_108[3:0];
  _RAND_109 = {1{`RANDOM}};
  memReg_15_core_prfDest = _RAND_109[5:0];
  _RAND_110 = {1{`RANDOM}};
  memReg_15_branch_valid = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  memReg_15_branch_mask = _RAND_111[4:0];
  _RAND_112 = {1{`RANDOM}};
  readPtr = _RAND_112[3:0];
  _RAND_113 = {1{`RANDOM}};
  emptyReg = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  writePtr = _RAND_114[3:0];
  _RAND_115 = {1{`RANDOM}};
  fullReg = _RAND_115[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module fifoWithBranchOps(
  input         clock,
  input         reset,
  output        write_ready,
  input         write_data_valid,
  input  [31:0] write_data_address,
  input  [31:0] write_data_core_instruction,
  input  [3:0]  write_data_core_robAddr,
  input  [5:0]  write_data_core_prfDest,
  input         write_data_branch_valid,
  input  [4:0]  write_data_branch_mask,
  input         write_data_writeData_valid,
  input  [63:0] write_data_writeData_data,
  input  [1:0]  write_data_cacheLine_response,
  input         read_ready,
  output        read_data_valid,
  output [31:0] read_data_address,
  output [31:0] read_data_core_instruction,
  output [3:0]  read_data_core_robAddr,
  output [5:0]  read_data_core_prfDest,
  output        read_data_branch_valid,
  output [4:0]  read_data_branch_mask,
  output        read_data_writeData_valid,
  output [63:0] read_data_writeData_data,
  output [1:0]  read_data_cacheLine_response,
  output        isEmpty,
  input         branchOps_valid,
  input  [4:0]  branchOps_branchMask,
  input         branchOps_passed
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [63:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [63:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [63:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [63:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
`endif // RANDOMIZE_REG_INIT
  reg  memReg_0_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_0_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_0_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_0_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_0_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_0_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_0_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_0_writeData_valid; // @[fifo.scala 27:33]
  reg [63:0] memReg_0_writeData_data; // @[fifo.scala 27:33]
  reg [1:0] memReg_0_cacheLine_response; // @[fifo.scala 27:33]
  reg  memReg_1_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_1_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_1_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_1_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_1_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_1_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_1_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_1_writeData_valid; // @[fifo.scala 27:33]
  reg [63:0] memReg_1_writeData_data; // @[fifo.scala 27:33]
  reg [1:0] memReg_1_cacheLine_response; // @[fifo.scala 27:33]
  reg  memReg_2_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_2_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_2_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_2_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_2_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_2_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_2_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_2_writeData_valid; // @[fifo.scala 27:33]
  reg [63:0] memReg_2_writeData_data; // @[fifo.scala 27:33]
  reg [1:0] memReg_2_cacheLine_response; // @[fifo.scala 27:33]
  reg  memReg_3_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_3_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_3_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_3_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_3_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_3_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_3_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_3_writeData_valid; // @[fifo.scala 27:33]
  reg [63:0] memReg_3_writeData_data; // @[fifo.scala 27:33]
  reg [1:0] memReg_3_cacheLine_response; // @[fifo.scala 27:33]
  reg  memReg_4_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_4_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_4_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_4_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_4_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_4_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_4_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_4_writeData_valid; // @[fifo.scala 27:33]
  reg [63:0] memReg_4_writeData_data; // @[fifo.scala 27:33]
  reg [1:0] memReg_4_cacheLine_response; // @[fifo.scala 27:33]
  reg  memReg_5_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_5_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_5_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_5_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_5_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_5_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_5_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_5_writeData_valid; // @[fifo.scala 27:33]
  reg [63:0] memReg_5_writeData_data; // @[fifo.scala 27:33]
  reg [1:0] memReg_5_cacheLine_response; // @[fifo.scala 27:33]
  reg  memReg_6_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_6_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_6_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_6_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_6_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_6_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_6_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_6_writeData_valid; // @[fifo.scala 27:33]
  reg [63:0] memReg_6_writeData_data; // @[fifo.scala 27:33]
  reg [1:0] memReg_6_cacheLine_response; // @[fifo.scala 27:33]
  reg  memReg_7_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_7_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_7_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_7_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_7_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_7_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_7_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_7_writeData_valid; // @[fifo.scala 27:33]
  reg [63:0] memReg_7_writeData_data; // @[fifo.scala 27:33]
  reg [1:0] memReg_7_cacheLine_response; // @[fifo.scala 27:33]
  reg  memReg_8_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_8_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_8_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_8_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_8_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_8_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_8_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_8_writeData_valid; // @[fifo.scala 27:33]
  reg [63:0] memReg_8_writeData_data; // @[fifo.scala 27:33]
  reg [1:0] memReg_8_cacheLine_response; // @[fifo.scala 27:33]
  reg  memReg_9_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_9_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_9_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_9_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_9_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_9_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_9_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_9_writeData_valid; // @[fifo.scala 27:33]
  reg [63:0] memReg_9_writeData_data; // @[fifo.scala 27:33]
  reg [1:0] memReg_9_cacheLine_response; // @[fifo.scala 27:33]
  reg  memReg_10_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_10_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_10_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_10_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_10_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_10_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_10_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_10_writeData_valid; // @[fifo.scala 27:33]
  reg [63:0] memReg_10_writeData_data; // @[fifo.scala 27:33]
  reg [1:0] memReg_10_cacheLine_response; // @[fifo.scala 27:33]
  reg  memReg_11_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_11_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_11_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_11_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_11_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_11_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_11_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_11_writeData_valid; // @[fifo.scala 27:33]
  reg [63:0] memReg_11_writeData_data; // @[fifo.scala 27:33]
  reg [1:0] memReg_11_cacheLine_response; // @[fifo.scala 27:33]
  reg  memReg_12_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_12_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_12_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_12_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_12_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_12_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_12_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_12_writeData_valid; // @[fifo.scala 27:33]
  reg [63:0] memReg_12_writeData_data; // @[fifo.scala 27:33]
  reg [1:0] memReg_12_cacheLine_response; // @[fifo.scala 27:33]
  reg  memReg_13_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_13_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_13_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_13_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_13_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_13_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_13_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_13_writeData_valid; // @[fifo.scala 27:33]
  reg [63:0] memReg_13_writeData_data; // @[fifo.scala 27:33]
  reg [1:0] memReg_13_cacheLine_response; // @[fifo.scala 27:33]
  reg  memReg_14_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_14_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_14_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_14_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_14_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_14_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_14_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_14_writeData_valid; // @[fifo.scala 27:33]
  reg [63:0] memReg_14_writeData_data; // @[fifo.scala 27:33]
  reg [1:0] memReg_14_cacheLine_response; // @[fifo.scala 27:33]
  reg  memReg_15_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_15_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_15_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_15_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_15_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_15_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_15_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_15_writeData_valid; // @[fifo.scala 27:33]
  reg [63:0] memReg_15_writeData_data; // @[fifo.scala 27:33]
  reg [1:0] memReg_15_cacheLine_response; // @[fifo.scala 27:33]
  reg [3:0] readPtr; // @[fifo.scala 33:25]
  wire [3:0] _nextVal_T_2 = readPtr + 4'h1; // @[fifo.scala 34:60]
  wire [3:0] nextRead = readPtr == 4'hf ? 4'h0 : _nextVal_T_2; // @[fifo.scala 34:22]
  wire [1:0] op = {write_data_valid,read_ready}; // @[fifo.scala 46:29]
  reg  emptyReg; // @[fifo.scala 43:25]
  wire  _T_2 = ~emptyReg; // @[fifo.scala 52:12]
  wire  _GEN_21 = 2'h2 == op ? 1'h0 : 2'h3 == op & _T_2; // @[fifo.scala 49:14]
  wire  _GEN_24 = 2'h1 == op ? _T_2 : _GEN_21; // @[fifo.scala 49:14]
  wire  incrRead = 2'h0 == op ? 1'h0 : _GEN_24; // @[fifo.scala 49:14]
  reg [3:0] writePtr; // @[fifo.scala 33:25]
  wire [3:0] _nextVal_T_5 = writePtr + 4'h1; // @[fifo.scala 34:60]
  wire [3:0] nextWrite = writePtr == 4'hf ? 4'h0 : _nextVal_T_5; // @[fifo.scala 34:22]
  reg  fullReg; // @[fifo.scala 44:34]
  wire  _T_4 = ~fullReg; // @[fifo.scala 59:12]
  wire  _GEN_18 = 2'h2 == op ? _T_4 : 2'h3 == op & _T_4; // @[fifo.scala 49:14]
  wire  _GEN_25 = 2'h1 == op ? 1'h0 : _GEN_18; // @[fifo.scala 49:14]
  wire  incrWrite = 2'h0 == op ? 1'h0 : _GEN_25; // @[fifo.scala 49:14]
  wire  _GEN_3 = ~emptyReg ? nextRead == writePtr : emptyReg; // @[fifo.scala 52:23 54:18 43:25]
  wire  _GEN_6 = ~fullReg ? 1'h0 : emptyReg; // @[fifo.scala 59:22 61:18 43:25]
  wire  _GEN_7 = ~fullReg ? nextWrite == readPtr : fullReg; // @[fifo.scala 59:22 62:17 44:34]
  wire  _fullReg_T_2 = emptyReg ? 1'h0 : nextWrite == nextRead; // @[fifo.scala 70:23]
  wire  _GEN_10 = _T_4 ? _fullReg_T_2 : fullReg; // @[fifo.scala 67:22 70:17 44:34]
  wire  _emptyReg_T_2 = fullReg ? 1'h0 : nextRead == nextWrite; // @[fifo.scala 75:24]
  wire  _GEN_11 = _T_2 ? 1'h0 : _GEN_10; // @[fifo.scala 73:23 74:17]
  wire  _GEN_12 = _T_2 ? _emptyReg_T_2 : _GEN_6; // @[fifo.scala 73:23 75:18]
  wire  _GEN_15 = 2'h3 == op ? _GEN_12 : emptyReg; // @[fifo.scala 49:14 43:25]
  wire  _GEN_16 = 2'h3 == op ? _GEN_11 : fullReg; // @[fifo.scala 49:14 44:34]
  wire  _GEN_19 = 2'h2 == op ? _GEN_6 : _GEN_15; // @[fifo.scala 49:14]
  wire  _GEN_23 = 2'h1 == op ? _GEN_3 : _GEN_19; // @[fifo.scala 49:14]
  wire  _GEN_27 = 2'h0 == op ? emptyReg : _GEN_23; // @[fifo.scala 49:14 43:25]
  wire  _GEN_110 = 4'h0 == writePtr ? write_data_branch_valid : memReg_0_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_111 = 4'h1 == writePtr ? write_data_branch_valid : memReg_1_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_112 = 4'h2 == writePtr ? write_data_branch_valid : memReg_2_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_113 = 4'h3 == writePtr ? write_data_branch_valid : memReg_3_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_114 = 4'h4 == writePtr ? write_data_branch_valid : memReg_4_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_115 = 4'h5 == writePtr ? write_data_branch_valid : memReg_5_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_116 = 4'h6 == writePtr ? write_data_branch_valid : memReg_6_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_117 = 4'h7 == writePtr ? write_data_branch_valid : memReg_7_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_118 = 4'h8 == writePtr ? write_data_branch_valid : memReg_8_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_119 = 4'h9 == writePtr ? write_data_branch_valid : memReg_9_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_120 = 4'ha == writePtr ? write_data_branch_valid : memReg_10_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_121 = 4'hb == writePtr ? write_data_branch_valid : memReg_11_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_122 = 4'hc == writePtr ? write_data_branch_valid : memReg_12_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_123 = 4'hd == writePtr ? write_data_branch_valid : memReg_13_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_124 = 4'he == writePtr ? write_data_branch_valid : memReg_14_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_125 = 4'hf == writePtr ? write_data_branch_valid : memReg_15_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_126 = 4'h0 == writePtr ? write_data_branch_mask : memReg_0_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_127 = 4'h1 == writePtr ? write_data_branch_mask : memReg_1_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_128 = 4'h2 == writePtr ? write_data_branch_mask : memReg_2_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_129 = 4'h3 == writePtr ? write_data_branch_mask : memReg_3_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_130 = 4'h4 == writePtr ? write_data_branch_mask : memReg_4_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_131 = 4'h5 == writePtr ? write_data_branch_mask : memReg_5_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_132 = 4'h6 == writePtr ? write_data_branch_mask : memReg_6_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_133 = 4'h7 == writePtr ? write_data_branch_mask : memReg_7_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_134 = 4'h8 == writePtr ? write_data_branch_mask : memReg_8_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_135 = 4'h9 == writePtr ? write_data_branch_mask : memReg_9_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_136 = 4'ha == writePtr ? write_data_branch_mask : memReg_10_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_137 = 4'hb == writePtr ? write_data_branch_mask : memReg_11_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_138 = 4'hc == writePtr ? write_data_branch_mask : memReg_12_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_139 = 4'hd == writePtr ? write_data_branch_mask : memReg_13_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_140 = 4'he == writePtr ? write_data_branch_mask : memReg_14_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_141 = 4'hf == writePtr ? write_data_branch_mask : memReg_15_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_302 = incrWrite ? _GEN_110 : memReg_0_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_303 = incrWrite ? _GEN_111 : memReg_1_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_304 = incrWrite ? _GEN_112 : memReg_2_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_305 = incrWrite ? _GEN_113 : memReg_3_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_306 = incrWrite ? _GEN_114 : memReg_4_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_307 = incrWrite ? _GEN_115 : memReg_5_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_308 = incrWrite ? _GEN_116 : memReg_6_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_309 = incrWrite ? _GEN_117 : memReg_7_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_310 = incrWrite ? _GEN_118 : memReg_8_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_311 = incrWrite ? _GEN_119 : memReg_9_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_312 = incrWrite ? _GEN_120 : memReg_10_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_313 = incrWrite ? _GEN_121 : memReg_11_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_314 = incrWrite ? _GEN_122 : memReg_12_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_315 = incrWrite ? _GEN_123 : memReg_13_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_316 = incrWrite ? _GEN_124 : memReg_14_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_317 = incrWrite ? _GEN_125 : memReg_15_branch_valid; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_318 = incrWrite ? _GEN_126 : memReg_0_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_319 = incrWrite ? _GEN_127 : memReg_1_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_320 = incrWrite ? _GEN_128 : memReg_2_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_321 = incrWrite ? _GEN_129 : memReg_3_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_322 = incrWrite ? _GEN_130 : memReg_4_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_323 = incrWrite ? _GEN_131 : memReg_5_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_324 = incrWrite ? _GEN_132 : memReg_6_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_325 = incrWrite ? _GEN_133 : memReg_7_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_326 = incrWrite ? _GEN_134 : memReg_8_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_327 = incrWrite ? _GEN_135 : memReg_9_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_328 = incrWrite ? _GEN_136 : memReg_10_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_329 = incrWrite ? _GEN_137 : memReg_11_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_330 = incrWrite ? _GEN_138 : memReg_12_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_331 = incrWrite ? _GEN_139 : memReg_13_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_332 = incrWrite ? _GEN_140 : memReg_14_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_333 = incrWrite ? _GEN_141 : memReg_15_branch_mask; // @[fifo.scala 81:17 27:33]
  wire  _GEN_415 = 4'h1 == readPtr ? memReg_1_valid : memReg_0_valid; // @[fifo.scala 86:{13,13}]
  wire  _GEN_416 = 4'h2 == readPtr ? memReg_2_valid : _GEN_415; // @[fifo.scala 86:{13,13}]
  wire  _GEN_417 = 4'h3 == readPtr ? memReg_3_valid : _GEN_416; // @[fifo.scala 86:{13,13}]
  wire  _GEN_418 = 4'h4 == readPtr ? memReg_4_valid : _GEN_417; // @[fifo.scala 86:{13,13}]
  wire  _GEN_419 = 4'h5 == readPtr ? memReg_5_valid : _GEN_418; // @[fifo.scala 86:{13,13}]
  wire  _GEN_420 = 4'h6 == readPtr ? memReg_6_valid : _GEN_419; // @[fifo.scala 86:{13,13}]
  wire  _GEN_421 = 4'h7 == readPtr ? memReg_7_valid : _GEN_420; // @[fifo.scala 86:{13,13}]
  wire  _GEN_422 = 4'h8 == readPtr ? memReg_8_valid : _GEN_421; // @[fifo.scala 86:{13,13}]
  wire  _GEN_423 = 4'h9 == readPtr ? memReg_9_valid : _GEN_422; // @[fifo.scala 86:{13,13}]
  wire  _GEN_424 = 4'ha == readPtr ? memReg_10_valid : _GEN_423; // @[fifo.scala 86:{13,13}]
  wire  _GEN_425 = 4'hb == readPtr ? memReg_11_valid : _GEN_424; // @[fifo.scala 86:{13,13}]
  wire  _GEN_426 = 4'hc == readPtr ? memReg_12_valid : _GEN_425; // @[fifo.scala 86:{13,13}]
  wire  _GEN_427 = 4'hd == readPtr ? memReg_13_valid : _GEN_426; // @[fifo.scala 86:{13,13}]
  wire  _GEN_428 = 4'he == readPtr ? memReg_14_valid : _GEN_427; // @[fifo.scala 86:{13,13}]
  wire  _GEN_429 = 4'hf == readPtr ? memReg_15_valid : _GEN_428; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_431 = 4'h1 == readPtr ? memReg_1_address : memReg_0_address; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_432 = 4'h2 == readPtr ? memReg_2_address : _GEN_431; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_433 = 4'h3 == readPtr ? memReg_3_address : _GEN_432; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_434 = 4'h4 == readPtr ? memReg_4_address : _GEN_433; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_435 = 4'h5 == readPtr ? memReg_5_address : _GEN_434; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_436 = 4'h6 == readPtr ? memReg_6_address : _GEN_435; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_437 = 4'h7 == readPtr ? memReg_7_address : _GEN_436; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_438 = 4'h8 == readPtr ? memReg_8_address : _GEN_437; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_439 = 4'h9 == readPtr ? memReg_9_address : _GEN_438; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_440 = 4'ha == readPtr ? memReg_10_address : _GEN_439; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_441 = 4'hb == readPtr ? memReg_11_address : _GEN_440; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_442 = 4'hc == readPtr ? memReg_12_address : _GEN_441; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_443 = 4'hd == readPtr ? memReg_13_address : _GEN_442; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_444 = 4'he == readPtr ? memReg_14_address : _GEN_443; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_447 = 4'h1 == readPtr ? memReg_1_core_instruction : memReg_0_core_instruction; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_448 = 4'h2 == readPtr ? memReg_2_core_instruction : _GEN_447; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_449 = 4'h3 == readPtr ? memReg_3_core_instruction : _GEN_448; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_450 = 4'h4 == readPtr ? memReg_4_core_instruction : _GEN_449; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_451 = 4'h5 == readPtr ? memReg_5_core_instruction : _GEN_450; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_452 = 4'h6 == readPtr ? memReg_6_core_instruction : _GEN_451; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_453 = 4'h7 == readPtr ? memReg_7_core_instruction : _GEN_452; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_454 = 4'h8 == readPtr ? memReg_8_core_instruction : _GEN_453; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_455 = 4'h9 == readPtr ? memReg_9_core_instruction : _GEN_454; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_456 = 4'ha == readPtr ? memReg_10_core_instruction : _GEN_455; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_457 = 4'hb == readPtr ? memReg_11_core_instruction : _GEN_456; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_458 = 4'hc == readPtr ? memReg_12_core_instruction : _GEN_457; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_459 = 4'hd == readPtr ? memReg_13_core_instruction : _GEN_458; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_460 = 4'he == readPtr ? memReg_14_core_instruction : _GEN_459; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_463 = 4'h1 == readPtr ? memReg_1_core_robAddr : memReg_0_core_robAddr; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_464 = 4'h2 == readPtr ? memReg_2_core_robAddr : _GEN_463; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_465 = 4'h3 == readPtr ? memReg_3_core_robAddr : _GEN_464; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_466 = 4'h4 == readPtr ? memReg_4_core_robAddr : _GEN_465; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_467 = 4'h5 == readPtr ? memReg_5_core_robAddr : _GEN_466; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_468 = 4'h6 == readPtr ? memReg_6_core_robAddr : _GEN_467; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_469 = 4'h7 == readPtr ? memReg_7_core_robAddr : _GEN_468; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_470 = 4'h8 == readPtr ? memReg_8_core_robAddr : _GEN_469; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_471 = 4'h9 == readPtr ? memReg_9_core_robAddr : _GEN_470; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_472 = 4'ha == readPtr ? memReg_10_core_robAddr : _GEN_471; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_473 = 4'hb == readPtr ? memReg_11_core_robAddr : _GEN_472; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_474 = 4'hc == readPtr ? memReg_12_core_robAddr : _GEN_473; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_475 = 4'hd == readPtr ? memReg_13_core_robAddr : _GEN_474; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_476 = 4'he == readPtr ? memReg_14_core_robAddr : _GEN_475; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_479 = 4'h1 == readPtr ? memReg_1_core_prfDest : memReg_0_core_prfDest; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_480 = 4'h2 == readPtr ? memReg_2_core_prfDest : _GEN_479; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_481 = 4'h3 == readPtr ? memReg_3_core_prfDest : _GEN_480; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_482 = 4'h4 == readPtr ? memReg_4_core_prfDest : _GEN_481; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_483 = 4'h5 == readPtr ? memReg_5_core_prfDest : _GEN_482; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_484 = 4'h6 == readPtr ? memReg_6_core_prfDest : _GEN_483; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_485 = 4'h7 == readPtr ? memReg_7_core_prfDest : _GEN_484; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_486 = 4'h8 == readPtr ? memReg_8_core_prfDest : _GEN_485; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_487 = 4'h9 == readPtr ? memReg_9_core_prfDest : _GEN_486; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_488 = 4'ha == readPtr ? memReg_10_core_prfDest : _GEN_487; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_489 = 4'hb == readPtr ? memReg_11_core_prfDest : _GEN_488; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_490 = 4'hc == readPtr ? memReg_12_core_prfDest : _GEN_489; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_491 = 4'hd == readPtr ? memReg_13_core_prfDest : _GEN_490; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_492 = 4'he == readPtr ? memReg_14_core_prfDest : _GEN_491; // @[fifo.scala 86:{13,13}]
  wire  _GEN_495 = 4'h1 == readPtr ? memReg_1_branch_valid : memReg_0_branch_valid; // @[fifo.scala 86:{13,13}]
  wire  _GEN_496 = 4'h2 == readPtr ? memReg_2_branch_valid : _GEN_495; // @[fifo.scala 86:{13,13}]
  wire  _GEN_497 = 4'h3 == readPtr ? memReg_3_branch_valid : _GEN_496; // @[fifo.scala 86:{13,13}]
  wire  _GEN_498 = 4'h4 == readPtr ? memReg_4_branch_valid : _GEN_497; // @[fifo.scala 86:{13,13}]
  wire  _GEN_499 = 4'h5 == readPtr ? memReg_5_branch_valid : _GEN_498; // @[fifo.scala 86:{13,13}]
  wire  _GEN_500 = 4'h6 == readPtr ? memReg_6_branch_valid : _GEN_499; // @[fifo.scala 86:{13,13}]
  wire  _GEN_501 = 4'h7 == readPtr ? memReg_7_branch_valid : _GEN_500; // @[fifo.scala 86:{13,13}]
  wire  _GEN_502 = 4'h8 == readPtr ? memReg_8_branch_valid : _GEN_501; // @[fifo.scala 86:{13,13}]
  wire  _GEN_503 = 4'h9 == readPtr ? memReg_9_branch_valid : _GEN_502; // @[fifo.scala 86:{13,13}]
  wire  _GEN_504 = 4'ha == readPtr ? memReg_10_branch_valid : _GEN_503; // @[fifo.scala 86:{13,13}]
  wire  _GEN_505 = 4'hb == readPtr ? memReg_11_branch_valid : _GEN_504; // @[fifo.scala 86:{13,13}]
  wire  _GEN_506 = 4'hc == readPtr ? memReg_12_branch_valid : _GEN_505; // @[fifo.scala 86:{13,13}]
  wire  _GEN_507 = 4'hd == readPtr ? memReg_13_branch_valid : _GEN_506; // @[fifo.scala 86:{13,13}]
  wire  _GEN_508 = 4'he == readPtr ? memReg_14_branch_valid : _GEN_507; // @[fifo.scala 86:{13,13}]
  wire  _GEN_509 = 4'hf == readPtr ? memReg_15_branch_valid : _GEN_508; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_511 = 4'h1 == readPtr ? memReg_1_branch_mask : memReg_0_branch_mask; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_512 = 4'h2 == readPtr ? memReg_2_branch_mask : _GEN_511; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_513 = 4'h3 == readPtr ? memReg_3_branch_mask : _GEN_512; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_514 = 4'h4 == readPtr ? memReg_4_branch_mask : _GEN_513; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_515 = 4'h5 == readPtr ? memReg_5_branch_mask : _GEN_514; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_516 = 4'h6 == readPtr ? memReg_6_branch_mask : _GEN_515; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_517 = 4'h7 == readPtr ? memReg_7_branch_mask : _GEN_516; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_518 = 4'h8 == readPtr ? memReg_8_branch_mask : _GEN_517; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_519 = 4'h9 == readPtr ? memReg_9_branch_mask : _GEN_518; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_520 = 4'ha == readPtr ? memReg_10_branch_mask : _GEN_519; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_521 = 4'hb == readPtr ? memReg_11_branch_mask : _GEN_520; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_522 = 4'hc == readPtr ? memReg_12_branch_mask : _GEN_521; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_523 = 4'hd == readPtr ? memReg_13_branch_mask : _GEN_522; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_524 = 4'he == readPtr ? memReg_14_branch_mask : _GEN_523; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_525 = 4'hf == readPtr ? memReg_15_branch_mask : _GEN_524; // @[fifo.scala 86:{13,13}]
  wire  _GEN_527 = 4'h1 == readPtr ? memReg_1_writeData_valid : memReg_0_writeData_valid; // @[fifo.scala 86:{13,13}]
  wire  _GEN_528 = 4'h2 == readPtr ? memReg_2_writeData_valid : _GEN_527; // @[fifo.scala 86:{13,13}]
  wire  _GEN_529 = 4'h3 == readPtr ? memReg_3_writeData_valid : _GEN_528; // @[fifo.scala 86:{13,13}]
  wire  _GEN_530 = 4'h4 == readPtr ? memReg_4_writeData_valid : _GEN_529; // @[fifo.scala 86:{13,13}]
  wire  _GEN_531 = 4'h5 == readPtr ? memReg_5_writeData_valid : _GEN_530; // @[fifo.scala 86:{13,13}]
  wire  _GEN_532 = 4'h6 == readPtr ? memReg_6_writeData_valid : _GEN_531; // @[fifo.scala 86:{13,13}]
  wire  _GEN_533 = 4'h7 == readPtr ? memReg_7_writeData_valid : _GEN_532; // @[fifo.scala 86:{13,13}]
  wire  _GEN_534 = 4'h8 == readPtr ? memReg_8_writeData_valid : _GEN_533; // @[fifo.scala 86:{13,13}]
  wire  _GEN_535 = 4'h9 == readPtr ? memReg_9_writeData_valid : _GEN_534; // @[fifo.scala 86:{13,13}]
  wire  _GEN_536 = 4'ha == readPtr ? memReg_10_writeData_valid : _GEN_535; // @[fifo.scala 86:{13,13}]
  wire  _GEN_537 = 4'hb == readPtr ? memReg_11_writeData_valid : _GEN_536; // @[fifo.scala 86:{13,13}]
  wire  _GEN_538 = 4'hc == readPtr ? memReg_12_writeData_valid : _GEN_537; // @[fifo.scala 86:{13,13}]
  wire  _GEN_539 = 4'hd == readPtr ? memReg_13_writeData_valid : _GEN_538; // @[fifo.scala 86:{13,13}]
  wire  _GEN_540 = 4'he == readPtr ? memReg_14_writeData_valid : _GEN_539; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_543 = 4'h1 == readPtr ? memReg_1_writeData_data : memReg_0_writeData_data; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_544 = 4'h2 == readPtr ? memReg_2_writeData_data : _GEN_543; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_545 = 4'h3 == readPtr ? memReg_3_writeData_data : _GEN_544; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_546 = 4'h4 == readPtr ? memReg_4_writeData_data : _GEN_545; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_547 = 4'h5 == readPtr ? memReg_5_writeData_data : _GEN_546; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_548 = 4'h6 == readPtr ? memReg_6_writeData_data : _GEN_547; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_549 = 4'h7 == readPtr ? memReg_7_writeData_data : _GEN_548; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_550 = 4'h8 == readPtr ? memReg_8_writeData_data : _GEN_549; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_551 = 4'h9 == readPtr ? memReg_9_writeData_data : _GEN_550; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_552 = 4'ha == readPtr ? memReg_10_writeData_data : _GEN_551; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_553 = 4'hb == readPtr ? memReg_11_writeData_data : _GEN_552; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_554 = 4'hc == readPtr ? memReg_12_writeData_data : _GEN_553; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_555 = 4'hd == readPtr ? memReg_13_writeData_data : _GEN_554; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_556 = 4'he == readPtr ? memReg_14_writeData_data : _GEN_555; // @[fifo.scala 86:{13,13}]
  wire [1:0] _GEN_575 = 4'h1 == readPtr ? memReg_1_cacheLine_response : memReg_0_cacheLine_response; // @[fifo.scala 86:{13,13}]
  wire [1:0] _GEN_576 = 4'h2 == readPtr ? memReg_2_cacheLine_response : _GEN_575; // @[fifo.scala 86:{13,13}]
  wire [1:0] _GEN_577 = 4'h3 == readPtr ? memReg_3_cacheLine_response : _GEN_576; // @[fifo.scala 86:{13,13}]
  wire [1:0] _GEN_578 = 4'h4 == readPtr ? memReg_4_cacheLine_response : _GEN_577; // @[fifo.scala 86:{13,13}]
  wire [1:0] _GEN_579 = 4'h5 == readPtr ? memReg_5_cacheLine_response : _GEN_578; // @[fifo.scala 86:{13,13}]
  wire [1:0] _GEN_580 = 4'h6 == readPtr ? memReg_6_cacheLine_response : _GEN_579; // @[fifo.scala 86:{13,13}]
  wire [1:0] _GEN_581 = 4'h7 == readPtr ? memReg_7_cacheLine_response : _GEN_580; // @[fifo.scala 86:{13,13}]
  wire [1:0] _GEN_582 = 4'h8 == readPtr ? memReg_8_cacheLine_response : _GEN_581; // @[fifo.scala 86:{13,13}]
  wire [1:0] _GEN_583 = 4'h9 == readPtr ? memReg_9_cacheLine_response : _GEN_582; // @[fifo.scala 86:{13,13}]
  wire [1:0] _GEN_584 = 4'ha == readPtr ? memReg_10_cacheLine_response : _GEN_583; // @[fifo.scala 86:{13,13}]
  wire [1:0] _GEN_585 = 4'hb == readPtr ? memReg_11_cacheLine_response : _GEN_584; // @[fifo.scala 86:{13,13}]
  wire [1:0] _GEN_586 = 4'hc == readPtr ? memReg_12_cacheLine_response : _GEN_585; // @[fifo.scala 86:{13,13}]
  wire [1:0] _GEN_587 = 4'hd == readPtr ? memReg_13_cacheLine_response : _GEN_586; // @[fifo.scala 86:{13,13}]
  wire [1:0] _GEN_588 = 4'he == readPtr ? memReg_14_cacheLine_response : _GEN_587; // @[fifo.scala 86:{13,13}]
  wire [4:0] _T_8 = write_data_branch_mask & branchOps_branchMask; // @[utils.scala 62:31]
  wire  _T_9 = |_T_8; // @[utils.scala 62:55]
  wire [4:0] _memReg_branch_mask_T = write_data_branch_mask ^ branchOps_branchMask; // @[utils.scala 63:42]
  wire [4:0] _GEN_606 = 4'h0 == writePtr ? _memReg_branch_mask_T : _GEN_318; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_607 = 4'h1 == writePtr ? _memReg_branch_mask_T : _GEN_319; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_608 = 4'h2 == writePtr ? _memReg_branch_mask_T : _GEN_320; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_609 = 4'h3 == writePtr ? _memReg_branch_mask_T : _GEN_321; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_610 = 4'h4 == writePtr ? _memReg_branch_mask_T : _GEN_322; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_611 = 4'h5 == writePtr ? _memReg_branch_mask_T : _GEN_323; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_612 = 4'h6 == writePtr ? _memReg_branch_mask_T : _GEN_324; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_613 = 4'h7 == writePtr ? _memReg_branch_mask_T : _GEN_325; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_614 = 4'h8 == writePtr ? _memReg_branch_mask_T : _GEN_326; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_615 = 4'h9 == writePtr ? _memReg_branch_mask_T : _GEN_327; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_616 = 4'ha == writePtr ? _memReg_branch_mask_T : _GEN_328; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_617 = 4'hb == writePtr ? _memReg_branch_mask_T : _GEN_329; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_618 = 4'hc == writePtr ? _memReg_branch_mask_T : _GEN_330; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_619 = 4'hd == writePtr ? _memReg_branch_mask_T : _GEN_331; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_620 = 4'he == writePtr ? _memReg_branch_mask_T : _GEN_332; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_621 = 4'hf == writePtr ? _memReg_branch_mask_T : _GEN_333; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_622 = 4'h0 == writePtr ? write_data_branch_mask : _GEN_318; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_623 = 4'h1 == writePtr ? write_data_branch_mask : _GEN_319; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_624 = 4'h2 == writePtr ? write_data_branch_mask : _GEN_320; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_625 = 4'h3 == writePtr ? write_data_branch_mask : _GEN_321; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_626 = 4'h4 == writePtr ? write_data_branch_mask : _GEN_322; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_627 = 4'h5 == writePtr ? write_data_branch_mask : _GEN_323; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_628 = 4'h6 == writePtr ? write_data_branch_mask : _GEN_324; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_629 = 4'h7 == writePtr ? write_data_branch_mask : _GEN_325; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_630 = 4'h8 == writePtr ? write_data_branch_mask : _GEN_326; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_631 = 4'h9 == writePtr ? write_data_branch_mask : _GEN_327; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_632 = 4'ha == writePtr ? write_data_branch_mask : _GEN_328; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_633 = 4'hb == writePtr ? write_data_branch_mask : _GEN_329; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_634 = 4'hc == writePtr ? write_data_branch_mask : _GEN_330; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_635 = 4'hd == writePtr ? write_data_branch_mask : _GEN_331; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_636 = 4'he == writePtr ? write_data_branch_mask : _GEN_332; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_637 = 4'hf == writePtr ? write_data_branch_mask : _GEN_333; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_638 = |_T_8 ? _GEN_606 : _GEN_622; // @[utils.scala 62:60]
  wire [4:0] _GEN_639 = |_T_8 ? _GEN_607 : _GEN_623; // @[utils.scala 62:60]
  wire [4:0] _GEN_640 = |_T_8 ? _GEN_608 : _GEN_624; // @[utils.scala 62:60]
  wire [4:0] _GEN_641 = |_T_8 ? _GEN_609 : _GEN_625; // @[utils.scala 62:60]
  wire [4:0] _GEN_642 = |_T_8 ? _GEN_610 : _GEN_626; // @[utils.scala 62:60]
  wire [4:0] _GEN_643 = |_T_8 ? _GEN_611 : _GEN_627; // @[utils.scala 62:60]
  wire [4:0] _GEN_644 = |_T_8 ? _GEN_612 : _GEN_628; // @[utils.scala 62:60]
  wire [4:0] _GEN_645 = |_T_8 ? _GEN_613 : _GEN_629; // @[utils.scala 62:60]
  wire [4:0] _GEN_646 = |_T_8 ? _GEN_614 : _GEN_630; // @[utils.scala 62:60]
  wire [4:0] _GEN_647 = |_T_8 ? _GEN_615 : _GEN_631; // @[utils.scala 62:60]
  wire [4:0] _GEN_648 = |_T_8 ? _GEN_616 : _GEN_632; // @[utils.scala 62:60]
  wire [4:0] _GEN_649 = |_T_8 ? _GEN_617 : _GEN_633; // @[utils.scala 62:60]
  wire [4:0] _GEN_650 = |_T_8 ? _GEN_618 : _GEN_634; // @[utils.scala 62:60]
  wire [4:0] _GEN_651 = |_T_8 ? _GEN_619 : _GEN_635; // @[utils.scala 62:60]
  wire [4:0] _GEN_652 = |_T_8 ? _GEN_620 : _GEN_636; // @[utils.scala 62:60]
  wire [4:0] _GEN_653 = |_T_8 ? _GEN_621 : _GEN_637; // @[utils.scala 62:60]
  wire  _GEN_654 = 4'h0 == writePtr ? write_data_branch_valid : _GEN_302; // @[utils.scala 67:{22,22}]
  wire  _GEN_655 = 4'h1 == writePtr ? write_data_branch_valid : _GEN_303; // @[utils.scala 67:{22,22}]
  wire  _GEN_656 = 4'h2 == writePtr ? write_data_branch_valid : _GEN_304; // @[utils.scala 67:{22,22}]
  wire  _GEN_657 = 4'h3 == writePtr ? write_data_branch_valid : _GEN_305; // @[utils.scala 67:{22,22}]
  wire  _GEN_658 = 4'h4 == writePtr ? write_data_branch_valid : _GEN_306; // @[utils.scala 67:{22,22}]
  wire  _GEN_659 = 4'h5 == writePtr ? write_data_branch_valid : _GEN_307; // @[utils.scala 67:{22,22}]
  wire  _GEN_660 = 4'h6 == writePtr ? write_data_branch_valid : _GEN_308; // @[utils.scala 67:{22,22}]
  wire  _GEN_661 = 4'h7 == writePtr ? write_data_branch_valid : _GEN_309; // @[utils.scala 67:{22,22}]
  wire  _GEN_662 = 4'h8 == writePtr ? write_data_branch_valid : _GEN_310; // @[utils.scala 67:{22,22}]
  wire  _GEN_663 = 4'h9 == writePtr ? write_data_branch_valid : _GEN_311; // @[utils.scala 67:{22,22}]
  wire  _GEN_664 = 4'ha == writePtr ? write_data_branch_valid : _GEN_312; // @[utils.scala 67:{22,22}]
  wire  _GEN_665 = 4'hb == writePtr ? write_data_branch_valid : _GEN_313; // @[utils.scala 67:{22,22}]
  wire  _GEN_666 = 4'hc == writePtr ? write_data_branch_valid : _GEN_314; // @[utils.scala 67:{22,22}]
  wire  _GEN_667 = 4'hd == writePtr ? write_data_branch_valid : _GEN_315; // @[utils.scala 67:{22,22}]
  wire  _GEN_668 = 4'he == writePtr ? write_data_branch_valid : _GEN_316; // @[utils.scala 67:{22,22}]
  wire  _GEN_669 = 4'hf == writePtr ? write_data_branch_valid : _GEN_317; // @[utils.scala 67:{22,22}]
  wire  _GEN_670 = 4'h0 == writePtr ? 1'h0 : _GEN_302; // @[utils.scala 71:{24,24}]
  wire  _GEN_671 = 4'h1 == writePtr ? 1'h0 : _GEN_303; // @[utils.scala 71:{24,24}]
  wire  _GEN_672 = 4'h2 == writePtr ? 1'h0 : _GEN_304; // @[utils.scala 71:{24,24}]
  wire  _GEN_673 = 4'h3 == writePtr ? 1'h0 : _GEN_305; // @[utils.scala 71:{24,24}]
  wire  _GEN_674 = 4'h4 == writePtr ? 1'h0 : _GEN_306; // @[utils.scala 71:{24,24}]
  wire  _GEN_675 = 4'h5 == writePtr ? 1'h0 : _GEN_307; // @[utils.scala 71:{24,24}]
  wire  _GEN_676 = 4'h6 == writePtr ? 1'h0 : _GEN_308; // @[utils.scala 71:{24,24}]
  wire  _GEN_677 = 4'h7 == writePtr ? 1'h0 : _GEN_309; // @[utils.scala 71:{24,24}]
  wire  _GEN_678 = 4'h8 == writePtr ? 1'h0 : _GEN_310; // @[utils.scala 71:{24,24}]
  wire  _GEN_679 = 4'h9 == writePtr ? 1'h0 : _GEN_311; // @[utils.scala 71:{24,24}]
  wire  _GEN_680 = 4'ha == writePtr ? 1'h0 : _GEN_312; // @[utils.scala 71:{24,24}]
  wire  _GEN_681 = 4'hb == writePtr ? 1'h0 : _GEN_313; // @[utils.scala 71:{24,24}]
  wire  _GEN_682 = 4'hc == writePtr ? 1'h0 : _GEN_314; // @[utils.scala 71:{24,24}]
  wire  _GEN_683 = 4'hd == writePtr ? 1'h0 : _GEN_315; // @[utils.scala 71:{24,24}]
  wire  _GEN_684 = 4'he == writePtr ? 1'h0 : _GEN_316; // @[utils.scala 71:{24,24}]
  wire  _GEN_685 = 4'hf == writePtr ? 1'h0 : _GEN_317; // @[utils.scala 71:{24,24}]
  wire [4:0] _GEN_686 = 4'h0 == writePtr ? 5'h0 : _GEN_318; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_687 = 4'h1 == writePtr ? 5'h0 : _GEN_319; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_688 = 4'h2 == writePtr ? 5'h0 : _GEN_320; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_689 = 4'h3 == writePtr ? 5'h0 : _GEN_321; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_690 = 4'h4 == writePtr ? 5'h0 : _GEN_322; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_691 = 4'h5 == writePtr ? 5'h0 : _GEN_323; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_692 = 4'h6 == writePtr ? 5'h0 : _GEN_324; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_693 = 4'h7 == writePtr ? 5'h0 : _GEN_325; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_694 = 4'h8 == writePtr ? 5'h0 : _GEN_326; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_695 = 4'h9 == writePtr ? 5'h0 : _GEN_327; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_696 = 4'ha == writePtr ? 5'h0 : _GEN_328; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_697 = 4'hb == writePtr ? 5'h0 : _GEN_329; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_698 = 4'hc == writePtr ? 5'h0 : _GEN_330; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_699 = 4'hd == writePtr ? 5'h0 : _GEN_331; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_700 = 4'he == writePtr ? 5'h0 : _GEN_332; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_701 = 4'hf == writePtr ? 5'h0 : _GEN_333; // @[utils.scala 72:{23,23}]
  wire  _GEN_734 = _T_9 ? _GEN_670 : _GEN_654; // @[utils.scala 70:60]
  wire  _GEN_735 = _T_9 ? _GEN_671 : _GEN_655; // @[utils.scala 70:60]
  wire  _GEN_736 = _T_9 ? _GEN_672 : _GEN_656; // @[utils.scala 70:60]
  wire  _GEN_737 = _T_9 ? _GEN_673 : _GEN_657; // @[utils.scala 70:60]
  wire  _GEN_738 = _T_9 ? _GEN_674 : _GEN_658; // @[utils.scala 70:60]
  wire  _GEN_739 = _T_9 ? _GEN_675 : _GEN_659; // @[utils.scala 70:60]
  wire  _GEN_740 = _T_9 ? _GEN_676 : _GEN_660; // @[utils.scala 70:60]
  wire  _GEN_741 = _T_9 ? _GEN_677 : _GEN_661; // @[utils.scala 70:60]
  wire  _GEN_742 = _T_9 ? _GEN_678 : _GEN_662; // @[utils.scala 70:60]
  wire  _GEN_743 = _T_9 ? _GEN_679 : _GEN_663; // @[utils.scala 70:60]
  wire  _GEN_744 = _T_9 ? _GEN_680 : _GEN_664; // @[utils.scala 70:60]
  wire  _GEN_745 = _T_9 ? _GEN_681 : _GEN_665; // @[utils.scala 70:60]
  wire  _GEN_746 = _T_9 ? _GEN_682 : _GEN_666; // @[utils.scala 70:60]
  wire  _GEN_747 = _T_9 ? _GEN_683 : _GEN_667; // @[utils.scala 70:60]
  wire  _GEN_748 = _T_9 ? _GEN_684 : _GEN_668; // @[utils.scala 70:60]
  wire  _GEN_749 = _T_9 ? _GEN_685 : _GEN_669; // @[utils.scala 70:60]
  wire [4:0] _GEN_750 = _T_9 ? _GEN_686 : _GEN_622; // @[utils.scala 70:60]
  wire [4:0] _GEN_751 = _T_9 ? _GEN_687 : _GEN_623; // @[utils.scala 70:60]
  wire [4:0] _GEN_752 = _T_9 ? _GEN_688 : _GEN_624; // @[utils.scala 70:60]
  wire [4:0] _GEN_753 = _T_9 ? _GEN_689 : _GEN_625; // @[utils.scala 70:60]
  wire [4:0] _GEN_754 = _T_9 ? _GEN_690 : _GEN_626; // @[utils.scala 70:60]
  wire [4:0] _GEN_755 = _T_9 ? _GEN_691 : _GEN_627; // @[utils.scala 70:60]
  wire [4:0] _GEN_756 = _T_9 ? _GEN_692 : _GEN_628; // @[utils.scala 70:60]
  wire [4:0] _GEN_757 = _T_9 ? _GEN_693 : _GEN_629; // @[utils.scala 70:60]
  wire [4:0] _GEN_758 = _T_9 ? _GEN_694 : _GEN_630; // @[utils.scala 70:60]
  wire [4:0] _GEN_759 = _T_9 ? _GEN_695 : _GEN_631; // @[utils.scala 70:60]
  wire [4:0] _GEN_760 = _T_9 ? _GEN_696 : _GEN_632; // @[utils.scala 70:60]
  wire [4:0] _GEN_761 = _T_9 ? _GEN_697 : _GEN_633; // @[utils.scala 70:60]
  wire [4:0] _GEN_762 = _T_9 ? _GEN_698 : _GEN_634; // @[utils.scala 70:60]
  wire [4:0] _GEN_763 = _T_9 ? _GEN_699 : _GEN_635; // @[utils.scala 70:60]
  wire [4:0] _GEN_764 = _T_9 ? _GEN_700 : _GEN_636; // @[utils.scala 70:60]
  wire [4:0] _GEN_765 = _T_9 ? _GEN_701 : _GEN_637; // @[utils.scala 70:60]
  wire [4:0] _GEN_766 = branchOps_passed ? _GEN_638 : _GEN_750; // @[utils.scala 60:30]
  wire [4:0] _GEN_767 = branchOps_passed ? _GEN_639 : _GEN_751; // @[utils.scala 60:30]
  wire [4:0] _GEN_768 = branchOps_passed ? _GEN_640 : _GEN_752; // @[utils.scala 60:30]
  wire [4:0] _GEN_769 = branchOps_passed ? _GEN_641 : _GEN_753; // @[utils.scala 60:30]
  wire [4:0] _GEN_770 = branchOps_passed ? _GEN_642 : _GEN_754; // @[utils.scala 60:30]
  wire [4:0] _GEN_771 = branchOps_passed ? _GEN_643 : _GEN_755; // @[utils.scala 60:30]
  wire [4:0] _GEN_772 = branchOps_passed ? _GEN_644 : _GEN_756; // @[utils.scala 60:30]
  wire [4:0] _GEN_773 = branchOps_passed ? _GEN_645 : _GEN_757; // @[utils.scala 60:30]
  wire [4:0] _GEN_774 = branchOps_passed ? _GEN_646 : _GEN_758; // @[utils.scala 60:30]
  wire [4:0] _GEN_775 = branchOps_passed ? _GEN_647 : _GEN_759; // @[utils.scala 60:30]
  wire [4:0] _GEN_776 = branchOps_passed ? _GEN_648 : _GEN_760; // @[utils.scala 60:30]
  wire [4:0] _GEN_777 = branchOps_passed ? _GEN_649 : _GEN_761; // @[utils.scala 60:30]
  wire [4:0] _GEN_778 = branchOps_passed ? _GEN_650 : _GEN_762; // @[utils.scala 60:30]
  wire [4:0] _GEN_779 = branchOps_passed ? _GEN_651 : _GEN_763; // @[utils.scala 60:30]
  wire [4:0] _GEN_780 = branchOps_passed ? _GEN_652 : _GEN_764; // @[utils.scala 60:30]
  wire [4:0] _GEN_781 = branchOps_passed ? _GEN_653 : _GEN_765; // @[utils.scala 60:30]
  wire  _GEN_782 = branchOps_passed ? _GEN_654 : _GEN_734; // @[utils.scala 60:30]
  wire  _GEN_783 = branchOps_passed ? _GEN_655 : _GEN_735; // @[utils.scala 60:30]
  wire  _GEN_784 = branchOps_passed ? _GEN_656 : _GEN_736; // @[utils.scala 60:30]
  wire  _GEN_785 = branchOps_passed ? _GEN_657 : _GEN_737; // @[utils.scala 60:30]
  wire  _GEN_786 = branchOps_passed ? _GEN_658 : _GEN_738; // @[utils.scala 60:30]
  wire  _GEN_787 = branchOps_passed ? _GEN_659 : _GEN_739; // @[utils.scala 60:30]
  wire  _GEN_788 = branchOps_passed ? _GEN_660 : _GEN_740; // @[utils.scala 60:30]
  wire  _GEN_789 = branchOps_passed ? _GEN_661 : _GEN_741; // @[utils.scala 60:30]
  wire  _GEN_790 = branchOps_passed ? _GEN_662 : _GEN_742; // @[utils.scala 60:30]
  wire  _GEN_791 = branchOps_passed ? _GEN_663 : _GEN_743; // @[utils.scala 60:30]
  wire  _GEN_792 = branchOps_passed ? _GEN_664 : _GEN_744; // @[utils.scala 60:30]
  wire  _GEN_793 = branchOps_passed ? _GEN_665 : _GEN_745; // @[utils.scala 60:30]
  wire  _GEN_794 = branchOps_passed ? _GEN_666 : _GEN_746; // @[utils.scala 60:30]
  wire  _GEN_795 = branchOps_passed ? _GEN_667 : _GEN_747; // @[utils.scala 60:30]
  wire  _GEN_796 = branchOps_passed ? _GEN_668 : _GEN_748; // @[utils.scala 60:30]
  wire  _GEN_797 = branchOps_passed ? _GEN_669 : _GEN_749; // @[utils.scala 60:30]
  wire [4:0] _GEN_830 = branchOps_valid ? _GEN_766 : _GEN_622; // @[utils.scala 59:26]
  wire [4:0] _GEN_831 = branchOps_valid ? _GEN_767 : _GEN_623; // @[utils.scala 59:26]
  wire [4:0] _GEN_832 = branchOps_valid ? _GEN_768 : _GEN_624; // @[utils.scala 59:26]
  wire [4:0] _GEN_833 = branchOps_valid ? _GEN_769 : _GEN_625; // @[utils.scala 59:26]
  wire [4:0] _GEN_834 = branchOps_valid ? _GEN_770 : _GEN_626; // @[utils.scala 59:26]
  wire [4:0] _GEN_835 = branchOps_valid ? _GEN_771 : _GEN_627; // @[utils.scala 59:26]
  wire [4:0] _GEN_836 = branchOps_valid ? _GEN_772 : _GEN_628; // @[utils.scala 59:26]
  wire [4:0] _GEN_837 = branchOps_valid ? _GEN_773 : _GEN_629; // @[utils.scala 59:26]
  wire [4:0] _GEN_838 = branchOps_valid ? _GEN_774 : _GEN_630; // @[utils.scala 59:26]
  wire [4:0] _GEN_839 = branchOps_valid ? _GEN_775 : _GEN_631; // @[utils.scala 59:26]
  wire [4:0] _GEN_840 = branchOps_valid ? _GEN_776 : _GEN_632; // @[utils.scala 59:26]
  wire [4:0] _GEN_841 = branchOps_valid ? _GEN_777 : _GEN_633; // @[utils.scala 59:26]
  wire [4:0] _GEN_842 = branchOps_valid ? _GEN_778 : _GEN_634; // @[utils.scala 59:26]
  wire [4:0] _GEN_843 = branchOps_valid ? _GEN_779 : _GEN_635; // @[utils.scala 59:26]
  wire [4:0] _GEN_844 = branchOps_valid ? _GEN_780 : _GEN_636; // @[utils.scala 59:26]
  wire [4:0] _GEN_845 = branchOps_valid ? _GEN_781 : _GEN_637; // @[utils.scala 59:26]
  wire  _GEN_846 = branchOps_valid ? _GEN_782 : _GEN_654; // @[utils.scala 59:26]
  wire  _GEN_847 = branchOps_valid ? _GEN_783 : _GEN_655; // @[utils.scala 59:26]
  wire  _GEN_848 = branchOps_valid ? _GEN_784 : _GEN_656; // @[utils.scala 59:26]
  wire  _GEN_849 = branchOps_valid ? _GEN_785 : _GEN_657; // @[utils.scala 59:26]
  wire  _GEN_850 = branchOps_valid ? _GEN_786 : _GEN_658; // @[utils.scala 59:26]
  wire  _GEN_851 = branchOps_valid ? _GEN_787 : _GEN_659; // @[utils.scala 59:26]
  wire  _GEN_852 = branchOps_valid ? _GEN_788 : _GEN_660; // @[utils.scala 59:26]
  wire  _GEN_853 = branchOps_valid ? _GEN_789 : _GEN_661; // @[utils.scala 59:26]
  wire  _GEN_854 = branchOps_valid ? _GEN_790 : _GEN_662; // @[utils.scala 59:26]
  wire  _GEN_855 = branchOps_valid ? _GEN_791 : _GEN_663; // @[utils.scala 59:26]
  wire  _GEN_856 = branchOps_valid ? _GEN_792 : _GEN_664; // @[utils.scala 59:26]
  wire  _GEN_857 = branchOps_valid ? _GEN_793 : _GEN_665; // @[utils.scala 59:26]
  wire  _GEN_858 = branchOps_valid ? _GEN_794 : _GEN_666; // @[utils.scala 59:26]
  wire  _GEN_859 = branchOps_valid ? _GEN_795 : _GEN_667; // @[utils.scala 59:26]
  wire  _GEN_860 = branchOps_valid ? _GEN_796 : _GEN_668; // @[utils.scala 59:26]
  wire  _GEN_861 = branchOps_valid ? _GEN_797 : _GEN_669; // @[utils.scala 59:26]
  wire [4:0] _GEN_862 = incrWrite ? _GEN_830 : _GEN_318; // @[fifo.scala 97:16]
  wire [4:0] _GEN_863 = incrWrite ? _GEN_831 : _GEN_319; // @[fifo.scala 97:16]
  wire [4:0] _GEN_864 = incrWrite ? _GEN_832 : _GEN_320; // @[fifo.scala 97:16]
  wire [4:0] _GEN_865 = incrWrite ? _GEN_833 : _GEN_321; // @[fifo.scala 97:16]
  wire [4:0] _GEN_866 = incrWrite ? _GEN_834 : _GEN_322; // @[fifo.scala 97:16]
  wire [4:0] _GEN_867 = incrWrite ? _GEN_835 : _GEN_323; // @[fifo.scala 97:16]
  wire [4:0] _GEN_868 = incrWrite ? _GEN_836 : _GEN_324; // @[fifo.scala 97:16]
  wire [4:0] _GEN_869 = incrWrite ? _GEN_837 : _GEN_325; // @[fifo.scala 97:16]
  wire [4:0] _GEN_870 = incrWrite ? _GEN_838 : _GEN_326; // @[fifo.scala 97:16]
  wire [4:0] _GEN_871 = incrWrite ? _GEN_839 : _GEN_327; // @[fifo.scala 97:16]
  wire [4:0] _GEN_872 = incrWrite ? _GEN_840 : _GEN_328; // @[fifo.scala 97:16]
  wire [4:0] _GEN_873 = incrWrite ? _GEN_841 : _GEN_329; // @[fifo.scala 97:16]
  wire [4:0] _GEN_874 = incrWrite ? _GEN_842 : _GEN_330; // @[fifo.scala 97:16]
  wire [4:0] _GEN_875 = incrWrite ? _GEN_843 : _GEN_331; // @[fifo.scala 97:16]
  wire [4:0] _GEN_876 = incrWrite ? _GEN_844 : _GEN_332; // @[fifo.scala 97:16]
  wire [4:0] _GEN_877 = incrWrite ? _GEN_845 : _GEN_333; // @[fifo.scala 97:16]
  wire  _GEN_878 = incrWrite ? _GEN_846 : _GEN_302; // @[fifo.scala 97:16]
  wire  _GEN_879 = incrWrite ? _GEN_847 : _GEN_303; // @[fifo.scala 97:16]
  wire  _GEN_880 = incrWrite ? _GEN_848 : _GEN_304; // @[fifo.scala 97:16]
  wire  _GEN_881 = incrWrite ? _GEN_849 : _GEN_305; // @[fifo.scala 97:16]
  wire  _GEN_882 = incrWrite ? _GEN_850 : _GEN_306; // @[fifo.scala 97:16]
  wire  _GEN_883 = incrWrite ? _GEN_851 : _GEN_307; // @[fifo.scala 97:16]
  wire  _GEN_884 = incrWrite ? _GEN_852 : _GEN_308; // @[fifo.scala 97:16]
  wire  _GEN_885 = incrWrite ? _GEN_853 : _GEN_309; // @[fifo.scala 97:16]
  wire  _GEN_886 = incrWrite ? _GEN_854 : _GEN_310; // @[fifo.scala 97:16]
  wire  _GEN_887 = incrWrite ? _GEN_855 : _GEN_311; // @[fifo.scala 97:16]
  wire  _GEN_888 = incrWrite ? _GEN_856 : _GEN_312; // @[fifo.scala 97:16]
  wire  _GEN_889 = incrWrite ? _GEN_857 : _GEN_313; // @[fifo.scala 97:16]
  wire  _GEN_890 = incrWrite ? _GEN_858 : _GEN_314; // @[fifo.scala 97:16]
  wire  _GEN_891 = incrWrite ? _GEN_859 : _GEN_315; // @[fifo.scala 97:16]
  wire  _GEN_892 = incrWrite ? _GEN_860 : _GEN_316; // @[fifo.scala 97:16]
  wire  _GEN_893 = incrWrite ? _GEN_861 : _GEN_317; // @[fifo.scala 97:16]
  wire [3:0] startPointer = read_ready ? _nextVal_T_2 : readPtr; // @[fifo.scala 102:25]
  wire [3:0] endPointer = writePtr - 4'h1; // @[fifo.scala 103:29]
  wire [4:0] _T_15 = memReg_0_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_16 = |_T_15; // @[fifo.scala 109:63]
  wire [4:0] _memReg_0_branch_mask_T = memReg_0_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _T_22 = memReg_1_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_23 = |_T_22; // @[fifo.scala 109:63]
  wire [4:0] _memReg_1_branch_mask_T = memReg_1_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_900 = |_T_22 ? _memReg_1_branch_mask_T : _GEN_863; // @[fifo.scala 109:68 110:35]
  wire  _GEN_901 = _T_23 ? 1'h0 : _GEN_879; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_29 = memReg_2_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_30 = |_T_29; // @[fifo.scala 109:63]
  wire [4:0] _memReg_2_branch_mask_T = memReg_2_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_906 = |_T_29 ? _memReg_2_branch_mask_T : _GEN_864; // @[fifo.scala 109:68 110:35]
  wire  _GEN_907 = _T_30 ? 1'h0 : _GEN_880; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_36 = memReg_3_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_37 = |_T_36; // @[fifo.scala 109:63]
  wire [4:0] _memReg_3_branch_mask_T = memReg_3_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_912 = |_T_36 ? _memReg_3_branch_mask_T : _GEN_865; // @[fifo.scala 109:68 110:35]
  wire  _GEN_913 = _T_37 ? 1'h0 : _GEN_881; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_43 = memReg_4_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_44 = |_T_43; // @[fifo.scala 109:63]
  wire [4:0] _memReg_4_branch_mask_T = memReg_4_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_918 = |_T_43 ? _memReg_4_branch_mask_T : _GEN_866; // @[fifo.scala 109:68 110:35]
  wire  _GEN_919 = _T_44 ? 1'h0 : _GEN_882; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_50 = memReg_5_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_51 = |_T_50; // @[fifo.scala 109:63]
  wire [4:0] _memReg_5_branch_mask_T = memReg_5_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_924 = |_T_50 ? _memReg_5_branch_mask_T : _GEN_867; // @[fifo.scala 109:68 110:35]
  wire  _GEN_925 = _T_51 ? 1'h0 : _GEN_883; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_57 = memReg_6_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_58 = |_T_57; // @[fifo.scala 109:63]
  wire [4:0] _memReg_6_branch_mask_T = memReg_6_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_930 = |_T_57 ? _memReg_6_branch_mask_T : _GEN_868; // @[fifo.scala 109:68 110:35]
  wire  _GEN_931 = _T_58 ? 1'h0 : _GEN_884; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_64 = memReg_7_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_65 = |_T_64; // @[fifo.scala 109:63]
  wire [4:0] _memReg_7_branch_mask_T = memReg_7_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_936 = |_T_64 ? _memReg_7_branch_mask_T : _GEN_869; // @[fifo.scala 109:68 110:35]
  wire  _GEN_937 = _T_65 ? 1'h0 : _GEN_885; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_71 = memReg_8_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_72 = |_T_71; // @[fifo.scala 109:63]
  wire [4:0] _memReg_8_branch_mask_T = memReg_8_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_942 = |_T_71 ? _memReg_8_branch_mask_T : _GEN_870; // @[fifo.scala 109:68 110:35]
  wire  _GEN_943 = _T_72 ? 1'h0 : _GEN_886; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_78 = memReg_9_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_79 = |_T_78; // @[fifo.scala 109:63]
  wire [4:0] _memReg_9_branch_mask_T = memReg_9_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_948 = |_T_78 ? _memReg_9_branch_mask_T : _GEN_871; // @[fifo.scala 109:68 110:35]
  wire  _GEN_949 = _T_79 ? 1'h0 : _GEN_887; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_85 = memReg_10_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_86 = |_T_85; // @[fifo.scala 109:63]
  wire [4:0] _memReg_10_branch_mask_T = memReg_10_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_954 = |_T_85 ? _memReg_10_branch_mask_T : _GEN_872; // @[fifo.scala 109:68 110:35]
  wire  _GEN_955 = _T_86 ? 1'h0 : _GEN_888; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_92 = memReg_11_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_93 = |_T_92; // @[fifo.scala 109:63]
  wire [4:0] _memReg_11_branch_mask_T = memReg_11_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_960 = |_T_92 ? _memReg_11_branch_mask_T : _GEN_873; // @[fifo.scala 109:68 110:35]
  wire  _GEN_961 = _T_93 ? 1'h0 : _GEN_889; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_99 = memReg_12_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_100 = |_T_99; // @[fifo.scala 109:63]
  wire [4:0] _memReg_12_branch_mask_T = memReg_12_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_966 = |_T_99 ? _memReg_12_branch_mask_T : _GEN_874; // @[fifo.scala 109:68 110:35]
  wire  _GEN_967 = _T_100 ? 1'h0 : _GEN_890; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_106 = memReg_13_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_107 = |_T_106; // @[fifo.scala 109:63]
  wire [4:0] _memReg_13_branch_mask_T = memReg_13_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_972 = |_T_106 ? _memReg_13_branch_mask_T : _GEN_875; // @[fifo.scala 109:68 110:35]
  wire  _GEN_973 = _T_107 ? 1'h0 : _GEN_891; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_113 = memReg_14_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_114 = |_T_113; // @[fifo.scala 109:63]
  wire [4:0] _memReg_14_branch_mask_T = memReg_14_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_978 = |_T_113 ? _memReg_14_branch_mask_T : _GEN_876; // @[fifo.scala 109:68 110:35]
  wire  _GEN_979 = _T_114 ? 1'h0 : _GEN_892; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_120 = memReg_15_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_121 = |_T_120; // @[fifo.scala 109:63]
  wire [4:0] _memReg_15_branch_mask_T = memReg_15_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _T_124 = _GEN_525 & branchOps_branchMask; // @[utils.scala 92:27]
  wire  _T_125 = |_T_124; // @[utils.scala 92:51]
  wire [4:0] _read_data_branch_mask_T = _GEN_525 ^ branchOps_branchMask; // @[utils.scala 93:42]
  wire [4:0] _GEN_1022 = |_T_124 ? _read_data_branch_mask_T : _GEN_525; // @[utils.scala 92:56 93:27 96:27]
  wire [4:0] _GEN_1023 = _T_125 ? 5'h0 : _GEN_525; // @[utils.scala 101:56 102:27 106:27]
  wire  _GEN_1024 = _T_125 ? 1'h0 : _GEN_509; // @[utils.scala 101:56 103:28 107:28]
  wire [4:0] _GEN_1025 = branchOps_passed ? _GEN_1022 : _GEN_1023; // @[utils.scala 90:30]
  wire  _GEN_1026 = branchOps_passed ? _GEN_509 : _GEN_1024; // @[utils.scala 90:30 98:26]
  assign write_ready = ~fullReg; // @[fifo.scala 88:18]
  assign read_data_valid = _T_2 & _GEN_429; // @[fifo.scala 122:32]
  assign read_data_address = 4'hf == readPtr ? memReg_15_address : _GEN_444; // @[fifo.scala 86:{13,13}]
  assign read_data_core_instruction = 4'hf == readPtr ? memReg_15_core_instruction : _GEN_460; // @[fifo.scala 86:{13,13}]
  assign read_data_core_robAddr = 4'hf == readPtr ? memReg_15_core_robAddr : _GEN_476; // @[fifo.scala 86:{13,13}]
  assign read_data_core_prfDest = 4'hf == readPtr ? memReg_15_core_prfDest : _GEN_492; // @[fifo.scala 86:{13,13}]
  assign read_data_branch_valid = branchOps_valid ? _GEN_1026 : _GEN_509; // @[utils.scala 112:24 89:27]
  assign read_data_branch_mask = branchOps_valid ? _GEN_1025 : _GEN_525; // @[utils.scala 111:23 89:27]
  assign read_data_writeData_valid = 4'hf == readPtr ? memReg_15_writeData_valid : _GEN_540; // @[fifo.scala 86:{13,13}]
  assign read_data_writeData_data = 4'hf == readPtr ? memReg_15_writeData_data : _GEN_556; // @[fifo.scala 86:{13,13}]
  assign read_data_cacheLine_response = 4'hf == readPtr ? memReg_15_cacheLine_response : _GEN_588; // @[fifo.scala 86:{13,13}]
  assign isEmpty = emptyReg; // @[fifo.scala 89:11]
  always @(posedge clock) begin
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (branchOps_passed) begin // @[fifo.scala 108:32]
        memReg_0_branch_valid <= _GEN_878;
      end else if (_T_16) begin // @[fifo.scala 113:68]
        memReg_0_branch_valid <= 1'h0; // @[fifo.scala 114:36]
      end else begin
        memReg_0_branch_valid <= _GEN_878;
      end
    end else begin
      memReg_0_branch_valid <= _GEN_878;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (branchOps_passed) begin // @[fifo.scala 108:32]
        if (|_T_15) begin // @[fifo.scala 109:68]
          memReg_0_branch_mask <= _memReg_0_branch_mask_T; // @[fifo.scala 110:35]
        end else begin
          memReg_0_branch_mask <= _GEN_862;
        end
      end else begin
        memReg_0_branch_mask <= _GEN_862;
      end
    end else begin
      memReg_0_branch_mask <= _GEN_862;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_writeData_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_writeData_valid <= write_data_writeData_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_cacheLine_response <= 2'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_cacheLine_response <= write_data_cacheLine_response; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h1 | 4'h1 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_1_branch_valid <= _GEN_879;
        end else begin
          memReg_1_branch_valid <= _GEN_901;
        end
      end else begin
        memReg_1_branch_valid <= _GEN_879;
      end
    end else begin
      memReg_1_branch_valid <= _GEN_879;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h1 | 4'h1 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_1_branch_mask <= _GEN_900;
        end else begin
          memReg_1_branch_mask <= _GEN_863;
        end
      end else begin
        memReg_1_branch_mask <= _GEN_863;
      end
    end else begin
      memReg_1_branch_mask <= _GEN_863;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_writeData_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_writeData_valid <= write_data_writeData_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_cacheLine_response <= 2'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_cacheLine_response <= write_data_cacheLine_response; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h2 | 4'h2 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_2_branch_valid <= _GEN_880;
        end else begin
          memReg_2_branch_valid <= _GEN_907;
        end
      end else begin
        memReg_2_branch_valid <= _GEN_880;
      end
    end else begin
      memReg_2_branch_valid <= _GEN_880;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h2 | 4'h2 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_2_branch_mask <= _GEN_906;
        end else begin
          memReg_2_branch_mask <= _GEN_864;
        end
      end else begin
        memReg_2_branch_mask <= _GEN_864;
      end
    end else begin
      memReg_2_branch_mask <= _GEN_864;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_writeData_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_writeData_valid <= write_data_writeData_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_cacheLine_response <= 2'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_cacheLine_response <= write_data_cacheLine_response; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h3 | 4'h3 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_3_branch_valid <= _GEN_881;
        end else begin
          memReg_3_branch_valid <= _GEN_913;
        end
      end else begin
        memReg_3_branch_valid <= _GEN_881;
      end
    end else begin
      memReg_3_branch_valid <= _GEN_881;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h3 | 4'h3 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_3_branch_mask <= _GEN_912;
        end else begin
          memReg_3_branch_mask <= _GEN_865;
        end
      end else begin
        memReg_3_branch_mask <= _GEN_865;
      end
    end else begin
      memReg_3_branch_mask <= _GEN_865;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_writeData_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_writeData_valid <= write_data_writeData_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_cacheLine_response <= 2'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_cacheLine_response <= write_data_cacheLine_response; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h4 | 4'h4 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_4_branch_valid <= _GEN_882;
        end else begin
          memReg_4_branch_valid <= _GEN_919;
        end
      end else begin
        memReg_4_branch_valid <= _GEN_882;
      end
    end else begin
      memReg_4_branch_valid <= _GEN_882;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h4 | 4'h4 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_4_branch_mask <= _GEN_918;
        end else begin
          memReg_4_branch_mask <= _GEN_866;
        end
      end else begin
        memReg_4_branch_mask <= _GEN_866;
      end
    end else begin
      memReg_4_branch_mask <= _GEN_866;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_writeData_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_writeData_valid <= write_data_writeData_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_cacheLine_response <= 2'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_cacheLine_response <= write_data_cacheLine_response; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h5 | 4'h5 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_5_branch_valid <= _GEN_883;
        end else begin
          memReg_5_branch_valid <= _GEN_925;
        end
      end else begin
        memReg_5_branch_valid <= _GEN_883;
      end
    end else begin
      memReg_5_branch_valid <= _GEN_883;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h5 | 4'h5 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_5_branch_mask <= _GEN_924;
        end else begin
          memReg_5_branch_mask <= _GEN_867;
        end
      end else begin
        memReg_5_branch_mask <= _GEN_867;
      end
    end else begin
      memReg_5_branch_mask <= _GEN_867;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_writeData_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_writeData_valid <= write_data_writeData_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_cacheLine_response <= 2'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_cacheLine_response <= write_data_cacheLine_response; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h6 | 4'h6 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_6_branch_valid <= _GEN_884;
        end else begin
          memReg_6_branch_valid <= _GEN_931;
        end
      end else begin
        memReg_6_branch_valid <= _GEN_884;
      end
    end else begin
      memReg_6_branch_valid <= _GEN_884;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h6 | 4'h6 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_6_branch_mask <= _GEN_930;
        end else begin
          memReg_6_branch_mask <= _GEN_868;
        end
      end else begin
        memReg_6_branch_mask <= _GEN_868;
      end
    end else begin
      memReg_6_branch_mask <= _GEN_868;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_writeData_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_writeData_valid <= write_data_writeData_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_cacheLine_response <= 2'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_cacheLine_response <= write_data_cacheLine_response; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h7 | 4'h7 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_7_branch_valid <= _GEN_885;
        end else begin
          memReg_7_branch_valid <= _GEN_937;
        end
      end else begin
        memReg_7_branch_valid <= _GEN_885;
      end
    end else begin
      memReg_7_branch_valid <= _GEN_885;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h7 | 4'h7 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_7_branch_mask <= _GEN_936;
        end else begin
          memReg_7_branch_mask <= _GEN_869;
        end
      end else begin
        memReg_7_branch_mask <= _GEN_869;
      end
    end else begin
      memReg_7_branch_mask <= _GEN_869;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_writeData_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_writeData_valid <= write_data_writeData_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_cacheLine_response <= 2'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_cacheLine_response <= write_data_cacheLine_response; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h8 | 4'h8 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_8_branch_valid <= _GEN_886;
        end else begin
          memReg_8_branch_valid <= _GEN_943;
        end
      end else begin
        memReg_8_branch_valid <= _GEN_886;
      end
    end else begin
      memReg_8_branch_valid <= _GEN_886;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h8 | 4'h8 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_8_branch_mask <= _GEN_942;
        end else begin
          memReg_8_branch_mask <= _GEN_870;
        end
      end else begin
        memReg_8_branch_mask <= _GEN_870;
      end
    end else begin
      memReg_8_branch_mask <= _GEN_870;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_writeData_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_writeData_valid <= write_data_writeData_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_cacheLine_response <= 2'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_cacheLine_response <= write_data_cacheLine_response; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h9 | 4'h9 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_9_branch_valid <= _GEN_887;
        end else begin
          memReg_9_branch_valid <= _GEN_949;
        end
      end else begin
        memReg_9_branch_valid <= _GEN_887;
      end
    end else begin
      memReg_9_branch_valid <= _GEN_887;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'h9 | 4'h9 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_9_branch_mask <= _GEN_948;
        end else begin
          memReg_9_branch_mask <= _GEN_871;
        end
      end else begin
        memReg_9_branch_mask <= _GEN_871;
      end
    end else begin
      memReg_9_branch_mask <= _GEN_871;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_writeData_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_writeData_valid <= write_data_writeData_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_cacheLine_response <= 2'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_cacheLine_response <= write_data_cacheLine_response; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'ha | 4'ha <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_10_branch_valid <= _GEN_888;
        end else begin
          memReg_10_branch_valid <= _GEN_955;
        end
      end else begin
        memReg_10_branch_valid <= _GEN_888;
      end
    end else begin
      memReg_10_branch_valid <= _GEN_888;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'ha | 4'ha <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_10_branch_mask <= _GEN_954;
        end else begin
          memReg_10_branch_mask <= _GEN_872;
        end
      end else begin
        memReg_10_branch_mask <= _GEN_872;
      end
    end else begin
      memReg_10_branch_mask <= _GEN_872;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_writeData_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_writeData_valid <= write_data_writeData_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_cacheLine_response <= 2'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_cacheLine_response <= write_data_cacheLine_response; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'hb | 4'hb <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_11_branch_valid <= _GEN_889;
        end else begin
          memReg_11_branch_valid <= _GEN_961;
        end
      end else begin
        memReg_11_branch_valid <= _GEN_889;
      end
    end else begin
      memReg_11_branch_valid <= _GEN_889;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'hb | 4'hb <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_11_branch_mask <= _GEN_960;
        end else begin
          memReg_11_branch_mask <= _GEN_873;
        end
      end else begin
        memReg_11_branch_mask <= _GEN_873;
      end
    end else begin
      memReg_11_branch_mask <= _GEN_873;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_writeData_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_writeData_valid <= write_data_writeData_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_cacheLine_response <= 2'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_cacheLine_response <= write_data_cacheLine_response; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'hc | 4'hc <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_12_branch_valid <= _GEN_890;
        end else begin
          memReg_12_branch_valid <= _GEN_967;
        end
      end else begin
        memReg_12_branch_valid <= _GEN_890;
      end
    end else begin
      memReg_12_branch_valid <= _GEN_890;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'hc | 4'hc <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_12_branch_mask <= _GEN_966;
        end else begin
          memReg_12_branch_mask <= _GEN_874;
        end
      end else begin
        memReg_12_branch_mask <= _GEN_874;
      end
    end else begin
      memReg_12_branch_mask <= _GEN_874;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_writeData_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_writeData_valid <= write_data_writeData_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_cacheLine_response <= 2'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_cacheLine_response <= write_data_cacheLine_response; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'hd | 4'hd <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_13_branch_valid <= _GEN_891;
        end else begin
          memReg_13_branch_valid <= _GEN_973;
        end
      end else begin
        memReg_13_branch_valid <= _GEN_891;
      end
    end else begin
      memReg_13_branch_valid <= _GEN_891;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'hd | 4'hd <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_13_branch_mask <= _GEN_972;
        end else begin
          memReg_13_branch_mask <= _GEN_875;
        end
      end else begin
        memReg_13_branch_mask <= _GEN_875;
      end
    end else begin
      memReg_13_branch_mask <= _GEN_875;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_writeData_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_writeData_valid <= write_data_writeData_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_cacheLine_response <= 2'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_cacheLine_response <= write_data_cacheLine_response; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'he | 4'he <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_14_branch_valid <= _GEN_892;
        end else begin
          memReg_14_branch_valid <= _GEN_979;
        end
      end else begin
        memReg_14_branch_valid <= _GEN_892;
      end
    end else begin
      memReg_14_branch_valid <= _GEN_892;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 4'he | 4'he <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_14_branch_mask <= _GEN_978;
        end else begin
          memReg_14_branch_mask <= _GEN_876;
        end
      end else begin
        memReg_14_branch_mask <= _GEN_876;
      end
    end else begin
      memReg_14_branch_mask <= _GEN_876;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_writeData_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_writeData_valid <= write_data_writeData_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_cacheLine_response <= 2'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_cacheLine_response <= write_data_cacheLine_response; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_valid <= write_data_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (branchOps_passed) begin // @[fifo.scala 108:32]
        memReg_15_branch_valid <= _GEN_893;
      end else if (_T_121) begin // @[fifo.scala 113:68]
        memReg_15_branch_valid <= 1'h0; // @[fifo.scala 114:36]
      end else begin
        memReg_15_branch_valid <= _GEN_893;
      end
    end else begin
      memReg_15_branch_valid <= _GEN_893;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (branchOps_passed) begin // @[fifo.scala 108:32]
        if (|_T_120) begin // @[fifo.scala 109:68]
          memReg_15_branch_mask <= _memReg_15_branch_mask_T; // @[fifo.scala 110:35]
        end else begin
          memReg_15_branch_mask <= _GEN_877;
        end
      end else begin
        memReg_15_branch_mask <= _GEN_877;
      end
    end else begin
      memReg_15_branch_mask <= _GEN_877;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_writeData_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_writeData_valid <= write_data_writeData_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_cacheLine_response <= 2'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_cacheLine_response <= write_data_cacheLine_response; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 33:25]
      readPtr <= 4'h0; // @[fifo.scala 33:25]
    end else if (incrRead) begin // @[fifo.scala 35:15]
      if (readPtr == 4'hf) begin // @[fifo.scala 34:22]
        readPtr <= 4'h0;
      end else begin
        readPtr <= _nextVal_T_2;
      end
    end
    emptyReg <= reset | _GEN_27; // @[fifo.scala 43:{25,25}]
    if (reset) begin // @[fifo.scala 33:25]
      writePtr <= 4'h0; // @[fifo.scala 33:25]
    end else if (incrWrite) begin // @[fifo.scala 35:15]
      if (writePtr == 4'hf) begin // @[fifo.scala 34:22]
        writePtr <= 4'h0;
      end else begin
        writePtr <= _nextVal_T_5;
      end
    end
    if (reset) begin // @[fifo.scala 44:34]
      fullReg <= 1'h0; // @[fifo.scala 44:34]
    end else if (!(2'h0 == op)) begin // @[fifo.scala 49:14]
      if (2'h1 == op) begin // @[fifo.scala 49:14]
        if (~emptyReg) begin // @[fifo.scala 52:23]
          fullReg <= 1'h0; // @[fifo.scala 53:17]
        end
      end else if (2'h2 == op) begin // @[fifo.scala 49:14]
        fullReg <= _GEN_7;
      end else begin
        fullReg <= _GEN_16;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  memReg_0_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  memReg_0_address = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  memReg_0_core_instruction = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  memReg_0_core_robAddr = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  memReg_0_core_prfDest = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  memReg_0_branch_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  memReg_0_branch_mask = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  memReg_0_writeData_valid = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  memReg_0_writeData_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  memReg_0_cacheLine_response = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  memReg_1_valid = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  memReg_1_address = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  memReg_1_core_instruction = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  memReg_1_core_robAddr = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  memReg_1_core_prfDest = _RAND_14[5:0];
  _RAND_15 = {1{`RANDOM}};
  memReg_1_branch_valid = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  memReg_1_branch_mask = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  memReg_1_writeData_valid = _RAND_17[0:0];
  _RAND_18 = {2{`RANDOM}};
  memReg_1_writeData_data = _RAND_18[63:0];
  _RAND_19 = {1{`RANDOM}};
  memReg_1_cacheLine_response = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  memReg_2_valid = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  memReg_2_address = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  memReg_2_core_instruction = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  memReg_2_core_robAddr = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  memReg_2_core_prfDest = _RAND_24[5:0];
  _RAND_25 = {1{`RANDOM}};
  memReg_2_branch_valid = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  memReg_2_branch_mask = _RAND_26[4:0];
  _RAND_27 = {1{`RANDOM}};
  memReg_2_writeData_valid = _RAND_27[0:0];
  _RAND_28 = {2{`RANDOM}};
  memReg_2_writeData_data = _RAND_28[63:0];
  _RAND_29 = {1{`RANDOM}};
  memReg_2_cacheLine_response = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  memReg_3_valid = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  memReg_3_address = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  memReg_3_core_instruction = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  memReg_3_core_robAddr = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  memReg_3_core_prfDest = _RAND_34[5:0];
  _RAND_35 = {1{`RANDOM}};
  memReg_3_branch_valid = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  memReg_3_branch_mask = _RAND_36[4:0];
  _RAND_37 = {1{`RANDOM}};
  memReg_3_writeData_valid = _RAND_37[0:0];
  _RAND_38 = {2{`RANDOM}};
  memReg_3_writeData_data = _RAND_38[63:0];
  _RAND_39 = {1{`RANDOM}};
  memReg_3_cacheLine_response = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  memReg_4_valid = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  memReg_4_address = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  memReg_4_core_instruction = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  memReg_4_core_robAddr = _RAND_43[3:0];
  _RAND_44 = {1{`RANDOM}};
  memReg_4_core_prfDest = _RAND_44[5:0];
  _RAND_45 = {1{`RANDOM}};
  memReg_4_branch_valid = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  memReg_4_branch_mask = _RAND_46[4:0];
  _RAND_47 = {1{`RANDOM}};
  memReg_4_writeData_valid = _RAND_47[0:0];
  _RAND_48 = {2{`RANDOM}};
  memReg_4_writeData_data = _RAND_48[63:0];
  _RAND_49 = {1{`RANDOM}};
  memReg_4_cacheLine_response = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  memReg_5_valid = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  memReg_5_address = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  memReg_5_core_instruction = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  memReg_5_core_robAddr = _RAND_53[3:0];
  _RAND_54 = {1{`RANDOM}};
  memReg_5_core_prfDest = _RAND_54[5:0];
  _RAND_55 = {1{`RANDOM}};
  memReg_5_branch_valid = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  memReg_5_branch_mask = _RAND_56[4:0];
  _RAND_57 = {1{`RANDOM}};
  memReg_5_writeData_valid = _RAND_57[0:0];
  _RAND_58 = {2{`RANDOM}};
  memReg_5_writeData_data = _RAND_58[63:0];
  _RAND_59 = {1{`RANDOM}};
  memReg_5_cacheLine_response = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  memReg_6_valid = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  memReg_6_address = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  memReg_6_core_instruction = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  memReg_6_core_robAddr = _RAND_63[3:0];
  _RAND_64 = {1{`RANDOM}};
  memReg_6_core_prfDest = _RAND_64[5:0];
  _RAND_65 = {1{`RANDOM}};
  memReg_6_branch_valid = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  memReg_6_branch_mask = _RAND_66[4:0];
  _RAND_67 = {1{`RANDOM}};
  memReg_6_writeData_valid = _RAND_67[0:0];
  _RAND_68 = {2{`RANDOM}};
  memReg_6_writeData_data = _RAND_68[63:0];
  _RAND_69 = {1{`RANDOM}};
  memReg_6_cacheLine_response = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  memReg_7_valid = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  memReg_7_address = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  memReg_7_core_instruction = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  memReg_7_core_robAddr = _RAND_73[3:0];
  _RAND_74 = {1{`RANDOM}};
  memReg_7_core_prfDest = _RAND_74[5:0];
  _RAND_75 = {1{`RANDOM}};
  memReg_7_branch_valid = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  memReg_7_branch_mask = _RAND_76[4:0];
  _RAND_77 = {1{`RANDOM}};
  memReg_7_writeData_valid = _RAND_77[0:0];
  _RAND_78 = {2{`RANDOM}};
  memReg_7_writeData_data = _RAND_78[63:0];
  _RAND_79 = {1{`RANDOM}};
  memReg_7_cacheLine_response = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  memReg_8_valid = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  memReg_8_address = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  memReg_8_core_instruction = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  memReg_8_core_robAddr = _RAND_83[3:0];
  _RAND_84 = {1{`RANDOM}};
  memReg_8_core_prfDest = _RAND_84[5:0];
  _RAND_85 = {1{`RANDOM}};
  memReg_8_branch_valid = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  memReg_8_branch_mask = _RAND_86[4:0];
  _RAND_87 = {1{`RANDOM}};
  memReg_8_writeData_valid = _RAND_87[0:0];
  _RAND_88 = {2{`RANDOM}};
  memReg_8_writeData_data = _RAND_88[63:0];
  _RAND_89 = {1{`RANDOM}};
  memReg_8_cacheLine_response = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  memReg_9_valid = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  memReg_9_address = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  memReg_9_core_instruction = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  memReg_9_core_robAddr = _RAND_93[3:0];
  _RAND_94 = {1{`RANDOM}};
  memReg_9_core_prfDest = _RAND_94[5:0];
  _RAND_95 = {1{`RANDOM}};
  memReg_9_branch_valid = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  memReg_9_branch_mask = _RAND_96[4:0];
  _RAND_97 = {1{`RANDOM}};
  memReg_9_writeData_valid = _RAND_97[0:0];
  _RAND_98 = {2{`RANDOM}};
  memReg_9_writeData_data = _RAND_98[63:0];
  _RAND_99 = {1{`RANDOM}};
  memReg_9_cacheLine_response = _RAND_99[1:0];
  _RAND_100 = {1{`RANDOM}};
  memReg_10_valid = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  memReg_10_address = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  memReg_10_core_instruction = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  memReg_10_core_robAddr = _RAND_103[3:0];
  _RAND_104 = {1{`RANDOM}};
  memReg_10_core_prfDest = _RAND_104[5:0];
  _RAND_105 = {1{`RANDOM}};
  memReg_10_branch_valid = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  memReg_10_branch_mask = _RAND_106[4:0];
  _RAND_107 = {1{`RANDOM}};
  memReg_10_writeData_valid = _RAND_107[0:0];
  _RAND_108 = {2{`RANDOM}};
  memReg_10_writeData_data = _RAND_108[63:0];
  _RAND_109 = {1{`RANDOM}};
  memReg_10_cacheLine_response = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  memReg_11_valid = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  memReg_11_address = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  memReg_11_core_instruction = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  memReg_11_core_robAddr = _RAND_113[3:0];
  _RAND_114 = {1{`RANDOM}};
  memReg_11_core_prfDest = _RAND_114[5:0];
  _RAND_115 = {1{`RANDOM}};
  memReg_11_branch_valid = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  memReg_11_branch_mask = _RAND_116[4:0];
  _RAND_117 = {1{`RANDOM}};
  memReg_11_writeData_valid = _RAND_117[0:0];
  _RAND_118 = {2{`RANDOM}};
  memReg_11_writeData_data = _RAND_118[63:0];
  _RAND_119 = {1{`RANDOM}};
  memReg_11_cacheLine_response = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  memReg_12_valid = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  memReg_12_address = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  memReg_12_core_instruction = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  memReg_12_core_robAddr = _RAND_123[3:0];
  _RAND_124 = {1{`RANDOM}};
  memReg_12_core_prfDest = _RAND_124[5:0];
  _RAND_125 = {1{`RANDOM}};
  memReg_12_branch_valid = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  memReg_12_branch_mask = _RAND_126[4:0];
  _RAND_127 = {1{`RANDOM}};
  memReg_12_writeData_valid = _RAND_127[0:0];
  _RAND_128 = {2{`RANDOM}};
  memReg_12_writeData_data = _RAND_128[63:0];
  _RAND_129 = {1{`RANDOM}};
  memReg_12_cacheLine_response = _RAND_129[1:0];
  _RAND_130 = {1{`RANDOM}};
  memReg_13_valid = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  memReg_13_address = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  memReg_13_core_instruction = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  memReg_13_core_robAddr = _RAND_133[3:0];
  _RAND_134 = {1{`RANDOM}};
  memReg_13_core_prfDest = _RAND_134[5:0];
  _RAND_135 = {1{`RANDOM}};
  memReg_13_branch_valid = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  memReg_13_branch_mask = _RAND_136[4:0];
  _RAND_137 = {1{`RANDOM}};
  memReg_13_writeData_valid = _RAND_137[0:0];
  _RAND_138 = {2{`RANDOM}};
  memReg_13_writeData_data = _RAND_138[63:0];
  _RAND_139 = {1{`RANDOM}};
  memReg_13_cacheLine_response = _RAND_139[1:0];
  _RAND_140 = {1{`RANDOM}};
  memReg_14_valid = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  memReg_14_address = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  memReg_14_core_instruction = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  memReg_14_core_robAddr = _RAND_143[3:0];
  _RAND_144 = {1{`RANDOM}};
  memReg_14_core_prfDest = _RAND_144[5:0];
  _RAND_145 = {1{`RANDOM}};
  memReg_14_branch_valid = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  memReg_14_branch_mask = _RAND_146[4:0];
  _RAND_147 = {1{`RANDOM}};
  memReg_14_writeData_valid = _RAND_147[0:0];
  _RAND_148 = {2{`RANDOM}};
  memReg_14_writeData_data = _RAND_148[63:0];
  _RAND_149 = {1{`RANDOM}};
  memReg_14_cacheLine_response = _RAND_149[1:0];
  _RAND_150 = {1{`RANDOM}};
  memReg_15_valid = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  memReg_15_address = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  memReg_15_core_instruction = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  memReg_15_core_robAddr = _RAND_153[3:0];
  _RAND_154 = {1{`RANDOM}};
  memReg_15_core_prfDest = _RAND_154[5:0];
  _RAND_155 = {1{`RANDOM}};
  memReg_15_branch_valid = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  memReg_15_branch_mask = _RAND_156[4:0];
  _RAND_157 = {1{`RANDOM}};
  memReg_15_writeData_valid = _RAND_157[0:0];
  _RAND_158 = {2{`RANDOM}};
  memReg_15_writeData_data = _RAND_158[63:0];
  _RAND_159 = {1{`RANDOM}};
  memReg_15_cacheLine_response = _RAND_159[1:0];
  _RAND_160 = {1{`RANDOM}};
  readPtr = _RAND_160[3:0];
  _RAND_161 = {1{`RANDOM}};
  emptyReg = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  writePtr = _RAND_162[3:0];
  _RAND_163 = {1{`RANDOM}};
  fullReg = _RAND_163[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module requestScheduler(
  input         clock,
  input         reset,
  input         requestIn_valid,
  input  [31:0] requestIn_address,
  input  [31:0] requestIn_core_instruction,
  input  [3:0]  requestIn_core_robAddr,
  input  [5:0]  requestIn_core_prfDest,
  input  [4:0]  requestIn_branch_mask,
  output        canAllocate,
  output        requestOut_valid,
  output [31:0] requestOut_address,
  output [31:0] requestOut_core_instruction,
  output [3:0]  requestOut_core_robAddr,
  output [5:0]  requestOut_core_prfDest,
  output        requestOut_branch_valid,
  output [4:0]  requestOut_branch_mask,
  output        requestOut_writeData_valid,
  output [63:0] requestOut_writeData_data,
  output        controlSignal_isSpeculative,
  input         controlSignal_inorderReady,
  input         controlSignal_speculativeReady,
  output        fenceReady,
  input         branchOps_valid,
  input  [4:0]  branchOps_branchMask,
  input         branchOps_passed
);
  wire  inorderQueue_clock; // @[requestScheduler.scala 30:28]
  wire  inorderQueue_reset; // @[requestScheduler.scala 30:28]
  wire  inorderQueue_write_ready; // @[requestScheduler.scala 30:28]
  wire  inorderQueue_write_data_valid; // @[requestScheduler.scala 30:28]
  wire [31:0] inorderQueue_write_data_address; // @[requestScheduler.scala 30:28]
  wire [31:0] inorderQueue_write_data_core_instruction; // @[requestScheduler.scala 30:28]
  wire [3:0] inorderQueue_write_data_core_robAddr; // @[requestScheduler.scala 30:28]
  wire [5:0] inorderQueue_write_data_core_prfDest; // @[requestScheduler.scala 30:28]
  wire  inorderQueue_write_data_branch_valid; // @[requestScheduler.scala 30:28]
  wire [4:0] inorderQueue_write_data_branch_mask; // @[requestScheduler.scala 30:28]
  wire  inorderQueue_read_ready; // @[requestScheduler.scala 30:28]
  wire  inorderQueue_read_data_valid; // @[requestScheduler.scala 30:28]
  wire [31:0] inorderQueue_read_data_address; // @[requestScheduler.scala 30:28]
  wire [31:0] inorderQueue_read_data_core_instruction; // @[requestScheduler.scala 30:28]
  wire [3:0] inorderQueue_read_data_core_robAddr; // @[requestScheduler.scala 30:28]
  wire [5:0] inorderQueue_read_data_core_prfDest; // @[requestScheduler.scala 30:28]
  wire  inorderQueue_read_data_branch_valid; // @[requestScheduler.scala 30:28]
  wire [4:0] inorderQueue_read_data_branch_mask; // @[requestScheduler.scala 30:28]
  wire  inorderQueue_isEmpty; // @[requestScheduler.scala 30:28]
  wire  inorderQueue_branchOps_valid; // @[requestScheduler.scala 30:28]
  wire [4:0] inorderQueue_branchOps_branchMask; // @[requestScheduler.scala 30:28]
  wire  inorderQueue_branchOps_passed; // @[requestScheduler.scala 30:28]
  wire [31:0] inorderQueue_checkAddress; // @[requestScheduler.scala 30:28]
  wire  inorderQueue_matchFound; // @[requestScheduler.scala 30:28]
  wire  speculativeQueue_clock; // @[requestScheduler.scala 35:32]
  wire  speculativeQueue_reset; // @[requestScheduler.scala 35:32]
  wire  speculativeQueue_write_ready; // @[requestScheduler.scala 35:32]
  wire  speculativeQueue_write_data_valid; // @[requestScheduler.scala 35:32]
  wire [31:0] speculativeQueue_write_data_address; // @[requestScheduler.scala 35:32]
  wire [31:0] speculativeQueue_write_data_core_instruction; // @[requestScheduler.scala 35:32]
  wire [3:0] speculativeQueue_write_data_core_robAddr; // @[requestScheduler.scala 35:32]
  wire [5:0] speculativeQueue_write_data_core_prfDest; // @[requestScheduler.scala 35:32]
  wire  speculativeQueue_write_data_branch_valid; // @[requestScheduler.scala 35:32]
  wire [4:0] speculativeQueue_write_data_branch_mask; // @[requestScheduler.scala 35:32]
  wire  speculativeQueue_write_data_writeData_valid; // @[requestScheduler.scala 35:32]
  wire [63:0] speculativeQueue_write_data_writeData_data; // @[requestScheduler.scala 35:32]
  wire [1:0] speculativeQueue_write_data_cacheLine_response; // @[requestScheduler.scala 35:32]
  wire  speculativeQueue_read_ready; // @[requestScheduler.scala 35:32]
  wire  speculativeQueue_read_data_valid; // @[requestScheduler.scala 35:32]
  wire [31:0] speculativeQueue_read_data_address; // @[requestScheduler.scala 35:32]
  wire [31:0] speculativeQueue_read_data_core_instruction; // @[requestScheduler.scala 35:32]
  wire [3:0] speculativeQueue_read_data_core_robAddr; // @[requestScheduler.scala 35:32]
  wire [5:0] speculativeQueue_read_data_core_prfDest; // @[requestScheduler.scala 35:32]
  wire  speculativeQueue_read_data_branch_valid; // @[requestScheduler.scala 35:32]
  wire [4:0] speculativeQueue_read_data_branch_mask; // @[requestScheduler.scala 35:32]
  wire  speculativeQueue_read_data_writeData_valid; // @[requestScheduler.scala 35:32]
  wire [63:0] speculativeQueue_read_data_writeData_data; // @[requestScheduler.scala 35:32]
  wire [1:0] speculativeQueue_read_data_cacheLine_response; // @[requestScheduler.scala 35:32]
  wire  speculativeQueue_isEmpty; // @[requestScheduler.scala 35:32]
  wire  speculativeQueue_branchOps_valid; // @[requestScheduler.scala 35:32]
  wire [4:0] speculativeQueue_branchOps_branchMask; // @[requestScheduler.scala 35:32]
  wire  speculativeQueue_branchOps_passed; // @[requestScheduler.scala 35:32]
  wire  speculativeEntryWire = requestIn_core_instruction[6:2] == 5'h0 & requestIn_address != 32'h40600000; // @[requestScheduler.scala 47:89]
  wire [4:0] _T_2 = requestIn_branch_mask & branchOps_branchMask; // @[utils.scala 92:27]
  wire  _T_3 = |_T_2; // @[utils.scala 92:51]
  wire [4:0] _inorderQueue_write_data_branch_mask_T = requestIn_branch_mask ^ branchOps_branchMask; // @[utils.scala 93:42]
  wire [4:0] _GEN_0 = |_T_2 ? _inorderQueue_write_data_branch_mask_T : requestIn_branch_mask; // @[utils.scala 92:56 93:27 96:27]
  wire [4:0] _GEN_1 = _T_3 ? 5'h0 : requestIn_branch_mask; // @[utils.scala 101:56 102:27 106:27]
  wire  _GEN_2 = _T_3 ? 1'h0 : 1'h1; // @[utils.scala 101:56 103:28 107:28]
  wire [4:0] _GEN_3 = branchOps_passed ? _GEN_0 : _GEN_1; // @[utils.scala 90:30]
  wire  _GEN_4 = branchOps_passed | _GEN_2; // @[utils.scala 90:30 98:26]
  wire [4:0] _GEN_5 = branchOps_valid ? _GEN_3 : requestIn_branch_mask; // @[utils.scala 111:23 89:27]
  wire  _GEN_6 = branchOps_valid ? _GEN_4 : 1'h1; // @[utils.scala 112:24 89:27]
  wire [4:0] _GEN_26 = speculativeEntryWire ? _GEN_5 : 5'h0; // @[requestScheduler.scala 54:38 utils.scala 49:41]
  wire  _GEN_27 = speculativeEntryWire & _GEN_6; // @[requestScheduler.scala 54:38 utils.scala 48:41]
  wire [5:0] _GEN_28 = speculativeEntryWire ? requestIn_core_prfDest : 6'h0; // @[requestScheduler.scala 54:38 55:35 utils.scala 49:41]
  wire [3:0] _GEN_29 = speculativeEntryWire ? requestIn_core_robAddr : 4'h0; // @[requestScheduler.scala 54:38 55:35 utils.scala 49:41]
  wire [31:0] _GEN_30 = speculativeEntryWire ? requestIn_core_instruction : 32'h0; // @[requestScheduler.scala 54:38 55:35 utils.scala 49:41]
  wire [31:0] _GEN_31 = speculativeEntryWire ? requestIn_address : 32'h0; // @[requestScheduler.scala 54:38 55:35 utils.scala 49:41]
  wire  _GEN_32 = speculativeEntryWire & requestIn_valid; // @[requestScheduler.scala 54:38 55:35 utils.scala 48:41]
  wire [4:0] _GEN_38 = speculativeEntryWire ? 5'h0 : _GEN_5; // @[requestScheduler.scala 54:38 utils.scala 49:41]
  wire  _GEN_39 = speculativeEntryWire ? 1'h0 : _GEN_6; // @[requestScheduler.scala 54:38 utils.scala 48:41]
  wire [5:0] _GEN_40 = speculativeEntryWire ? 6'h0 : requestIn_core_prfDest; // @[requestScheduler.scala 54:38 utils.scala 49:41 requestScheduler.scala 58:31]
  wire [3:0] _GEN_41 = speculativeEntryWire ? 4'h0 : requestIn_core_robAddr; // @[requestScheduler.scala 54:38 utils.scala 49:41 requestScheduler.scala 58:31]
  wire [31:0] _GEN_42 = speculativeEntryWire ? 32'h0 : requestIn_core_instruction; // @[requestScheduler.scala 54:38 utils.scala 49:41 requestScheduler.scala 58:31]
  wire [31:0] _GEN_43 = speculativeEntryWire ? 32'h0 : requestIn_address; // @[requestScheduler.scala 54:38 utils.scala 49:41 requestScheduler.scala 58:31]
  wire  _GEN_44 = speculativeEntryWire ? 1'h0 : requestIn_valid; // @[requestScheduler.scala 54:38 utils.scala 48:41 requestScheduler.scala 58:31]
  wire [4:0] _GEN_50 = speculativeEntryWire & inorderQueue_matchFound ? _GEN_5 : _GEN_38; // @[requestScheduler.scala 51:58]
  wire  _GEN_51 = speculativeEntryWire & inorderQueue_matchFound ? _GEN_6 : _GEN_39; // @[requestScheduler.scala 51:58]
  wire [5:0] _GEN_52 = speculativeEntryWire & inorderQueue_matchFound ? requestIn_core_prfDest : _GEN_40; // @[requestScheduler.scala 51:58 52:31]
  wire [3:0] _GEN_53 = speculativeEntryWire & inorderQueue_matchFound ? requestIn_core_robAddr : _GEN_41; // @[requestScheduler.scala 51:58 52:31]
  wire [31:0] _GEN_54 = speculativeEntryWire & inorderQueue_matchFound ? requestIn_core_instruction : _GEN_42; // @[requestScheduler.scala 51:58 52:31]
  wire [31:0] _GEN_55 = speculativeEntryWire & inorderQueue_matchFound ? requestIn_address : _GEN_43; // @[requestScheduler.scala 51:58 52:31]
  wire  _GEN_56 = speculativeEntryWire & inorderQueue_matchFound ? requestIn_valid : _GEN_44; // @[requestScheduler.scala 51:58 52:31]
  wire [4:0] _GEN_62 = speculativeEntryWire & inorderQueue_matchFound ? 5'h0 : _GEN_26; // @[requestScheduler.scala 51:58 utils.scala 49:41]
  wire  _GEN_63 = speculativeEntryWire & inorderQueue_matchFound ? 1'h0 : _GEN_27; // @[requestScheduler.scala 51:58 utils.scala 48:41]
  wire [5:0] _GEN_64 = speculativeEntryWire & inorderQueue_matchFound ? 6'h0 : _GEN_28; // @[requestScheduler.scala 51:58 utils.scala 49:41]
  wire [3:0] _GEN_65 = speculativeEntryWire & inorderQueue_matchFound ? 4'h0 : _GEN_29; // @[requestScheduler.scala 51:58 utils.scala 49:41]
  wire [31:0] _GEN_66 = speculativeEntryWire & inorderQueue_matchFound ? 32'h0 : _GEN_30; // @[requestScheduler.scala 51:58 utils.scala 49:41]
  wire [31:0] _GEN_67 = speculativeEntryWire & inorderQueue_matchFound ? 32'h0 : _GEN_31; // @[requestScheduler.scala 51:58 utils.scala 49:41]
  wire  _GEN_68 = speculativeEntryWire & inorderQueue_matchFound ? 1'h0 : _GEN_32; // @[requestScheduler.scala 51:58 utils.scala 48:41]
  wire  _speculativeBranchResolved_T_1 = |speculativeQueue_read_data_branch_mask[3:0]; // @[requestScheduler.scala 73:92]
  wire  _speculativeBranchResolved_T_3 = ~speculativeQueue_isEmpty; // @[requestScheduler.scala 73:99]
  wire  speculativeBranchResolved = ~(|speculativeQueue_read_data_branch_mask[3:0]) & ~speculativeQueue_isEmpty; // @[requestScheduler.scala 73:96]
  wire  speculativeBranchInvalidated = ~speculativeQueue_read_data_branch_valid & _speculativeBranchResolved_T_1 &
    _speculativeBranchResolved_T_3; // @[requestScheduler.scala 74:142]
  wire  _inorderBranchResolved_T_1 = |inorderQueue_read_data_branch_mask[3:0]; // @[requestScheduler.scala 75:84]
  wire  _inorderBranchResolved_T_3 = ~inorderQueue_isEmpty; // @[requestScheduler.scala 75:91]
  wire  inorderBranchResolved = ~(|inorderQueue_read_data_branch_mask[3:0]) & ~inorderQueue_isEmpty; // @[requestScheduler.scala 75:88]
  wire  inorderBranchInvalidated = ~inorderQueue_read_data_branch_valid & _inorderBranchResolved_T_1 &
    _inorderBranchResolved_T_3; // @[requestScheduler.scala 76:130]
  wire [1:0] _T_18 = {controlSignal_inorderReady,controlSignal_speculativeReady}; // @[requestScheduler.scala 79:39]
  wire  _T_22 = _speculativeBranchResolved_T_3 | speculativeBranchInvalidated; // @[requestScheduler.scala 82:40]
  wire  _GEN_93 = (_speculativeBranchResolved_T_3 | speculativeBranchInvalidated) & _speculativeBranchResolved_T_3; // @[requestScheduler.scala 44:31 82:72 83:38]
  wire  _GEN_95 = (_speculativeBranchResolved_T_3 | speculativeBranchInvalidated) & speculativeQueue_read_data_valid; // @[requestScheduler.scala 82:72 85:22 utils.scala 48:41]
  wire [31:0] _GEN_96 = _speculativeBranchResolved_T_3 | speculativeBranchInvalidated ?
    speculativeQueue_read_data_address : 32'h0; // @[requestScheduler.scala 82:72 85:22 utils.scala 49:41]
  wire [31:0] _GEN_97 = _speculativeBranchResolved_T_3 | speculativeBranchInvalidated ?
    speculativeQueue_read_data_core_instruction : 32'h0; // @[requestScheduler.scala 82:72 85:22 utils.scala 49:41]
  wire [3:0] _GEN_98 = _speculativeBranchResolved_T_3 | speculativeBranchInvalidated ?
    speculativeQueue_read_data_core_robAddr : 4'h0; // @[requestScheduler.scala 82:72 85:22 utils.scala 49:41]
  wire [5:0] _GEN_99 = _speculativeBranchResolved_T_3 | speculativeBranchInvalidated ?
    speculativeQueue_read_data_core_prfDest : 6'h0; // @[requestScheduler.scala 82:72 85:22 utils.scala 49:41]
  wire  _GEN_100 = (_speculativeBranchResolved_T_3 | speculativeBranchInvalidated) &
    speculativeQueue_read_data_branch_valid; // @[requestScheduler.scala 82:72 85:22 utils.scala 48:41]
  wire [4:0] _GEN_101 = _speculativeBranchResolved_T_3 | speculativeBranchInvalidated ?
    speculativeQueue_read_data_branch_mask : 5'h0; // @[requestScheduler.scala 82:72 85:22 utils.scala 49:41]
  wire  _GEN_102 = (_speculativeBranchResolved_T_3 | speculativeBranchInvalidated) &
    speculativeQueue_read_data_writeData_valid; // @[requestScheduler.scala 82:72 85:22 utils.scala 48:41]
  wire [63:0] _GEN_103 = _speculativeBranchResolved_T_3 | speculativeBranchInvalidated ?
    speculativeQueue_read_data_writeData_data : 64'h0; // @[requestScheduler.scala 82:72 85:22 utils.scala 49:41]
  wire  _T_24 = inorderBranchResolved | inorderBranchInvalidated; // @[requestScheduler.scala 89:36]
  wire  _GEN_107 = (inorderBranchResolved | inorderBranchInvalidated) & _inorderBranchResolved_T_3; // @[requestScheduler.scala 41:27 89:64 90:35]
  wire  _GEN_109 = (inorderBranchResolved | inorderBranchInvalidated) & inorderQueue_read_data_valid; // @[requestScheduler.scala 89:64 92:22 utils.scala 48:41]
  wire [31:0] _GEN_110 = inorderBranchResolved | inorderBranchInvalidated ? inorderQueue_read_data_address : 32'h0; // @[requestScheduler.scala 89:64 92:22 utils.scala 49:41]
  wire [31:0] _GEN_111 = inorderBranchResolved | inorderBranchInvalidated ? inorderQueue_read_data_core_instruction : 32'h0
    ; // @[requestScheduler.scala 89:64 92:22 utils.scala 49:41]
  wire [3:0] _GEN_112 = inorderBranchResolved | inorderBranchInvalidated ? inorderQueue_read_data_core_robAddr : 4'h0; // @[requestScheduler.scala 89:64 92:22 utils.scala 49:41]
  wire [5:0] _GEN_113 = inorderBranchResolved | inorderBranchInvalidated ? inorderQueue_read_data_core_prfDest : 6'h0; // @[requestScheduler.scala 89:64 92:22 utils.scala 49:41]
  wire  _GEN_114 = (inorderBranchResolved | inorderBranchInvalidated) & inorderQueue_read_data_branch_valid; // @[requestScheduler.scala 89:64 92:22 utils.scala 48:41]
  wire [4:0] _GEN_115 = inorderBranchResolved | inorderBranchInvalidated ? inorderQueue_read_data_branch_mask : 5'h0; // @[requestScheduler.scala 89:64 92:22 utils.scala 49:41]
  wire  _GEN_137 = _T_24 ? 1'h0 : _T_22; // @[requestScheduler.scala 101:71 104:40]
  wire  _GEN_138 = _T_24 ? inorderQueue_read_data_valid : _GEN_95; // @[requestScheduler.scala 101:71 105:22]
  wire [31:0] _GEN_139 = _T_24 ? inorderQueue_read_data_address : _GEN_96; // @[requestScheduler.scala 101:71 105:22]
  wire [31:0] _GEN_140 = _T_24 ? inorderQueue_read_data_core_instruction : _GEN_97; // @[requestScheduler.scala 101:71 105:22]
  wire [3:0] _GEN_141 = _T_24 ? inorderQueue_read_data_core_robAddr : _GEN_98; // @[requestScheduler.scala 101:71 105:22]
  wire [5:0] _GEN_142 = _T_24 ? inorderQueue_read_data_core_prfDest : _GEN_99; // @[requestScheduler.scala 101:71 105:22]
  wire  _GEN_143 = _T_24 ? inorderQueue_read_data_branch_valid : _GEN_100; // @[requestScheduler.scala 101:71 105:22]
  wire [4:0] _GEN_144 = _T_24 ? inorderQueue_read_data_branch_mask : _GEN_101; // @[requestScheduler.scala 101:71 105:22]
  wire  _GEN_145 = _T_24 ? 1'h0 : _GEN_102; // @[requestScheduler.scala 101:71 105:22]
  wire [63:0] _GEN_146 = _T_24 ? 64'h0 : _GEN_103; // @[requestScheduler.scala 101:71 105:22]
  wire  _GEN_150 = _T_24 ? 1'h0 : _GEN_93; // @[requestScheduler.scala 101:71 44:31]
  wire  _GEN_151 = speculativeBranchResolved | speculativeBranchInvalidated ? _speculativeBranchResolved_T_3 : _GEN_150; // @[requestScheduler.scala 96:72 98:38]
  wire  _GEN_152 = speculativeBranchResolved | speculativeBranchInvalidated | _GEN_137; // @[requestScheduler.scala 96:72 99:40]
  wire  _GEN_153 = speculativeBranchResolved | speculativeBranchInvalidated ? speculativeQueue_read_data_valid :
    _GEN_138; // @[requestScheduler.scala 100:22 96:72]
  wire [31:0] _GEN_154 = speculativeBranchResolved | speculativeBranchInvalidated ? speculativeQueue_read_data_address
     : _GEN_139; // @[requestScheduler.scala 100:22 96:72]
  wire [31:0] _GEN_155 = speculativeBranchResolved | speculativeBranchInvalidated ?
    speculativeQueue_read_data_core_instruction : _GEN_140; // @[requestScheduler.scala 100:22 96:72]
  wire [3:0] _GEN_156 = speculativeBranchResolved | speculativeBranchInvalidated ?
    speculativeQueue_read_data_core_robAddr : _GEN_141; // @[requestScheduler.scala 100:22 96:72]
  wire [5:0] _GEN_157 = speculativeBranchResolved | speculativeBranchInvalidated ?
    speculativeQueue_read_data_core_prfDest : _GEN_142; // @[requestScheduler.scala 100:22 96:72]
  wire  _GEN_158 = speculativeBranchResolved | speculativeBranchInvalidated ? speculativeQueue_read_data_branch_valid :
    _GEN_143; // @[requestScheduler.scala 100:22 96:72]
  wire [4:0] _GEN_159 = speculativeBranchResolved | speculativeBranchInvalidated ?
    speculativeQueue_read_data_branch_mask : _GEN_144; // @[requestScheduler.scala 100:22 96:72]
  wire  _GEN_160 = speculativeBranchResolved | speculativeBranchInvalidated ? speculativeQueue_read_data_writeData_valid
     : _GEN_145; // @[requestScheduler.scala 100:22 96:72]
  wire [63:0] _GEN_161 = speculativeBranchResolved | speculativeBranchInvalidated ?
    speculativeQueue_read_data_writeData_data : _GEN_146; // @[requestScheduler.scala 100:22 96:72]
  wire  _GEN_165 = speculativeBranchResolved | speculativeBranchInvalidated ? 1'h0 : _GEN_107; // @[requestScheduler.scala 41:27 96:72]
  wire  _GEN_167 = 2'h3 == _T_18 & _GEN_152; // @[requestScheduler.scala 27:31 79:73]
  wire  _GEN_168 = 2'h3 == _T_18 & _GEN_153; // @[requestScheduler.scala 79:73 utils.scala 48:41]
  wire [31:0] _GEN_169 = 2'h3 == _T_18 ? _GEN_154 : 32'h0; // @[requestScheduler.scala 79:73 utils.scala 49:41]
  wire [31:0] _GEN_170 = 2'h3 == _T_18 ? _GEN_155 : 32'h0; // @[requestScheduler.scala 79:73 utils.scala 49:41]
  wire [3:0] _GEN_171 = 2'h3 == _T_18 ? _GEN_156 : 4'h0; // @[requestScheduler.scala 79:73 utils.scala 49:41]
  wire [5:0] _GEN_172 = 2'h3 == _T_18 ? _GEN_157 : 6'h0; // @[requestScheduler.scala 79:73 utils.scala 49:41]
  wire  _GEN_173 = 2'h3 == _T_18 & _GEN_158; // @[requestScheduler.scala 79:73 utils.scala 48:41]
  wire [4:0] _GEN_174 = 2'h3 == _T_18 ? _GEN_159 : 5'h0; // @[requestScheduler.scala 79:73 utils.scala 49:41]
  wire  _GEN_175 = 2'h3 == _T_18 & _GEN_160; // @[requestScheduler.scala 79:73 utils.scala 48:41]
  wire [63:0] _GEN_176 = 2'h3 == _T_18 ? _GEN_161 : 64'h0; // @[requestScheduler.scala 79:73 utils.scala 49:41]
  wire  _GEN_180 = 2'h3 == _T_18 & _GEN_165; // @[requestScheduler.scala 41:27 79:73]
  wire  _GEN_181 = 2'h2 == _T_18 ? _GEN_107 : _GEN_180; // @[requestScheduler.scala 79:73]
  wire  _GEN_182 = 2'h2 == _T_18 ? 1'h0 : _GEN_167; // @[requestScheduler.scala 79:73]
  wire  _GEN_183 = 2'h2 == _T_18 ? _GEN_109 : _GEN_168; // @[requestScheduler.scala 79:73]
  wire [31:0] _GEN_184 = 2'h2 == _T_18 ? _GEN_110 : _GEN_169; // @[requestScheduler.scala 79:73]
  wire [31:0] _GEN_185 = 2'h2 == _T_18 ? _GEN_111 : _GEN_170; // @[requestScheduler.scala 79:73]
  wire [3:0] _GEN_186 = 2'h2 == _T_18 ? _GEN_112 : _GEN_171; // @[requestScheduler.scala 79:73]
  wire [5:0] _GEN_187 = 2'h2 == _T_18 ? _GEN_113 : _GEN_172; // @[requestScheduler.scala 79:73]
  wire  _GEN_188 = 2'h2 == _T_18 ? _GEN_114 : _GEN_173; // @[requestScheduler.scala 79:73]
  wire [4:0] _GEN_189 = 2'h2 == _T_18 ? _GEN_115 : _GEN_174; // @[requestScheduler.scala 79:73]
  wire  _GEN_190 = 2'h2 == _T_18 ? 1'h0 : _GEN_175; // @[requestScheduler.scala 79:73]
  wire [63:0] _GEN_191 = 2'h2 == _T_18 ? 64'h0 : _GEN_176; // @[requestScheduler.scala 79:73]
  wire  _GEN_195 = 2'h2 == _T_18 ? 1'h0 : 2'h3 == _T_18 & _GEN_151; // @[requestScheduler.scala 44:31 79:73]
  wire  _GEN_196 = 2'h1 == _T_18 ? _GEN_93 : _GEN_195; // @[requestScheduler.scala 79:73]
  wire  _GEN_197 = 2'h1 == _T_18 ? _T_22 : _GEN_182; // @[requestScheduler.scala 79:73]
  wire  _GEN_198 = 2'h1 == _T_18 ? _GEN_95 : _GEN_183; // @[requestScheduler.scala 79:73]
  wire [31:0] _GEN_199 = 2'h1 == _T_18 ? _GEN_96 : _GEN_184; // @[requestScheduler.scala 79:73]
  wire [31:0] _GEN_200 = 2'h1 == _T_18 ? _GEN_97 : _GEN_185; // @[requestScheduler.scala 79:73]
  wire [3:0] _GEN_201 = 2'h1 == _T_18 ? _GEN_98 : _GEN_186; // @[requestScheduler.scala 79:73]
  wire [5:0] _GEN_202 = 2'h1 == _T_18 ? _GEN_99 : _GEN_187; // @[requestScheduler.scala 79:73]
  wire  _GEN_203 = 2'h1 == _T_18 ? _GEN_100 : _GEN_188; // @[requestScheduler.scala 79:73]
  wire [4:0] _GEN_204 = 2'h1 == _T_18 ? _GEN_101 : _GEN_189; // @[requestScheduler.scala 79:73]
  wire  _GEN_205 = 2'h1 == _T_18 ? _GEN_102 : _GEN_190; // @[requestScheduler.scala 79:73]
  wire [63:0] _GEN_206 = 2'h1 == _T_18 ? _GEN_103 : _GEN_191; // @[requestScheduler.scala 79:73]
  wire  _GEN_210 = 2'h1 == _T_18 ? 1'h0 : _GEN_181; // @[requestScheduler.scala 41:27 79:73]
  wire  _GEN_211 = 2'h0 == _T_18 ? 1'h0 : _GEN_196; // @[requestScheduler.scala 44:31 79:73]
  wire  _GEN_212 = 2'h0 == _T_18 ? 1'h0 : _GEN_197; // @[requestScheduler.scala 27:31 79:73]
  wire  _GEN_213 = 2'h0 == _T_18 ? 1'h0 : _GEN_198; // @[requestScheduler.scala 79:73 utils.scala 48:41]
  wire [31:0] _GEN_214 = 2'h0 == _T_18 ? 32'h0 : _GEN_199; // @[requestScheduler.scala 79:73 utils.scala 49:41]
  wire [31:0] _GEN_215 = 2'h0 == _T_18 ? 32'h0 : _GEN_200; // @[requestScheduler.scala 79:73 utils.scala 49:41]
  wire [3:0] _GEN_216 = 2'h0 == _T_18 ? 4'h0 : _GEN_201; // @[requestScheduler.scala 79:73 utils.scala 49:41]
  wire [5:0] _GEN_217 = 2'h0 == _T_18 ? 6'h0 : _GEN_202; // @[requestScheduler.scala 79:73 utils.scala 49:41]
  wire  _GEN_218 = 2'h0 == _T_18 ? 1'h0 : _GEN_203; // @[requestScheduler.scala 79:73 utils.scala 48:41]
  wire [4:0] _GEN_219 = 2'h0 == _T_18 ? 5'h0 : _GEN_204; // @[requestScheduler.scala 79:73 utils.scala 49:41]
  wire  _GEN_220 = 2'h0 == _T_18 ? 1'h0 : _GEN_205; // @[requestScheduler.scala 79:73 utils.scala 48:41]
  wire [63:0] _GEN_221 = 2'h0 == _T_18 ? 64'h0 : _GEN_206; // @[requestScheduler.scala 79:73 utils.scala 49:41]
  wire  _GEN_225 = 2'h0 == _T_18 ? 1'h0 : _GEN_210; // @[requestScheduler.scala 41:27 79:73]
  fifoWithAddrCheck inorderQueue ( // @[requestScheduler.scala 30:28]
    .clock(inorderQueue_clock),
    .reset(inorderQueue_reset),
    .write_ready(inorderQueue_write_ready),
    .write_data_valid(inorderQueue_write_data_valid),
    .write_data_address(inorderQueue_write_data_address),
    .write_data_core_instruction(inorderQueue_write_data_core_instruction),
    .write_data_core_robAddr(inorderQueue_write_data_core_robAddr),
    .write_data_core_prfDest(inorderQueue_write_data_core_prfDest),
    .write_data_branch_valid(inorderQueue_write_data_branch_valid),
    .write_data_branch_mask(inorderQueue_write_data_branch_mask),
    .read_ready(inorderQueue_read_ready),
    .read_data_valid(inorderQueue_read_data_valid),
    .read_data_address(inorderQueue_read_data_address),
    .read_data_core_instruction(inorderQueue_read_data_core_instruction),
    .read_data_core_robAddr(inorderQueue_read_data_core_robAddr),
    .read_data_core_prfDest(inorderQueue_read_data_core_prfDest),
    .read_data_branch_valid(inorderQueue_read_data_branch_valid),
    .read_data_branch_mask(inorderQueue_read_data_branch_mask),
    .isEmpty(inorderQueue_isEmpty),
    .branchOps_valid(inorderQueue_branchOps_valid),
    .branchOps_branchMask(inorderQueue_branchOps_branchMask),
    .branchOps_passed(inorderQueue_branchOps_passed),
    .checkAddress(inorderQueue_checkAddress),
    .matchFound(inorderQueue_matchFound)
  );
  fifoWithBranchOps speculativeQueue ( // @[requestScheduler.scala 35:32]
    .clock(speculativeQueue_clock),
    .reset(speculativeQueue_reset),
    .write_ready(speculativeQueue_write_ready),
    .write_data_valid(speculativeQueue_write_data_valid),
    .write_data_address(speculativeQueue_write_data_address),
    .write_data_core_instruction(speculativeQueue_write_data_core_instruction),
    .write_data_core_robAddr(speculativeQueue_write_data_core_robAddr),
    .write_data_core_prfDest(speculativeQueue_write_data_core_prfDest),
    .write_data_branch_valid(speculativeQueue_write_data_branch_valid),
    .write_data_branch_mask(speculativeQueue_write_data_branch_mask),
    .write_data_writeData_valid(speculativeQueue_write_data_writeData_valid),
    .write_data_writeData_data(speculativeQueue_write_data_writeData_data),
    .write_data_cacheLine_response(speculativeQueue_write_data_cacheLine_response),
    .read_ready(speculativeQueue_read_ready),
    .read_data_valid(speculativeQueue_read_data_valid),
    .read_data_address(speculativeQueue_read_data_address),
    .read_data_core_instruction(speculativeQueue_read_data_core_instruction),
    .read_data_core_robAddr(speculativeQueue_read_data_core_robAddr),
    .read_data_core_prfDest(speculativeQueue_read_data_core_prfDest),
    .read_data_branch_valid(speculativeQueue_read_data_branch_valid),
    .read_data_branch_mask(speculativeQueue_read_data_branch_mask),
    .read_data_writeData_valid(speculativeQueue_read_data_writeData_valid),
    .read_data_writeData_data(speculativeQueue_read_data_writeData_data),
    .read_data_cacheLine_response(speculativeQueue_read_data_cacheLine_response),
    .isEmpty(speculativeQueue_isEmpty),
    .branchOps_valid(speculativeQueue_branchOps_valid),
    .branchOps_branchMask(speculativeQueue_branchOps_branchMask),
    .branchOps_passed(speculativeQueue_branchOps_passed)
  );
  assign canAllocate = inorderQueue_write_ready & speculativeQueue_write_ready; // @[requestScheduler.scala 120:43]
  assign requestOut_valid = (controlSignal_inorderReady | controlSignal_speculativeReady) & _GEN_213; // @[requestScheduler.scala 78:113 utils.scala 48:41]
  assign requestOut_address = controlSignal_inorderReady | controlSignal_speculativeReady ? _GEN_214 : 32'h0; // @[requestScheduler.scala 78:113 utils.scala 49:41]
  assign requestOut_core_instruction = controlSignal_inorderReady | controlSignal_speculativeReady ? _GEN_215 : 32'h0; // @[requestScheduler.scala 78:113 utils.scala 49:41]
  assign requestOut_core_robAddr = controlSignal_inorderReady | controlSignal_speculativeReady ? _GEN_216 : 4'h0; // @[requestScheduler.scala 78:113 utils.scala 49:41]
  assign requestOut_core_prfDest = controlSignal_inorderReady | controlSignal_speculativeReady ? _GEN_217 : 6'h0; // @[requestScheduler.scala 78:113 utils.scala 49:41]
  assign requestOut_branch_valid = (controlSignal_inorderReady | controlSignal_speculativeReady) & _GEN_218; // @[requestScheduler.scala 78:113 utils.scala 48:41]
  assign requestOut_branch_mask = controlSignal_inorderReady | controlSignal_speculativeReady ? _GEN_219 : 5'h0; // @[requestScheduler.scala 78:113 utils.scala 49:41]
  assign requestOut_writeData_valid = (controlSignal_inorderReady | controlSignal_speculativeReady) & _GEN_220; // @[requestScheduler.scala 78:113 utils.scala 48:41]
  assign requestOut_writeData_data = controlSignal_inorderReady | controlSignal_speculativeReady ? _GEN_221 : 64'h0; // @[requestScheduler.scala 78:113 utils.scala 49:41]
  assign controlSignal_isSpeculative = (controlSignal_inorderReady | controlSignal_speculativeReady) & _GEN_212; // @[requestScheduler.scala 78:113 27:31]
  assign fenceReady = inorderQueue_isEmpty & speculativeQueue_isEmpty; // @[requestScheduler.scala 121:38]
  assign inorderQueue_clock = clock;
  assign inorderQueue_reset = reset;
  assign inorderQueue_write_data_valid = requestIn_valid & _GEN_56; // @[requestScheduler.scala 50:50 62:35]
  assign inorderQueue_write_data_address = requestIn_valid ? _GEN_55 : 32'h0; // @[requestScheduler.scala 50:50 utils.scala 49:41]
  assign inorderQueue_write_data_core_instruction = requestIn_valid ? _GEN_54 : 32'h0; // @[requestScheduler.scala 50:50 utils.scala 49:41]
  assign inorderQueue_write_data_core_robAddr = requestIn_valid ? _GEN_53 : 4'h0; // @[requestScheduler.scala 50:50 utils.scala 49:41]
  assign inorderQueue_write_data_core_prfDest = requestIn_valid ? _GEN_52 : 6'h0; // @[requestScheduler.scala 50:50 utils.scala 49:41]
  assign inorderQueue_write_data_branch_valid = requestIn_valid & _GEN_51; // @[requestScheduler.scala 50:50 utils.scala 48:41]
  assign inorderQueue_write_data_branch_mask = requestIn_valid ? _GEN_50 : 5'h0; // @[requestScheduler.scala 50:50 utils.scala 49:41]
  assign inorderQueue_read_ready = (controlSignal_inorderReady | controlSignal_speculativeReady) & _GEN_225; // @[requestScheduler.scala 78:113 41:27]
  assign inorderQueue_branchOps_valid = branchOps_valid; // @[requestScheduler.scala 65:26]
  assign inorderQueue_branchOps_branchMask = branchOps_branchMask; // @[requestScheduler.scala 65:26]
  assign inorderQueue_branchOps_passed = branchOps_passed; // @[requestScheduler.scala 65:26]
  assign inorderQueue_checkAddress = requestIn_address; // @[requestScheduler.scala 40:29]
  assign speculativeQueue_clock = clock;
  assign speculativeQueue_reset = reset;
  assign speculativeQueue_write_data_valid = requestIn_valid & _GEN_68; // @[requestScheduler.scala 50:50 63:39]
  assign speculativeQueue_write_data_address = requestIn_valid ? _GEN_67 : 32'h0; // @[requestScheduler.scala 50:50 utils.scala 49:41]
  assign speculativeQueue_write_data_core_instruction = requestIn_valid ? _GEN_66 : 32'h0; // @[requestScheduler.scala 50:50 utils.scala 49:41]
  assign speculativeQueue_write_data_core_robAddr = requestIn_valid ? _GEN_65 : 4'h0; // @[requestScheduler.scala 50:50 utils.scala 49:41]
  assign speculativeQueue_write_data_core_prfDest = requestIn_valid ? _GEN_64 : 6'h0; // @[requestScheduler.scala 50:50 utils.scala 49:41]
  assign speculativeQueue_write_data_branch_valid = requestIn_valid & _GEN_63; // @[requestScheduler.scala 50:50 utils.scala 48:41]
  assign speculativeQueue_write_data_branch_mask = requestIn_valid ? _GEN_62 : 5'h0; // @[requestScheduler.scala 50:50 utils.scala 49:41]
  assign speculativeQueue_write_data_writeData_valid = 1'h0; // @[requestScheduler.scala 50:50 utils.scala 48:41]
  assign speculativeQueue_write_data_writeData_data = 64'h0; // @[requestScheduler.scala 50:50 utils.scala 49:41]
  assign speculativeQueue_write_data_cacheLine_response = 2'h0; // @[requestScheduler.scala 126:50]
  assign speculativeQueue_read_ready = (controlSignal_inorderReady | controlSignal_speculativeReady) & _GEN_211; // @[requestScheduler.scala 78:113 44:31]
  assign speculativeQueue_branchOps_valid = branchOps_valid; // @[requestScheduler.scala 66:30]
  assign speculativeQueue_branchOps_branchMask = branchOps_branchMask; // @[requestScheduler.scala 66:30]
  assign speculativeQueue_branchOps_passed = branchOps_passed; // @[requestScheduler.scala 66:30]
endmodule
module arbiter(
  input          clock,
  input          reset,
  input          request_request_valid,
  input  [31:0]  request_request_address,
  input  [31:0]  request_request_core_instruction,
  input  [3:0]   request_request_core_robAddr,
  input  [5:0]   request_request_core_prfDest,
  input          request_request_branch_valid,
  input  [4:0]   request_request_branch_mask,
  input          request_request_writeData_valid,
  input  [63:0]  request_request_writeData_data,
  input          request_isSpeculative,
  output         request_inorderReady,
  output         request_speculativeReady,
  input          toPeripheral_ready,
  output         toPeripheral_request_valid,
  output [31:0]  toPeripheral_request_address,
  output [31:0]  toPeripheral_request_core_instruction,
  output [3:0]   toPeripheral_request_core_robAddr,
  output [5:0]   toPeripheral_request_core_prfDest,
  output         toPeripheral_request_branch_valid,
  output [4:0]   toPeripheral_request_branch_mask,
  output         toPeripheral_request_writeData_valid,
  output [63:0]  toPeripheral_request_writeData_data,
  input          toCacheLookup_ready,
  input          toCacheLookup_holdInOrder,
  output [1:0]   toCacheLookup_requestType,
  output         toCacheLookup_request_valid,
  output [31:0]  toCacheLookup_request_address,
  output [31:0]  toCacheLookup_request_core_instruction,
  output [3:0]   toCacheLookup_request_core_robAddr,
  output [5:0]   toCacheLookup_request_core_prfDest,
  output         toCacheLookup_request_branch_valid,
  output [4:0]   toCacheLookup_request_branch_mask,
  output         toCacheLookup_request_writeData_valid,
  output [63:0]  toCacheLookup_request_writeData_data,
  output [511:0] toCacheLookup_request_cacheLine_cacheLine,
  output [1:0]   toCacheLookup_request_cacheLine_response,
  output         replayRequest_ready,
  input          replayRequest_request_valid,
  input  [31:0]  replayRequest_request_address,
  input  [31:0]  replayRequest_request_core_instruction,
  input  [3:0]   replayRequest_request_core_robAddr,
  input  [5:0]   replayRequest_request_core_prfDest,
  input          replayRequest_request_branch_valid,
  input  [4:0]   replayRequest_request_branch_mask,
  input          replayRequest_request_writeData_valid,
  input  [63:0]  replayRequest_request_writeData_data,
  input  [511:0] replayRequest_request_cacheLine_cacheLine,
  input  [1:0]   replayRequest_request_cacheLine_response,
  output         coherencyRequest_ready,
  input          coherencyRequest_request_valid,
  input  [31:0]  coherencyRequest_request_address,
  input  [1:0]   coherencyRequest_request_response,
  input          writeDataIn_valid,
  input  [63:0]  writeDataIn_data,
  output         writeCommit_ready,
  input          writeCommit_fired,
  input          branchOps_valid,
  input  [4:0]   branchOps_branchMask,
  input          branchOps_passed,
  input          responseOut_valid,
  input  [31:0]  responseOut_instruction,
  output         fenceReady,
  input          writeInstuctionCommitFired
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
`endif // RANDOMIZE_REG_INIT
  reg  speculativeBuffer_valid; // @[arbiter.scala 62:34]
  reg [31:0] speculativeBuffer_address; // @[arbiter.scala 62:34]
  reg [31:0] speculativeBuffer_core_instruction; // @[arbiter.scala 62:34]
  reg [3:0] speculativeBuffer_core_robAddr; // @[arbiter.scala 62:34]
  reg [5:0] speculativeBuffer_core_prfDest; // @[arbiter.scala 62:34]
  reg  speculativeBuffer_branch_valid; // @[arbiter.scala 62:34]
  reg [4:0] speculativeBuffer_branch_mask; // @[arbiter.scala 62:34]
  reg  inorderBuffer_valid; // @[arbiter.scala 63:30]
  reg [31:0] inorderBuffer_address; // @[arbiter.scala 63:30]
  reg [31:0] inorderBuffer_core_instruction; // @[arbiter.scala 63:30]
  reg [3:0] inorderBuffer_core_robAddr; // @[arbiter.scala 63:30]
  reg [5:0] inorderBuffer_core_prfDest; // @[arbiter.scala 63:30]
  reg  inorderBuffer_branch_valid; // @[arbiter.scala 63:30]
  reg [4:0] inorderBuffer_branch_mask; // @[arbiter.scala 63:30]
  reg  inorderBuffer_writeData_valid; // @[arbiter.scala 63:30]
  reg [63:0] inorderBuffer_writeData_data; // @[arbiter.scala 63:30]
  reg  operationBuffer_valid; // @[arbiter.scala 64:32]
  reg [31:0] operationBuffer_address; // @[arbiter.scala 64:32]
  reg [31:0] operationBuffer_core_instruction; // @[arbiter.scala 64:32]
  reg [3:0] operationBuffer_core_robAddr; // @[arbiter.scala 64:32]
  reg [5:0] operationBuffer_core_prfDest; // @[arbiter.scala 64:32]
  reg  operationBuffer_branch_valid; // @[arbiter.scala 64:32]
  reg [4:0] operationBuffer_branch_mask; // @[arbiter.scala 64:32]
  reg  operationBuffer_writeData_valid; // @[arbiter.scala 64:32]
  reg [63:0] operationBuffer_writeData_data; // @[arbiter.scala 64:32]
  wire  _speculativeBufferReadyWire_T = ~speculativeBuffer_valid; // @[arbiter.scala 67:48]
  wire  _operationBufferReadyWire_T = ~operationBuffer_valid; // @[arbiter.scala 68:47]
  wire  operationBufferReadyWire = ~operationBuffer_valid | operationBuffer_valid & ~operationBuffer_branch_valid; // @[arbiter.scala 68:70]
  wire  _inorderBufferReadyWire_T = ~inorderBuffer_valid; // @[arbiter.scala 69:32]
  wire  inorderBufferReadyWire = ~inorderBuffer_valid | inorderBuffer_valid & ~inorderBuffer_branch_valid; // @[arbiter.scala 69:53]
  wire  _GEN_0 = request_isSpeculative ? request_request_valid : speculativeBuffer_valid; // @[arbiter.scala 76:32 77:24 62:34]
  wire  _GEN_5 = request_isSpeculative ? request_request_branch_valid : speculativeBuffer_branch_valid; // @[arbiter.scala 76:32 77:24 62:34]
  wire [4:0] _GEN_6 = request_isSpeculative ? request_request_branch_mask : speculativeBuffer_branch_mask; // @[arbiter.scala 76:32 77:24 62:34]
  wire  _GEN_12 = request_isSpeculative ? operationBuffer_valid : request_request_valid; // @[arbiter.scala 64:32 76:32 79:23]
  wire  _GEN_17 = request_isSpeculative ? operationBuffer_branch_valid : request_request_branch_valid; // @[arbiter.scala 64:32 76:32 79:23]
  wire [4:0] _GEN_18 = request_isSpeculative ? operationBuffer_branch_mask : request_request_branch_mask; // @[arbiter.scala 64:32 76:32 79:23]
  wire  _GEN_24 = request_request_valid & request_request_branch_valid ? _GEN_0 : speculativeBuffer_valid; // @[arbiter.scala 62:34 75:62]
  wire  _GEN_29 = request_request_valid & request_request_branch_valid ? _GEN_5 : speculativeBuffer_branch_valid; // @[arbiter.scala 62:34 75:62]
  wire [4:0] _GEN_30 = request_request_valid & request_request_branch_valid ? _GEN_6 : speculativeBuffer_branch_mask; // @[arbiter.scala 62:34 75:62]
  wire  _GEN_36 = request_request_valid & request_request_branch_valid ? _GEN_12 : operationBuffer_valid; // @[arbiter.scala 64:32 75:62]
  wire  _GEN_41 = request_request_valid & request_request_branch_valid ? _GEN_17 : operationBuffer_branch_valid; // @[arbiter.scala 64:32 75:62]
  wire [4:0] _GEN_42 = request_request_valid & request_request_branch_valid ? _GEN_18 : operationBuffer_branch_mask; // @[arbiter.scala 64:32 75:62]
  reg [2:0] operationState; // @[arbiter.scala 85:31]
  wire  operationWires_isRead = operationBuffer_core_instruction[6:0] == 7'h3; // @[arbiter.scala 99:66]
  wire  operationWires_isWrite = operationBuffer_core_instruction[6:0] == 7'h23; // @[arbiter.scala 100:67]
  wire  operationWires_rAtomics = operationBuffer_core_instruction[6:0] == 7'h2f; // @[arbiter.scala 101:68]
  wire  operationWires_isLR = operationBuffer_core_instruction[31:27] == 5'h2 & operationWires_rAtomics; // @[arbiter.scala 102:81]
  wire  operationWires_isSC = operationBuffer_core_instruction[31:27] == 5'h3 & operationWires_rAtomics; // @[arbiter.scala 103:81]
  wire  operationWires_isPeriRead = operationWires_isRead & operationBuffer_address == 32'h40600000; // @[arbiter.scala 104:87]
  wire  operationWires_isPeriWrite = operationWires_isWrite & operationBuffer_address == 32'h40600004; // @[arbiter.scala 105:88]
  wire  _GEN_48 = operationWires_isLR | operationWires_isSC | operationWires_rAtomics ? operationBuffer_valid :
    inorderBuffer_valid; // @[arbiter.scala 118:91 120:25 63:30]
  wire [31:0] _GEN_49 = operationWires_isLR | operationWires_isSC | operationWires_rAtomics ? operationBuffer_address :
    inorderBuffer_address; // @[arbiter.scala 118:91 120:25 63:30]
  wire [31:0] _GEN_50 = operationWires_isLR | operationWires_isSC | operationWires_rAtomics ?
    operationBuffer_core_instruction : inorderBuffer_core_instruction; // @[arbiter.scala 118:91 120:25 63:30]
  wire [3:0] _GEN_51 = operationWires_isLR | operationWires_isSC | operationWires_rAtomics ?
    operationBuffer_core_robAddr : inorderBuffer_core_robAddr; // @[arbiter.scala 118:91 120:25 63:30]
  wire [5:0] _GEN_52 = operationWires_isLR | operationWires_isSC | operationWires_rAtomics ?
    operationBuffer_core_prfDest : inorderBuffer_core_prfDest; // @[arbiter.scala 118:91 120:25 63:30]
  wire  _GEN_53 = operationWires_isLR | operationWires_isSC | operationWires_rAtomics ? operationBuffer_branch_valid :
    inorderBuffer_branch_valid; // @[arbiter.scala 118:91 120:25 63:30]
  wire [4:0] _GEN_54 = operationWires_isLR | operationWires_isSC | operationWires_rAtomics ? operationBuffer_branch_mask
     : inorderBuffer_branch_mask; // @[arbiter.scala 118:91 120:25 63:30]
  wire  _GEN_55 = operationWires_isLR | operationWires_isSC | operationWires_rAtomics ? 1'h0 :
    inorderBuffer_writeData_valid; // @[arbiter.scala 118:91 121:41 63:30]
  wire [63:0] _GEN_56 = operationWires_isLR | operationWires_isSC | operationWires_rAtomics ?
    operationBuffer_writeData_data : inorderBuffer_writeData_data; // @[arbiter.scala 118:91 120:25 63:30]
  wire [2:0] _GEN_60 = operationWires_isLR | operationWires_isSC | operationWires_rAtomics ? 3'h3 : operationState; // @[arbiter.scala 118:91 122:26 85:31]
  wire  _GEN_61 = (operationWires_isLR | operationWires_isSC | operationWires_rAtomics) & _GEN_36; // @[arbiter.scala 118:91 125:33]
  wire [2:0] _GEN_62 = operationWires_isWrite ? 3'h1 : _GEN_60; // @[arbiter.scala 115:44 117:26]
  wire  _GEN_63 = operationWires_isWrite ? inorderBuffer_valid : _GEN_48; // @[arbiter.scala 115:44 63:30]
  wire [31:0] _GEN_64 = operationWires_isWrite ? inorderBuffer_address : _GEN_49; // @[arbiter.scala 115:44 63:30]
  wire [31:0] _GEN_65 = operationWires_isWrite ? inorderBuffer_core_instruction : _GEN_50; // @[arbiter.scala 115:44 63:30]
  wire [3:0] _GEN_66 = operationWires_isWrite ? inorderBuffer_core_robAddr : _GEN_51; // @[arbiter.scala 115:44 63:30]
  wire [5:0] _GEN_67 = operationWires_isWrite ? inorderBuffer_core_prfDest : _GEN_52; // @[arbiter.scala 115:44 63:30]
  wire  _GEN_68 = operationWires_isWrite ? inorderBuffer_branch_valid : _GEN_53; // @[arbiter.scala 115:44 63:30]
  wire [4:0] _GEN_69 = operationWires_isWrite ? inorderBuffer_branch_mask : _GEN_54; // @[arbiter.scala 115:44 63:30]
  wire  _GEN_70 = operationWires_isWrite ? inorderBuffer_writeData_valid : _GEN_55; // @[arbiter.scala 115:44 63:30]
  wire [63:0] _GEN_71 = operationWires_isWrite ? inorderBuffer_writeData_data : _GEN_56; // @[arbiter.scala 115:44 63:30]
  wire  _GEN_75 = operationWires_isWrite ? _GEN_36 : _GEN_61; // @[arbiter.scala 115:44]
  wire  _GEN_76 = operationWires_isRead ? operationBuffer_valid : _GEN_63; // @[arbiter.scala 111:36 113:25]
  wire  _GEN_81 = operationWires_isRead ? operationBuffer_branch_valid : _GEN_68; // @[arbiter.scala 111:36 113:25]
  wire [4:0] _GEN_82 = operationWires_isRead ? operationBuffer_branch_mask : _GEN_69; // @[arbiter.scala 111:36 113:25]
  wire  _GEN_90 = operationBuffer_valid ? _GEN_76 : inorderBuffer_valid; // @[arbiter.scala 110:33 63:30]
  wire  _GEN_95 = operationBuffer_valid ? _GEN_81 : inorderBuffer_branch_valid; // @[arbiter.scala 110:33 63:30]
  wire [4:0] _GEN_96 = operationBuffer_valid ? _GEN_82 : inorderBuffer_branch_mask; // @[arbiter.scala 110:33 63:30]
  wire  _GEN_104 = writeDataIn_valid ? operationBuffer_valid : inorderBuffer_valid; // @[arbiter.scala 135:30 137:23 63:30]
  wire [31:0] _GEN_105 = writeDataIn_valid ? operationBuffer_address : inorderBuffer_address; // @[arbiter.scala 135:30 137:23 63:30]
  wire [31:0] _GEN_106 = writeDataIn_valid ? operationBuffer_core_instruction : inorderBuffer_core_instruction; // @[arbiter.scala 135:30 137:23 63:30]
  wire [3:0] _GEN_107 = writeDataIn_valid ? operationBuffer_core_robAddr : inorderBuffer_core_robAddr; // @[arbiter.scala 135:30 137:23 63:30]
  wire [5:0] _GEN_108 = writeDataIn_valid ? operationBuffer_core_prfDest : inorderBuffer_core_prfDest; // @[arbiter.scala 135:30 137:23 63:30]
  wire  _GEN_109 = writeDataIn_valid ? operationBuffer_branch_valid : inorderBuffer_branch_valid; // @[arbiter.scala 135:30 137:23 63:30]
  wire [4:0] _GEN_110 = writeDataIn_valid ? operationBuffer_branch_mask : inorderBuffer_branch_mask; // @[arbiter.scala 135:30 137:23 63:30]
  wire  _GEN_111 = writeDataIn_valid ? writeDataIn_valid : inorderBuffer_writeData_valid; // @[arbiter.scala 135:30 139:39 63:30]
  wire [63:0] _GEN_112 = writeDataIn_valid ? writeDataIn_data : inorderBuffer_writeData_data; // @[arbiter.scala 135:30 138:38 63:30]
  wire  _GEN_116 = writeDataIn_valid ? 1'h0 : _GEN_36; // @[arbiter.scala 135:30 140:31]
  wire [2:0] _GEN_117 = writeDataIn_valid ? 3'h4 : operationState; // @[arbiter.scala 135:30 141:24 85:31]
  wire [2:0] _operationState_T_3 = responseOut_valid & responseOut_instruction == operationBuffer_core_instruction ? 3'h1
     : 3'h3; // @[arbiter.scala 145:28]
  wire [2:0] _operationState_T_4 = writeInstuctionCommitFired ? 3'h0 : 3'h4; // @[arbiter.scala 149:28]
  wire [2:0] _GEN_118 = 3'h4 == operationState ? _operationState_T_4 : operationState; // @[arbiter.scala 107:25 149:22 85:31]
  wire [2:0] _GEN_119 = 3'h3 == operationState ? _operationState_T_3 : _GEN_118; // @[arbiter.scala 107:25 145:22]
  wire  _GEN_120 = 3'h2 == operationState ? _GEN_104 : inorderBuffer_valid; // @[arbiter.scala 107:25 63:30]
  wire  _GEN_125 = 3'h2 == operationState ? _GEN_109 : inorderBuffer_branch_valid; // @[arbiter.scala 107:25 63:30]
  wire [4:0] _GEN_126 = 3'h2 == operationState ? _GEN_110 : inorderBuffer_branch_mask; // @[arbiter.scala 107:25 63:30]
  wire  _GEN_136 = 3'h1 == operationState ? inorderBuffer_valid : _GEN_120; // @[arbiter.scala 107:25 63:30]
  wire  _GEN_141 = 3'h1 == operationState ? inorderBuffer_branch_valid : _GEN_125; // @[arbiter.scala 107:25 63:30]
  wire [4:0] _GEN_142 = 3'h1 == operationState ? inorderBuffer_branch_mask : _GEN_126; // @[arbiter.scala 107:25 63:30]
  wire  _GEN_150 = 3'h0 == operationState ? _GEN_90 : _GEN_136; // @[arbiter.scala 107:25]
  wire  _GEN_155 = 3'h0 == operationState ? _GEN_95 : _GEN_141; // @[arbiter.scala 107:25]
  wire [4:0] _GEN_156 = 3'h0 == operationState ? _GEN_96 : _GEN_142; // @[arbiter.scala 107:25]
  reg  atomicBusyState; // @[arbiter.scala 175:32]
  wire  _T_24 = ~toCacheLookup_holdInOrder; // @[arbiter.scala 178:29]
  wire  _T_26 = operationWires_isPeriRead | operationWires_isPeriWrite; // @[arbiter.scala 179:63]
  wire  _T_27 = ~(operationWires_isPeriRead | operationWires_isPeriWrite); // @[arbiter.scala 179:35]
  wire [1:0] _GEN_224 = inorderBuffer_valid & ~(operationWires_isPeriRead | operationWires_isPeriWrite) ? 2'h1 : 2'h0; // @[arbiter.scala 179:94 183:25]
  wire  _GEN_267 = inorderBuffer_valid & _T_24 & _T_27 | speculativeBuffer_valid; // @[arbiter.scala 201:130 205:23]
  wire [1:0] _GEN_283 = replayRequest_request_valid ? 2'h2 : {{1'd0}, _GEN_267}; // @[arbiter.scala 196:44 199:23]
  wire [1:0] _GEN_292 = coherencyRequest_request_valid ? 2'h3 : _GEN_283; // @[arbiter.scala 188:47 195:23]
  wire [1:0] _GEN_318 = atomicBusyState & ~toCacheLookup_holdInOrder ? _GEN_224 : _GEN_292; // @[arbiter.scala 178:56]
  wire [1:0] requestTypeWire = toCacheLookup_ready ? _GEN_318 : 2'h0; // @[arbiter.scala 177:72]
  wire [4:0] _T_9 = speculativeBuffer_branch_mask & branchOps_branchMask; // @[utils.scala 122:29]
  wire  _T_10 = |_T_9; // @[utils.scala 122:53]
  wire [4:0] _speculativeBuffer_branch_mask_T = speculativeBuffer_branch_mask ^ branchOps_branchMask; // @[utils.scala 123:40]
  wire [4:0] _GEN_165 = |_T_9 ? _speculativeBuffer_branch_mask_T : _GEN_30; // @[utils.scala 122:58 123:25]
  wire  _GEN_166 = _T_10 ? 1'h0 : _GEN_29; // @[utils.scala 127:58 128:26]
  wire [4:0] _GEN_167 = _T_10 ? 5'h0 : _GEN_30; // @[utils.scala 127:58 129:25]
  wire [4:0] _GEN_168 = branchOps_passed ? _GEN_165 : _GEN_167; // @[utils.scala 121:32]
  wire  _GEN_169 = branchOps_passed ? speculativeBuffer_branch_valid : _GEN_166; // @[utils.scala 121:32 125:24]
  wire [4:0] _GEN_170 = branchOps_valid ? _GEN_168 : _GEN_30; // @[utils.scala 120:29]
  wire  _GEN_171 = branchOps_valid ? _GEN_169 : _GEN_29; // @[utils.scala 120:29]
  wire [4:0] _T_13 = operationBuffer_branch_mask & branchOps_branchMask; // @[utils.scala 122:29]
  wire  _T_14 = |_T_13; // @[utils.scala 122:53]
  wire [4:0] _operationBuffer_branch_mask_T = operationBuffer_branch_mask ^ branchOps_branchMask; // @[utils.scala 123:40]
  wire [4:0] _GEN_176 = |_T_13 ? _operationBuffer_branch_mask_T : _GEN_42; // @[utils.scala 122:58 123:25]
  wire  _GEN_177 = _T_14 ? 1'h0 : _GEN_41; // @[utils.scala 127:58 128:26]
  wire [4:0] _GEN_178 = _T_14 ? 5'h0 : _GEN_42; // @[utils.scala 127:58 129:25]
  wire [4:0] _GEN_179 = branchOps_passed ? _GEN_176 : _GEN_178; // @[utils.scala 121:32]
  wire  _GEN_180 = branchOps_passed ? operationBuffer_branch_valid : _GEN_177; // @[utils.scala 121:32 125:24]
  wire [4:0] _GEN_181 = branchOps_valid ? _GEN_179 : _GEN_42; // @[utils.scala 120:29]
  wire  _GEN_182 = branchOps_valid ? _GEN_180 : _GEN_41; // @[utils.scala 120:29]
  wire [4:0] _T_17 = inorderBuffer_branch_mask & branchOps_branchMask; // @[utils.scala 122:29]
  wire  _T_18 = |_T_17; // @[utils.scala 122:53]
  wire [4:0] _inorderBuffer_branch_mask_T = inorderBuffer_branch_mask ^ branchOps_branchMask; // @[utils.scala 123:40]
  wire [4:0] _GEN_187 = |_T_17 ? _inorderBuffer_branch_mask_T : _GEN_156; // @[utils.scala 122:58 123:25]
  wire  _GEN_188 = _T_18 ? 1'h0 : _GEN_155; // @[utils.scala 127:58 128:26]
  wire [4:0] _GEN_189 = _T_18 ? 5'h0 : _GEN_156; // @[utils.scala 127:58 129:25]
  wire [4:0] _GEN_190 = branchOps_passed ? _GEN_187 : _GEN_189; // @[utils.scala 121:32]
  wire  _GEN_191 = branchOps_passed ? inorderBuffer_branch_valid : _GEN_188; // @[utils.scala 121:32 125:24]
  wire [4:0] _GEN_192 = branchOps_valid ? _GEN_190 : _GEN_156; // @[utils.scala 120:29]
  wire  _GEN_193 = branchOps_valid ? _GEN_191 : _GEN_155; // @[utils.scala 120:29]
  wire [4:0] _GEN_204 = _T_18 ? _inorderBuffer_branch_mask_T : inorderBuffer_branch_mask; // @[utils.scala 92:56 93:27 96:27]
  wire [4:0] _GEN_205 = _T_18 ? 5'h0 : inorderBuffer_branch_mask; // @[utils.scala 101:56 102:27 106:27]
  wire  _GEN_206 = _T_18 ? 1'h0 : inorderBuffer_branch_valid; // @[utils.scala 101:56 103:28 107:28]
  wire [4:0] _GEN_207 = branchOps_passed ? _GEN_204 : _GEN_205; // @[utils.scala 90:30]
  wire  _GEN_208 = branchOps_passed ? inorderBuffer_branch_valid : _GEN_206; // @[utils.scala 90:30 98:26]
  wire [4:0] _GEN_209 = branchOps_valid ? _GEN_207 : inorderBuffer_branch_mask; // @[utils.scala 111:23 89:27]
  wire  _GEN_210 = branchOps_valid ? _GEN_208 : inorderBuffer_branch_valid; // @[utils.scala 112:24 89:27]
  wire  _GEN_211 = inorderBuffer_valid & ~(operationWires_isPeriRead | operationWires_isPeriWrite) ? 1'h0 : _GEN_150; // @[arbiter.scala 179:94 180:29]
  wire  _GEN_212 = inorderBuffer_valid & ~(operationWires_isPeriRead | operationWires_isPeriWrite) & inorderBuffer_valid
    ; // @[arbiter.scala 179:94 182:31 utils.scala 48:41]
  wire [31:0] _GEN_213 = inorderBuffer_valid & ~(operationWires_isPeriRead | operationWires_isPeriWrite) ?
    inorderBuffer_address : 32'h0; // @[arbiter.scala 179:94 182:31 utils.scala 49:41]
  wire [31:0] _GEN_214 = inorderBuffer_valid & ~(operationWires_isPeriRead | operationWires_isPeriWrite) ?
    inorderBuffer_core_instruction : 32'h0; // @[arbiter.scala 179:94 182:31 utils.scala 49:41]
  wire [3:0] _GEN_215 = inorderBuffer_valid & ~(operationWires_isPeriRead | operationWires_isPeriWrite) ?
    inorderBuffer_core_robAddr : 4'h0; // @[arbiter.scala 179:94 182:31 utils.scala 49:41]
  wire [5:0] _GEN_216 = inorderBuffer_valid & ~(operationWires_isPeriRead | operationWires_isPeriWrite) ?
    inorderBuffer_core_prfDest : 6'h0; // @[arbiter.scala 179:94 182:31 utils.scala 49:41]
  wire  _GEN_217 = inorderBuffer_valid & ~(operationWires_isPeriRead | operationWires_isPeriWrite) & _GEN_210; // @[arbiter.scala 179:94 utils.scala 48:41]
  wire [4:0] _GEN_218 = inorderBuffer_valid & ~(operationWires_isPeriRead | operationWires_isPeriWrite) ? _GEN_209 : 5'h0
    ; // @[arbiter.scala 179:94 utils.scala 49:41]
  wire  _GEN_219 = inorderBuffer_valid & ~(operationWires_isPeriRead | operationWires_isPeriWrite) &
    inorderBuffer_writeData_valid; // @[arbiter.scala 179:94 182:31 utils.scala 48:41]
  wire [63:0] _GEN_220 = inorderBuffer_valid & ~(operationWires_isPeriRead | operationWires_isPeriWrite) ?
    inorderBuffer_writeData_data : 64'h0; // @[arbiter.scala 179:94 182:31 utils.scala 49:41]
  wire [4:0] _GEN_233 = _T_10 ? _speculativeBuffer_branch_mask_T : speculativeBuffer_branch_mask; // @[utils.scala 92:56 93:27 96:27]
  wire [4:0] _GEN_234 = _T_10 ? 5'h0 : speculativeBuffer_branch_mask; // @[utils.scala 101:56 102:27 106:27]
  wire  _GEN_235 = _T_10 ? 1'h0 : speculativeBuffer_branch_valid; // @[utils.scala 101:56 103:28 107:28]
  wire [4:0] _GEN_236 = branchOps_passed ? _GEN_233 : _GEN_234; // @[utils.scala 90:30]
  wire  _GEN_237 = branchOps_passed ? speculativeBuffer_branch_valid : _GEN_235; // @[utils.scala 90:30 98:26]
  wire [4:0] _GEN_238 = branchOps_valid ? _GEN_236 : speculativeBuffer_branch_mask; // @[utils.scala 111:23 89:27]
  wire  _GEN_239 = branchOps_valid ? _GEN_237 : speculativeBuffer_branch_valid; // @[utils.scala 112:24 89:27]
  wire  _GEN_240 = speculativeBuffer_valid ? 1'h0 : _GEN_24; // @[arbiter.scala 210:42 211:31]
  wire [31:0] _GEN_242 = speculativeBuffer_valid ? speculativeBuffer_address : 32'h0; // @[arbiter.scala 210:42 213:29 utils.scala 49:41]
  wire [31:0] _GEN_243 = speculativeBuffer_valid ? speculativeBuffer_core_instruction : 32'h0; // @[arbiter.scala 210:42 213:29 utils.scala 49:41]
  wire [3:0] _GEN_244 = speculativeBuffer_valid ? speculativeBuffer_core_robAddr : 4'h0; // @[arbiter.scala 210:42 213:29 utils.scala 49:41]
  wire [5:0] _GEN_245 = speculativeBuffer_valid ? speculativeBuffer_core_prfDest : 6'h0; // @[arbiter.scala 210:42 213:29 utils.scala 49:41]
  wire  _GEN_246 = speculativeBuffer_valid & _GEN_239; // @[arbiter.scala 210:42 utils.scala 48:41]
  wire [4:0] _GEN_247 = speculativeBuffer_valid ? _GEN_238 : 5'h0; // @[arbiter.scala 210:42 utils.scala 49:41]
  wire  _GEN_254 = inorderBuffer_valid & _T_24 & _T_27 ? 1'h0 : _GEN_150; // @[arbiter.scala 201:130 202:27]
  wire  _GEN_255 = inorderBuffer_valid & _T_24 & _T_27 ? inorderBuffer_valid : speculativeBuffer_valid; // @[arbiter.scala 201:130 204:29]
  wire [31:0] _GEN_256 = inorderBuffer_valid & _T_24 & _T_27 ? inorderBuffer_address : _GEN_242; // @[arbiter.scala 201:130 204:29]
  wire [31:0] _GEN_257 = inorderBuffer_valid & _T_24 & _T_27 ? inorderBuffer_core_instruction : _GEN_243; // @[arbiter.scala 201:130 204:29]
  wire [3:0] _GEN_258 = inorderBuffer_valid & _T_24 & _T_27 ? inorderBuffer_core_robAddr : _GEN_244; // @[arbiter.scala 201:130 204:29]
  wire [5:0] _GEN_259 = inorderBuffer_valid & _T_24 & _T_27 ? inorderBuffer_core_prfDest : _GEN_245; // @[arbiter.scala 201:130 204:29]
  wire  _GEN_260 = inorderBuffer_valid & _T_24 & _T_27 ? _GEN_210 : _GEN_246; // @[arbiter.scala 201:130]
  wire [4:0] _GEN_261 = inorderBuffer_valid & _T_24 & _T_27 ? _GEN_209 : _GEN_247; // @[arbiter.scala 201:130]
  wire  _GEN_262 = inorderBuffer_valid & _T_24 & _T_27 & inorderBuffer_writeData_valid; // @[arbiter.scala 201:130 204:29]
  wire [63:0] _GEN_263 = inorderBuffer_valid & _T_24 & _T_27 ? inorderBuffer_writeData_data : 64'h0; // @[arbiter.scala 201:130 204:29]
  wire  _GEN_268 = inorderBuffer_valid & _T_24 & _T_27 ? operationWires_rAtomics & ~inorderBuffer_writeData_valid :
    atomicBusyState; // @[arbiter.scala 201:130 208:23 175:32]
  wire  _GEN_269 = inorderBuffer_valid & _T_24 & _T_27 ? _GEN_24 : _GEN_240; // @[arbiter.scala 201:130]
  wire  _GEN_271 = replayRequest_request_valid ? replayRequest_request_valid : _GEN_255; // @[arbiter.scala 196:44 198:29]
  wire [31:0] _GEN_272 = replayRequest_request_valid ? replayRequest_request_address : _GEN_256; // @[arbiter.scala 196:44 198:29]
  wire [31:0] _GEN_273 = replayRequest_request_valid ? replayRequest_request_core_instruction : _GEN_257; // @[arbiter.scala 196:44 198:29]
  wire [3:0] _GEN_274 = replayRequest_request_valid ? replayRequest_request_core_robAddr : _GEN_258; // @[arbiter.scala 196:44 198:29]
  wire [5:0] _GEN_275 = replayRequest_request_valid ? replayRequest_request_core_prfDest : _GEN_259; // @[arbiter.scala 196:44 198:29]
  wire  _GEN_276 = replayRequest_request_valid ? replayRequest_request_branch_valid : _GEN_260; // @[arbiter.scala 196:44 198:29]
  wire [4:0] _GEN_277 = replayRequest_request_valid ? replayRequest_request_branch_mask : _GEN_261; // @[arbiter.scala 196:44 198:29]
  wire  _GEN_278 = replayRequest_request_valid ? replayRequest_request_writeData_valid : _GEN_262; // @[arbiter.scala 196:44 198:29]
  wire [63:0] _GEN_279 = replayRequest_request_valid ? replayRequest_request_writeData_data : _GEN_263; // @[arbiter.scala 196:44 198:29]
  wire [511:0] _GEN_280 = replayRequest_request_valid ? replayRequest_request_cacheLine_cacheLine : 512'h0; // @[arbiter.scala 196:44 198:29]
  wire [1:0] _GEN_281 = replayRequest_request_valid ? replayRequest_request_cacheLine_response : 2'h0; // @[arbiter.scala 196:44 198:29]
  wire  _GEN_284 = replayRequest_request_valid ? _GEN_150 : _GEN_254; // @[arbiter.scala 196:44]
  wire  _GEN_285 = replayRequest_request_valid ? atomicBusyState : _GEN_268; // @[arbiter.scala 175:32 196:44]
  wire  _GEN_286 = replayRequest_request_valid ? _GEN_24 : _GEN_269; // @[arbiter.scala 196:44]
  wire  _GEN_288 = coherencyRequest_request_valid ? coherencyRequest_request_valid : _GEN_271; // @[arbiter.scala 188:47 191:35]
  wire [31:0] _GEN_289 = coherencyRequest_request_valid ? coherencyRequest_request_address : _GEN_272; // @[arbiter.scala 188:47 192:37]
  wire [1:0] _GEN_290 = coherencyRequest_request_valid ? coherencyRequest_request_response : _GEN_281; // @[arbiter.scala 188:47 193:48]
  wire  _GEN_291 = coherencyRequest_request_valid | _GEN_276; // @[arbiter.scala 188:47 194:42]
  wire  _GEN_293 = coherencyRequest_request_valid ? 1'h0 : replayRequest_request_valid; // @[arbiter.scala 188:47 57:23]
  wire [31:0] _GEN_294 = coherencyRequest_request_valid ? 32'h0 : _GEN_273; // @[arbiter.scala 188:47 utils.scala 49:41]
  wire [3:0] _GEN_295 = coherencyRequest_request_valid ? 4'h0 : _GEN_274; // @[arbiter.scala 188:47 utils.scala 49:41]
  wire [5:0] _GEN_296 = coherencyRequest_request_valid ? 6'h0 : _GEN_275; // @[arbiter.scala 188:47 utils.scala 49:41]
  wire [4:0] _GEN_297 = coherencyRequest_request_valid ? 5'h0 : _GEN_277; // @[arbiter.scala 188:47 utils.scala 49:41]
  wire  _GEN_298 = coherencyRequest_request_valid ? 1'h0 : _GEN_278; // @[arbiter.scala 188:47 utils.scala 48:41]
  wire [63:0] _GEN_299 = coherencyRequest_request_valid ? 64'h0 : _GEN_279; // @[arbiter.scala 188:47 utils.scala 49:41]
  wire [511:0] _GEN_300 = coherencyRequest_request_valid ? 512'h0 : _GEN_280; // @[arbiter.scala 188:47 utils.scala 49:41]
  wire  _GEN_302 = coherencyRequest_request_valid ? _GEN_150 : _GEN_284; // @[arbiter.scala 188:47]
  wire  _GEN_306 = atomicBusyState & ~toCacheLookup_holdInOrder ? _GEN_212 : _GEN_288; // @[arbiter.scala 178:56]
  wire [31:0] _GEN_307 = atomicBusyState & ~toCacheLookup_holdInOrder ? _GEN_213 : _GEN_289; // @[arbiter.scala 178:56]
  wire [31:0] _GEN_308 = atomicBusyState & ~toCacheLookup_holdInOrder ? _GEN_214 : _GEN_294; // @[arbiter.scala 178:56]
  wire [3:0] _GEN_309 = atomicBusyState & ~toCacheLookup_holdInOrder ? _GEN_215 : _GEN_295; // @[arbiter.scala 178:56]
  wire [5:0] _GEN_310 = atomicBusyState & ~toCacheLookup_holdInOrder ? _GEN_216 : _GEN_296; // @[arbiter.scala 178:56]
  wire  _GEN_311 = atomicBusyState & ~toCacheLookup_holdInOrder ? _GEN_217 : _GEN_291; // @[arbiter.scala 178:56]
  wire [4:0] _GEN_312 = atomicBusyState & ~toCacheLookup_holdInOrder ? _GEN_218 : _GEN_297; // @[arbiter.scala 178:56]
  wire  _GEN_313 = atomicBusyState & ~toCacheLookup_holdInOrder ? _GEN_219 : _GEN_298; // @[arbiter.scala 178:56]
  wire [63:0] _GEN_314 = atomicBusyState & ~toCacheLookup_holdInOrder ? _GEN_220 : _GEN_299; // @[arbiter.scala 178:56]
  wire [511:0] _GEN_315 = atomicBusyState & ~toCacheLookup_holdInOrder ? 512'h0 : _GEN_300; // @[arbiter.scala 178:56]
  wire [1:0] _GEN_316 = atomicBusyState & ~toCacheLookup_holdInOrder ? 2'h0 : _GEN_290; // @[arbiter.scala 178:56]
  wire  _GEN_320 = atomicBusyState & ~toCacheLookup_holdInOrder ? 1'h0 : coherencyRequest_request_valid; // @[arbiter.scala 178:56 58:26]
  wire  _GEN_321 = atomicBusyState & ~toCacheLookup_holdInOrder ? 1'h0 : _GEN_293; // @[arbiter.scala 178:56 57:23]
  wire  _GEN_329 = toCacheLookup_ready & _GEN_311; // @[arbiter.scala 177:72 utils.scala 48:41]
  wire [4:0] _GEN_330 = toCacheLookup_ready ? _GEN_312 : 5'h0; // @[arbiter.scala 177:72 utils.scala 49:41]
  assign request_inorderReady = inorderBufferReadyWire & operationBufferReadyWire; // @[arbiter.scala 72:51]
  assign request_speculativeReady = ~speculativeBuffer_valid | speculativeBuffer_valid & ~speculativeBuffer_branch_valid
    ; // @[arbiter.scala 67:73]
  assign toPeripheral_request_valid = toPeripheral_ready & _T_26 & inorderBuffer_valid & inorderBuffer_valid; // @[arbiter.scala 223:112 225:26 utils.scala 48:41]
  assign toPeripheral_request_address = toPeripheral_ready & _T_26 & inorderBuffer_valid ? inorderBuffer_address : 32'h0
    ; // @[arbiter.scala 223:112 225:26 utils.scala 49:41]
  assign toPeripheral_request_core_instruction = toPeripheral_ready & _T_26 & inorderBuffer_valid ?
    inorderBuffer_core_instruction : 32'h0; // @[arbiter.scala 223:112 225:26 utils.scala 49:41]
  assign toPeripheral_request_core_robAddr = toPeripheral_ready & _T_26 & inorderBuffer_valid ?
    inorderBuffer_core_robAddr : 4'h0; // @[arbiter.scala 223:112 225:26 utils.scala 49:41]
  assign toPeripheral_request_core_prfDest = toPeripheral_ready & _T_26 & inorderBuffer_valid ?
    inorderBuffer_core_prfDest : 6'h0; // @[arbiter.scala 223:112 225:26 utils.scala 49:41]
  assign toPeripheral_request_branch_valid = toPeripheral_ready & _T_26 & inorderBuffer_valid &
    inorderBuffer_branch_valid; // @[arbiter.scala 223:112 225:26 utils.scala 48:41]
  assign toPeripheral_request_branch_mask = toPeripheral_ready & _T_26 & inorderBuffer_valid ? inorderBuffer_branch_mask
     : 5'h0; // @[arbiter.scala 223:112 225:26 utils.scala 49:41]
  assign toPeripheral_request_writeData_valid = toPeripheral_ready & _T_26 & inorderBuffer_valid &
    inorderBuffer_writeData_valid; // @[arbiter.scala 223:112 225:26 utils.scala 48:41]
  assign toPeripheral_request_writeData_data = toPeripheral_ready & _T_26 & inorderBuffer_valid ?
    inorderBuffer_writeData_data : 64'h0; // @[arbiter.scala 223:112 225:26 utils.scala 49:41]
  assign toCacheLookup_requestType = toCacheLookup_ready ? requestTypeWire : 2'h0; // @[arbiter.scala 177:72 221:31 56:29]
  assign toCacheLookup_request_valid = toCacheLookup_ready & _GEN_306; // @[arbiter.scala 177:72 utils.scala 48:41]
  assign toCacheLookup_request_address = toCacheLookup_ready ? _GEN_307 : 32'h0; // @[arbiter.scala 177:72 utils.scala 49:41]
  assign toCacheLookup_request_core_instruction = toCacheLookup_ready ? _GEN_308 : 32'h0; // @[arbiter.scala 177:72 utils.scala 49:41]
  assign toCacheLookup_request_core_robAddr = toCacheLookup_ready ? _GEN_309 : 4'h0; // @[arbiter.scala 177:72 utils.scala 49:41]
  assign toCacheLookup_request_core_prfDest = toCacheLookup_ready ? _GEN_310 : 6'h0; // @[arbiter.scala 177:72 utils.scala 49:41]
  assign toCacheLookup_request_branch_valid = toPeripheral_ready & _T_26 & inorderBuffer_valid ? _GEN_210 : _GEN_329; // @[arbiter.scala 223:112]
  assign toCacheLookup_request_branch_mask = toPeripheral_ready & _T_26 & inorderBuffer_valid ? _GEN_209 : _GEN_330; // @[arbiter.scala 223:112]
  assign toCacheLookup_request_writeData_valid = toCacheLookup_ready & _GEN_313; // @[arbiter.scala 177:72 utils.scala 48:41]
  assign toCacheLookup_request_writeData_data = toCacheLookup_ready ? _GEN_314 : 64'h0; // @[arbiter.scala 177:72 utils.scala 49:41]
  assign toCacheLookup_request_cacheLine_cacheLine = toCacheLookup_ready ? _GEN_315 : 512'h0; // @[arbiter.scala 177:72 utils.scala 49:41]
  assign toCacheLookup_request_cacheLine_response = toCacheLookup_ready ? _GEN_316 : 2'h0; // @[arbiter.scala 177:72 utils.scala 49:41]
  assign replayRequest_ready = toCacheLookup_ready & _GEN_321; // @[arbiter.scala 177:72 57:23]
  assign coherencyRequest_ready = toCacheLookup_ready & _GEN_320; // @[arbiter.scala 177:72 58:26]
  assign writeCommit_ready = 3'h0 == operationState ? 1'h0 : 3'h1 == operationState; // @[arbiter.scala 107:25 59:21]
  assign fenceReady = _speculativeBufferReadyWire_T & _inorderBufferReadyWire_T & _operationBufferReadyWire_T; // @[arbiter.scala 230:67]
  always @(posedge clock) begin
    if (reset) begin // @[arbiter.scala 62:34]
      speculativeBuffer_valid <= 1'h0; // @[arbiter.scala 62:34]
    end else if (toCacheLookup_ready) begin // @[arbiter.scala 177:72]
      if (atomicBusyState & ~toCacheLookup_holdInOrder) begin // @[arbiter.scala 178:56]
        speculativeBuffer_valid <= _GEN_24;
      end else if (coherencyRequest_request_valid) begin // @[arbiter.scala 188:47]
        speculativeBuffer_valid <= _GEN_24;
      end else begin
        speculativeBuffer_valid <= _GEN_286;
      end
    end else begin
      speculativeBuffer_valid <= _GEN_24;
    end
    if (reset) begin // @[arbiter.scala 62:34]
      speculativeBuffer_address <= 32'h0; // @[arbiter.scala 62:34]
    end else if (request_request_valid & request_request_branch_valid) begin // @[arbiter.scala 75:62]
      if (request_isSpeculative) begin // @[arbiter.scala 76:32]
        speculativeBuffer_address <= request_request_address; // @[arbiter.scala 77:24]
      end
    end
    if (reset) begin // @[arbiter.scala 62:34]
      speculativeBuffer_core_instruction <= 32'h0; // @[arbiter.scala 62:34]
    end else if (request_request_valid & request_request_branch_valid) begin // @[arbiter.scala 75:62]
      if (request_isSpeculative) begin // @[arbiter.scala 76:32]
        speculativeBuffer_core_instruction <= request_request_core_instruction; // @[arbiter.scala 77:24]
      end
    end
    if (reset) begin // @[arbiter.scala 62:34]
      speculativeBuffer_core_robAddr <= 4'h0; // @[arbiter.scala 62:34]
    end else if (request_request_valid & request_request_branch_valid) begin // @[arbiter.scala 75:62]
      if (request_isSpeculative) begin // @[arbiter.scala 76:32]
        speculativeBuffer_core_robAddr <= request_request_core_robAddr; // @[arbiter.scala 77:24]
      end
    end
    if (reset) begin // @[arbiter.scala 62:34]
      speculativeBuffer_core_prfDest <= 6'h0; // @[arbiter.scala 62:34]
    end else if (request_request_valid & request_request_branch_valid) begin // @[arbiter.scala 75:62]
      if (request_isSpeculative) begin // @[arbiter.scala 76:32]
        speculativeBuffer_core_prfDest <= request_request_core_prfDest; // @[arbiter.scala 77:24]
      end
    end
    if (reset) begin // @[arbiter.scala 62:34]
      speculativeBuffer_branch_valid <= 1'h0; // @[arbiter.scala 62:34]
    end else if (requestTypeWire != 2'h1) begin // @[arbiter.scala 153:32]
      if (speculativeBuffer_valid) begin // @[arbiter.scala 154:34]
        if (speculativeBuffer_branch_valid) begin // @[utils.scala 119:24]
          speculativeBuffer_branch_valid <= _GEN_171;
        end else begin
          speculativeBuffer_branch_valid <= _GEN_29;
        end
      end else begin
        speculativeBuffer_branch_valid <= _GEN_29;
      end
    end else begin
      speculativeBuffer_branch_valid <= _GEN_29;
    end
    if (reset) begin // @[arbiter.scala 62:34]
      speculativeBuffer_branch_mask <= 5'h0; // @[arbiter.scala 62:34]
    end else if (requestTypeWire != 2'h1) begin // @[arbiter.scala 153:32]
      if (speculativeBuffer_valid) begin // @[arbiter.scala 154:34]
        if (speculativeBuffer_branch_valid) begin // @[utils.scala 119:24]
          speculativeBuffer_branch_mask <= _GEN_170;
        end else begin
          speculativeBuffer_branch_mask <= _GEN_30;
        end
      end else begin
        speculativeBuffer_branch_mask <= _GEN_30;
      end
    end else begin
      speculativeBuffer_branch_mask <= _GEN_30;
    end
    if (reset) begin // @[arbiter.scala 63:30]
      inorderBuffer_valid <= 1'h0; // @[arbiter.scala 63:30]
    end else if (toPeripheral_ready & _T_26 & inorderBuffer_valid) begin // @[arbiter.scala 223:112]
      inorderBuffer_valid <= 1'h0; // @[arbiter.scala 224:25]
    end else if (toCacheLookup_ready) begin // @[arbiter.scala 177:72]
      if (atomicBusyState & ~toCacheLookup_holdInOrder) begin // @[arbiter.scala 178:56]
        inorderBuffer_valid <= _GEN_211;
      end else begin
        inorderBuffer_valid <= _GEN_302;
      end
    end else if (3'h0 == operationState) begin // @[arbiter.scala 107:25]
      inorderBuffer_valid <= _GEN_90;
    end else begin
      inorderBuffer_valid <= _GEN_136;
    end
    if (reset) begin // @[arbiter.scala 63:30]
      inorderBuffer_address <= 32'h0; // @[arbiter.scala 63:30]
    end else if (3'h0 == operationState) begin // @[arbiter.scala 107:25]
      if (operationBuffer_valid) begin // @[arbiter.scala 110:33]
        if (operationWires_isRead) begin // @[arbiter.scala 111:36]
          inorderBuffer_address <= operationBuffer_address; // @[arbiter.scala 113:25]
        end else begin
          inorderBuffer_address <= _GEN_64;
        end
      end
    end else if (!(3'h1 == operationState)) begin // @[arbiter.scala 107:25]
      if (3'h2 == operationState) begin // @[arbiter.scala 107:25]
        inorderBuffer_address <= _GEN_105;
      end
    end
    if (reset) begin // @[arbiter.scala 63:30]
      inorderBuffer_core_instruction <= 32'h0; // @[arbiter.scala 63:30]
    end else if (3'h0 == operationState) begin // @[arbiter.scala 107:25]
      if (operationBuffer_valid) begin // @[arbiter.scala 110:33]
        if (operationWires_isRead) begin // @[arbiter.scala 111:36]
          inorderBuffer_core_instruction <= operationBuffer_core_instruction; // @[arbiter.scala 113:25]
        end else begin
          inorderBuffer_core_instruction <= _GEN_65;
        end
      end
    end else if (!(3'h1 == operationState)) begin // @[arbiter.scala 107:25]
      if (3'h2 == operationState) begin // @[arbiter.scala 107:25]
        inorderBuffer_core_instruction <= _GEN_106;
      end
    end
    if (reset) begin // @[arbiter.scala 63:30]
      inorderBuffer_core_robAddr <= 4'h0; // @[arbiter.scala 63:30]
    end else if (3'h0 == operationState) begin // @[arbiter.scala 107:25]
      if (operationBuffer_valid) begin // @[arbiter.scala 110:33]
        if (operationWires_isRead) begin // @[arbiter.scala 111:36]
          inorderBuffer_core_robAddr <= operationBuffer_core_robAddr; // @[arbiter.scala 113:25]
        end else begin
          inorderBuffer_core_robAddr <= _GEN_66;
        end
      end
    end else if (!(3'h1 == operationState)) begin // @[arbiter.scala 107:25]
      if (3'h2 == operationState) begin // @[arbiter.scala 107:25]
        inorderBuffer_core_robAddr <= _GEN_107;
      end
    end
    if (reset) begin // @[arbiter.scala 63:30]
      inorderBuffer_core_prfDest <= 6'h0; // @[arbiter.scala 63:30]
    end else if (3'h0 == operationState) begin // @[arbiter.scala 107:25]
      if (operationBuffer_valid) begin // @[arbiter.scala 110:33]
        if (operationWires_isRead) begin // @[arbiter.scala 111:36]
          inorderBuffer_core_prfDest <= operationBuffer_core_prfDest; // @[arbiter.scala 113:25]
        end else begin
          inorderBuffer_core_prfDest <= _GEN_67;
        end
      end
    end else if (!(3'h1 == operationState)) begin // @[arbiter.scala 107:25]
      if (3'h2 == operationState) begin // @[arbiter.scala 107:25]
        inorderBuffer_core_prfDest <= _GEN_108;
      end
    end
    if (reset) begin // @[arbiter.scala 63:30]
      inorderBuffer_branch_valid <= 1'h0; // @[arbiter.scala 63:30]
    end else if (requestTypeWire != 2'h1) begin // @[arbiter.scala 153:32]
      if (inorderBuffer_valid) begin // @[arbiter.scala 160:30]
        if (inorderBuffer_branch_valid) begin // @[utils.scala 119:24]
          inorderBuffer_branch_valid <= _GEN_193;
        end else begin
          inorderBuffer_branch_valid <= _GEN_155;
        end
      end else begin
        inorderBuffer_branch_valid <= _GEN_155;
      end
    end else begin
      inorderBuffer_branch_valid <= _GEN_155;
    end
    if (reset) begin // @[arbiter.scala 63:30]
      inorderBuffer_branch_mask <= 5'h0; // @[arbiter.scala 63:30]
    end else if (requestTypeWire != 2'h1) begin // @[arbiter.scala 153:32]
      if (inorderBuffer_valid) begin // @[arbiter.scala 160:30]
        if (inorderBuffer_branch_valid) begin // @[utils.scala 119:24]
          inorderBuffer_branch_mask <= _GEN_192;
        end else begin
          inorderBuffer_branch_mask <= _GEN_156;
        end
      end else begin
        inorderBuffer_branch_mask <= _GEN_156;
      end
    end else begin
      inorderBuffer_branch_mask <= _GEN_156;
    end
    if (reset) begin // @[arbiter.scala 63:30]
      inorderBuffer_writeData_valid <= 1'h0; // @[arbiter.scala 63:30]
    end else if (3'h0 == operationState) begin // @[arbiter.scala 107:25]
      if (operationBuffer_valid) begin // @[arbiter.scala 110:33]
        if (operationWires_isRead) begin // @[arbiter.scala 111:36]
          inorderBuffer_writeData_valid <= operationBuffer_writeData_valid; // @[arbiter.scala 113:25]
        end else begin
          inorderBuffer_writeData_valid <= _GEN_70;
        end
      end
    end else if (!(3'h1 == operationState)) begin // @[arbiter.scala 107:25]
      if (3'h2 == operationState) begin // @[arbiter.scala 107:25]
        inorderBuffer_writeData_valid <= _GEN_111;
      end
    end
    if (reset) begin // @[arbiter.scala 63:30]
      inorderBuffer_writeData_data <= 64'h0; // @[arbiter.scala 63:30]
    end else if (3'h0 == operationState) begin // @[arbiter.scala 107:25]
      if (operationBuffer_valid) begin // @[arbiter.scala 110:33]
        if (operationWires_isRead) begin // @[arbiter.scala 111:36]
          inorderBuffer_writeData_data <= operationBuffer_writeData_data; // @[arbiter.scala 113:25]
        end else begin
          inorderBuffer_writeData_data <= _GEN_71;
        end
      end
    end else if (!(3'h1 == operationState)) begin // @[arbiter.scala 107:25]
      if (3'h2 == operationState) begin // @[arbiter.scala 107:25]
        inorderBuffer_writeData_data <= _GEN_112;
      end
    end
    if (reset) begin // @[arbiter.scala 64:32]
      operationBuffer_valid <= 1'h0; // @[arbiter.scala 64:32]
    end else if (3'h0 == operationState) begin // @[arbiter.scala 107:25]
      if (operationBuffer_valid) begin // @[arbiter.scala 110:33]
        if (operationWires_isRead) begin // @[arbiter.scala 111:36]
          operationBuffer_valid <= 1'h0; // @[arbiter.scala 114:33]
        end else begin
          operationBuffer_valid <= _GEN_75;
        end
      end else begin
        operationBuffer_valid <= _GEN_36;
      end
    end else if (3'h1 == operationState) begin // @[arbiter.scala 107:25]
      operationBuffer_valid <= _GEN_36;
    end else if (3'h2 == operationState) begin // @[arbiter.scala 107:25]
      operationBuffer_valid <= _GEN_116;
    end else begin
      operationBuffer_valid <= _GEN_36;
    end
    if (reset) begin // @[arbiter.scala 64:32]
      operationBuffer_address <= 32'h0; // @[arbiter.scala 64:32]
    end else if (request_request_valid & request_request_branch_valid) begin // @[arbiter.scala 75:62]
      if (!(request_isSpeculative)) begin // @[arbiter.scala 76:32]
        operationBuffer_address <= request_request_address; // @[arbiter.scala 79:23]
      end
    end
    if (reset) begin // @[arbiter.scala 64:32]
      operationBuffer_core_instruction <= 32'h0; // @[arbiter.scala 64:32]
    end else if (request_request_valid & request_request_branch_valid) begin // @[arbiter.scala 75:62]
      if (!(request_isSpeculative)) begin // @[arbiter.scala 76:32]
        operationBuffer_core_instruction <= request_request_core_instruction; // @[arbiter.scala 79:23]
      end
    end
    if (reset) begin // @[arbiter.scala 64:32]
      operationBuffer_core_robAddr <= 4'h0; // @[arbiter.scala 64:32]
    end else if (request_request_valid & request_request_branch_valid) begin // @[arbiter.scala 75:62]
      if (!(request_isSpeculative)) begin // @[arbiter.scala 76:32]
        operationBuffer_core_robAddr <= request_request_core_robAddr; // @[arbiter.scala 79:23]
      end
    end
    if (reset) begin // @[arbiter.scala 64:32]
      operationBuffer_core_prfDest <= 6'h0; // @[arbiter.scala 64:32]
    end else if (request_request_valid & request_request_branch_valid) begin // @[arbiter.scala 75:62]
      if (!(request_isSpeculative)) begin // @[arbiter.scala 76:32]
        operationBuffer_core_prfDest <= request_request_core_prfDest; // @[arbiter.scala 79:23]
      end
    end
    if (reset) begin // @[arbiter.scala 64:32]
      operationBuffer_branch_valid <= 1'h0; // @[arbiter.scala 64:32]
    end else if (requestTypeWire != 2'h1) begin // @[arbiter.scala 153:32]
      if (operationBuffer_valid) begin // @[arbiter.scala 157:32]
        if (operationBuffer_branch_valid) begin // @[utils.scala 119:24]
          operationBuffer_branch_valid <= _GEN_182;
        end else begin
          operationBuffer_branch_valid <= _GEN_41;
        end
      end else begin
        operationBuffer_branch_valid <= _GEN_41;
      end
    end else begin
      operationBuffer_branch_valid <= _GEN_41;
    end
    if (reset) begin // @[arbiter.scala 64:32]
      operationBuffer_branch_mask <= 5'h0; // @[arbiter.scala 64:32]
    end else if (requestTypeWire != 2'h1) begin // @[arbiter.scala 153:32]
      if (operationBuffer_valid) begin // @[arbiter.scala 157:32]
        if (operationBuffer_branch_valid) begin // @[utils.scala 119:24]
          operationBuffer_branch_mask <= _GEN_181;
        end else begin
          operationBuffer_branch_mask <= _GEN_42;
        end
      end else begin
        operationBuffer_branch_mask <= _GEN_42;
      end
    end else begin
      operationBuffer_branch_mask <= _GEN_42;
    end
    if (reset) begin // @[arbiter.scala 64:32]
      operationBuffer_writeData_valid <= 1'h0; // @[arbiter.scala 64:32]
    end else if (3'h0 == operationState) begin // @[arbiter.scala 107:25]
      operationBuffer_writeData_valid <= 1'h0; // @[arbiter.scala 109:38]
    end else if (request_request_valid & request_request_branch_valid) begin // @[arbiter.scala 75:62]
      if (!(request_isSpeculative)) begin // @[arbiter.scala 76:32]
        operationBuffer_writeData_valid <= request_request_writeData_valid; // @[arbiter.scala 79:23]
      end
    end
    if (reset) begin // @[arbiter.scala 64:32]
      operationBuffer_writeData_data <= 64'h0; // @[arbiter.scala 64:32]
    end else if (request_request_valid & request_request_branch_valid) begin // @[arbiter.scala 75:62]
      if (!(request_isSpeculative)) begin // @[arbiter.scala 76:32]
        operationBuffer_writeData_data <= request_request_writeData_data; // @[arbiter.scala 79:23]
      end
    end
    if (reset) begin // @[arbiter.scala 85:31]
      operationState <= 3'h0; // @[arbiter.scala 85:31]
    end else if (3'h0 == operationState) begin // @[arbiter.scala 107:25]
      if (operationBuffer_valid) begin // @[arbiter.scala 110:33]
        if (!(operationWires_isRead)) begin // @[arbiter.scala 111:36]
          operationState <= _GEN_62;
        end
      end
    end else if (3'h1 == operationState) begin // @[arbiter.scala 107:25]
      if (writeCommit_fired) begin // @[arbiter.scala 132:28]
        operationState <= 3'h2;
      end else begin
        operationState <= 3'h1;
      end
    end else if (3'h2 == operationState) begin // @[arbiter.scala 107:25]
      operationState <= _GEN_117;
    end else begin
      operationState <= _GEN_119;
    end
    if (reset) begin // @[arbiter.scala 175:32]
      atomicBusyState <= 1'h0; // @[arbiter.scala 175:32]
    end else if (toCacheLookup_ready) begin // @[arbiter.scala 177:72]
      if (atomicBusyState & ~toCacheLookup_holdInOrder) begin // @[arbiter.scala 178:56]
        if (inorderBuffer_valid & ~(operationWires_isPeriRead | operationWires_isPeriWrite)) begin // @[arbiter.scala 179:94]
          atomicBusyState <= 1'h0; // @[arbiter.scala 186:25]
        end
      end else if (!(coherencyRequest_request_valid)) begin // @[arbiter.scala 188:47]
        atomicBusyState <= _GEN_285;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  speculativeBuffer_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  speculativeBuffer_address = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  speculativeBuffer_core_instruction = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  speculativeBuffer_core_robAddr = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  speculativeBuffer_core_prfDest = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  speculativeBuffer_branch_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  speculativeBuffer_branch_mask = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  inorderBuffer_valid = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  inorderBuffer_address = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  inorderBuffer_core_instruction = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  inorderBuffer_core_robAddr = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  inorderBuffer_core_prfDest = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  inorderBuffer_branch_valid = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  inorderBuffer_branch_mask = _RAND_13[4:0];
  _RAND_14 = {1{`RANDOM}};
  inorderBuffer_writeData_valid = _RAND_14[0:0];
  _RAND_15 = {2{`RANDOM}};
  inorderBuffer_writeData_data = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  operationBuffer_valid = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  operationBuffer_address = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  operationBuffer_core_instruction = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  operationBuffer_core_robAddr = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  operationBuffer_core_prfDest = _RAND_20[5:0];
  _RAND_21 = {1{`RANDOM}};
  operationBuffer_branch_valid = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  operationBuffer_branch_mask = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  operationBuffer_writeData_valid = _RAND_23[0:0];
  _RAND_24 = {2{`RANDOM}};
  operationBuffer_writeData_data = _RAND_24[63:0];
  _RAND_25 = {1{`RANDOM}};
  operationState = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  atomicBusyState = _RAND_26[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module moduleForwardingMemory(
  input          clock,
  input  [6:0]   rdAddr,
  output [511:0] rdData,
  input  [6:0]   wrAddr,
  input  [511:0] wrData,
  input          wrEna
);
`ifdef RANDOMIZE_MEM_INIT
  reg [511:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [511:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [511:0] mem [0:127]; // @[utils.scala 30:25]
  wire  mem_memData_en; // @[utils.scala 30:25]
  wire [6:0] mem_memData_addr; // @[utils.scala 30:25]
  wire [511:0] mem_memData_data; // @[utils.scala 30:25]
  wire [511:0] mem_MPORT_data; // @[utils.scala 30:25]
  wire [6:0] mem_MPORT_addr; // @[utils.scala 30:25]
  wire  mem_MPORT_mask; // @[utils.scala 30:25]
  wire  mem_MPORT_en; // @[utils.scala 30:25]
  reg  mem_memData_en_pipe_0;
  reg [6:0] mem_memData_addr_pipe_0;
  reg [511:0] wrDataReg; // @[utils.scala 32:27]
  reg  doForwardReg; // @[utils.scala 33:30]
  assign mem_memData_en = mem_memData_en_pipe_0;
  assign mem_memData_addr = mem_memData_addr_pipe_0;
  assign mem_memData_data = mem[mem_memData_addr]; // @[utils.scala 30:25]
  assign mem_MPORT_data = wrData;
  assign mem_MPORT_addr = wrAddr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = wrEna;
  assign rdData = doForwardReg ? wrDataReg : mem_memData_data; // @[utils.scala 40:15]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[utils.scala 30:25]
    end
    mem_memData_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      mem_memData_addr_pipe_0 <= rdAddr;
    end
    wrDataReg <= wrData; // @[utils.scala 32:27]
    doForwardReg <= wrAddr == rdAddr & wrEna; // @[utils.scala 33:49]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {16{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    mem[initvar] = _RAND_0[511:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_memData_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_memData_addr_pipe_0 = _RAND_2[6:0];
  _RAND_3 = {16{`RANDOM}};
  wrDataReg = _RAND_3[511:0];
  _RAND_4 = {1{`RANDOM}};
  doForwardReg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module moduleForwardingMemory_4(
  input         clock,
  input  [6:0]  rdAddr,
  output [91:0] rdData,
  input  [6:0]  wrAddr,
  input  [91:0] wrData,
  input         wrEna
);
`ifdef RANDOMIZE_MEM_INIT
  reg [95:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [95:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [91:0] mem [0:127]; // @[utils.scala 30:25]
  wire  mem_memData_en; // @[utils.scala 30:25]
  wire [6:0] mem_memData_addr; // @[utils.scala 30:25]
  wire [91:0] mem_memData_data; // @[utils.scala 30:25]
  wire [91:0] mem_MPORT_data; // @[utils.scala 30:25]
  wire [6:0] mem_MPORT_addr; // @[utils.scala 30:25]
  wire  mem_MPORT_mask; // @[utils.scala 30:25]
  wire  mem_MPORT_en; // @[utils.scala 30:25]
  reg  mem_memData_en_pipe_0;
  reg [6:0] mem_memData_addr_pipe_0;
  reg [91:0] wrDataReg; // @[utils.scala 32:27]
  reg  doForwardReg; // @[utils.scala 33:30]
  assign mem_memData_en = mem_memData_en_pipe_0;
  assign mem_memData_addr = mem_memData_addr_pipe_0;
  assign mem_memData_data = mem[mem_memData_addr]; // @[utils.scala 30:25]
  assign mem_MPORT_data = wrData;
  assign mem_MPORT_addr = wrAddr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = wrEna;
  assign rdData = doForwardReg ? wrDataReg : mem_memData_data; // @[utils.scala 40:15]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[utils.scala 30:25]
    end
    mem_memData_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      mem_memData_addr_pipe_0 <= rdAddr;
    end
    wrDataReg <= wrData; // @[utils.scala 32:27]
    doForwardReg <= wrAddr == rdAddr & wrEna; // @[utils.scala 33:49]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {3{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    mem[initvar] = _RAND_0[91:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_memData_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_memData_addr_pipe_0 = _RAND_2[6:0];
  _RAND_3 = {3{`RANDOM}};
  wrDataReg = _RAND_3[91:0];
  _RAND_4 = {1{`RANDOM}};
  doForwardReg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module cacheLookupUnit(
  input          clock,
  input          reset,
  output         request_ready,
  output         request_holdInOrder,
  input  [1:0]   request_requestType,
  input          request_request_valid,
  input  [31:0]  request_request_address,
  input  [31:0]  request_request_core_instruction,
  input  [3:0]   request_request_core_robAddr,
  input  [5:0]   request_request_core_prfDest,
  input          request_request_branch_valid,
  input  [4:0]   request_request_branch_mask,
  input          request_request_writeData_valid,
  input  [63:0]  request_request_writeData_data,
  input  [511:0] request_request_cacheLine_cacheLine,
  input  [1:0]   request_request_cacheLine_response,
  input          toReplay_ready,
  output         toReplay_request_valid,
  output [31:0]  toReplay_request_address,
  output [31:0]  toReplay_request_core_instruction,
  output [3:0]   toReplay_request_core_robAddr,
  output [5:0]   toReplay_request_core_prfDest,
  output         toReplay_request_branch_valid,
  output [4:0]   toReplay_request_branch_mask,
  output         toReplay_request_writeData_valid,
  output [63:0]  toReplay_request_writeData_data,
  output [1:0]   toReplay_request_cacheLine_response,
  input          toWriteBack_ready,
  output         toWriteBack_request_valid,
  output [31:0]  toWriteBack_request_address,
  output [511:0] toWriteBack_request_data,
  input          toCoherency_ready,
  output         toCoherency_request_valid,
  output [1:0]   toCoherency_request_response,
  output [511:0] toCoherency_request_cacheLine,
  output         toCoherency_request_dataValid,
  output         toResponse_request_valid,
  output [31:0]  toResponse_request_address,
  output [31:0]  toResponse_request_core_instruction,
  output [3:0]   toResponse_request_core_robAddr,
  output [5:0]   toResponse_request_core_prfDest,
  output         toResponse_request_branch_valid,
  output [4:0]   toResponse_request_branch_mask,
  output [63:0]  toResponse_request_writeData_data,
  output         writeInstructionCommit_ready,
  input          writeInstructionCommit_fired,
  input          branchOps_valid,
  input  [4:0]   branchOps_branchMask,
  input          branchOps_passed
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [511:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [511:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [511:0] _RAND_47;
  reg [31:0] _RAND_48;
`endif // RANDOMIZE_REG_INIT
  wire  dataBRAM_0_clock; // @[cacheLookupUnit.scala 60:39]
  wire [6:0] dataBRAM_0_rdAddr; // @[cacheLookupUnit.scala 60:39]
  wire [511:0] dataBRAM_0_rdData; // @[cacheLookupUnit.scala 60:39]
  wire [6:0] dataBRAM_0_wrAddr; // @[cacheLookupUnit.scala 60:39]
  wire [511:0] dataBRAM_0_wrData; // @[cacheLookupUnit.scala 60:39]
  wire  dataBRAM_0_wrEna; // @[cacheLookupUnit.scala 60:39]
  wire  dataBRAM_1_clock; // @[cacheLookupUnit.scala 60:39]
  wire [6:0] dataBRAM_1_rdAddr; // @[cacheLookupUnit.scala 60:39]
  wire [511:0] dataBRAM_1_rdData; // @[cacheLookupUnit.scala 60:39]
  wire [6:0] dataBRAM_1_wrAddr; // @[cacheLookupUnit.scala 60:39]
  wire [511:0] dataBRAM_1_wrData; // @[cacheLookupUnit.scala 60:39]
  wire  dataBRAM_1_wrEna; // @[cacheLookupUnit.scala 60:39]
  wire  dataBRAM_2_clock; // @[cacheLookupUnit.scala 60:39]
  wire [6:0] dataBRAM_2_rdAddr; // @[cacheLookupUnit.scala 60:39]
  wire [511:0] dataBRAM_2_rdData; // @[cacheLookupUnit.scala 60:39]
  wire [6:0] dataBRAM_2_wrAddr; // @[cacheLookupUnit.scala 60:39]
  wire [511:0] dataBRAM_2_wrData; // @[cacheLookupUnit.scala 60:39]
  wire  dataBRAM_2_wrEna; // @[cacheLookupUnit.scala 60:39]
  wire  dataBRAM_3_clock; // @[cacheLookupUnit.scala 60:39]
  wire [6:0] dataBRAM_3_rdAddr; // @[cacheLookupUnit.scala 60:39]
  wire [511:0] dataBRAM_3_rdData; // @[cacheLookupUnit.scala 60:39]
  wire [6:0] dataBRAM_3_wrAddr; // @[cacheLookupUnit.scala 60:39]
  wire [511:0] dataBRAM_3_wrData; // @[cacheLookupUnit.scala 60:39]
  wire  dataBRAM_3_wrEna; // @[cacheLookupUnit.scala 60:39]
  wire  tagBRAM_clock; // @[cacheLookupUnit.scala 110:23]
  wire [6:0] tagBRAM_rdAddr; // @[cacheLookupUnit.scala 110:23]
  wire [91:0] tagBRAM_rdData; // @[cacheLookupUnit.scala 110:23]
  wire [6:0] tagBRAM_wrAddr; // @[cacheLookupUnit.scala 110:23]
  wire [91:0] tagBRAM_wrData; // @[cacheLookupUnit.scala 110:23]
  wire  tagBRAM_wrEna; // @[cacheLookupUnit.scala 110:23]
  wire  _operationValid_T_1 = request_ready & request_request_valid & request_request_branch_valid; // @[cacheLookupUnit.scala 52:71]
  reg  operationValid; // @[cacheLookupUnit.scala 52:31]
  reg [31:0] reservationRegister_address; // @[cacheLookupUnit.scala 121:36]
  reg  reservationRegister_reserved; // @[cacheLookupUnit.scala 121:36]
  reg  reservationRegister_size; // @[cacheLookupUnit.scala 121:36]
  reg  lastMissRecordRegister_valid; // @[cacheLookupUnit.scala 130:39]
  reg [31:0] lastMissRecordRegister_address; // @[cacheLookupUnit.scala 130:39]
  reg [31:0] lastMissRecordRegister_core_instruction; // @[cacheLookupUnit.scala 130:39]
  reg [3:0] lastMissRecordRegister_core_robAddr; // @[cacheLookupUnit.scala 130:39]
  reg [5:0] lastMissRecordRegister_core_prfDest; // @[cacheLookupUnit.scala 130:39]
  reg  lastMissRecordRegister_branch_valid; // @[cacheLookupUnit.scala 130:39]
  reg [4:0] lastMissRecordRegister_branch_mask; // @[cacheLookupUnit.scala 130:39]
  wire  _replayMatch_T_1 = request_request_core_instruction == lastMissRecordRegister_core_instruction; // @[cacheLookupUnit.scala 136:41]
  wire  _replayMatch_T_2 = request_request_address == lastMissRecordRegister_address & _replayMatch_T_1; // @[cacheLookupUnit.scala 135:68]
  wire  _replayMatch_T_3 = request_request_core_robAddr == lastMissRecordRegister_core_robAddr; // @[cacheLookupUnit.scala 137:37]
  wire  _replayMatch_T_4 = _replayMatch_T_2 & _replayMatch_T_3; // @[cacheLookupUnit.scala 136:86]
  wire  _replayMatch_T_5 = request_request_core_prfDest == lastMissRecordRegister_core_prfDest; // @[cacheLookupUnit.scala 138:37]
  wire  replayMatch = _replayMatch_T_4 & _replayMatch_T_5; // @[cacheLookupUnit.scala 137:78]
  wire  _GEN_0 = replayMatch ? 1'h0 : lastMissRecordRegister_valid; // @[cacheLookupUnit.scala 140:22 141:36 130:39]
  wire  _GEN_1 = _operationValid_T_1 & lastMissRecordRegister_valid ? _GEN_0 : lastMissRecordRegister_valid; // @[cacheLookupUnit.scala 133:111 130:39]
  reg  readBuffer_valid; // @[cacheLookupUnit.scala 146:27]
  reg [31:0] readBuffer_address; // @[cacheLookupUnit.scala 146:27]
  reg [31:0] readBuffer_core_instruction; // @[cacheLookupUnit.scala 146:27]
  reg [3:0] readBuffer_core_robAddr; // @[cacheLookupUnit.scala 146:27]
  reg [5:0] readBuffer_core_prfDest; // @[cacheLookupUnit.scala 146:27]
  reg  readBuffer_branch_valid; // @[cacheLookupUnit.scala 146:27]
  reg [4:0] readBuffer_branch_mask; // @[cacheLookupUnit.scala 146:27]
  reg  readBuffer_writeData_valid; // @[cacheLookupUnit.scala 146:27]
  reg [63:0] readBuffer_writeData_data; // @[cacheLookupUnit.scala 146:27]
  reg [511:0] readBuffer_cacheLine_cacheLine; // @[cacheLookupUnit.scala 146:27]
  reg [1:0] readBuffer_cacheLine_response; // @[cacheLookupUnit.scala 146:27]
  reg [1:0] requestType; // @[cacheLookupUnit.scala 147:28]
  reg  replayBuffer_valid; // @[cacheLookupUnit.scala 153:29]
  reg [31:0] replayBuffer_address; // @[cacheLookupUnit.scala 153:29]
  reg [31:0] replayBuffer_core_instruction; // @[cacheLookupUnit.scala 153:29]
  reg [3:0] replayBuffer_core_robAddr; // @[cacheLookupUnit.scala 153:29]
  reg [5:0] replayBuffer_core_prfDest; // @[cacheLookupUnit.scala 153:29]
  reg  replayBuffer_branch_valid; // @[cacheLookupUnit.scala 153:29]
  reg [4:0] replayBuffer_branch_mask; // @[cacheLookupUnit.scala 153:29]
  reg  replayBuffer_writeData_valid; // @[cacheLookupUnit.scala 153:29]
  reg [63:0] replayBuffer_writeData_data; // @[cacheLookupUnit.scala 153:29]
  reg [1:0] replayBuffer_cacheLine_response; // @[cacheLookupUnit.scala 153:29]
  wire  _GEN_14 = toReplay_ready ? 1'h0 : replayBuffer_valid; // @[cacheLookupUnit.scala 155:23 157:24 153:29]
  reg  memoryResponseBuffer_valid; // @[cacheLookupUnit.scala 160:37]
  reg [31:0] memoryResponseBuffer_address; // @[cacheLookupUnit.scala 160:37]
  reg [31:0] memoryResponseBuffer_core_instruction; // @[cacheLookupUnit.scala 160:37]
  reg [3:0] memoryResponseBuffer_core_robAddr; // @[cacheLookupUnit.scala 160:37]
  reg [5:0] memoryResponseBuffer_core_prfDest; // @[cacheLookupUnit.scala 160:37]
  reg  memoryResponseBuffer_branch_valid; // @[cacheLookupUnit.scala 160:37]
  reg [4:0] memoryResponseBuffer_branch_mask; // @[cacheLookupUnit.scala 160:37]
  reg [63:0] memoryResponseBuffer_writeData_data; // @[cacheLookupUnit.scala 160:37]
  wire [4:0] _T_4 = memoryResponseBuffer_branch_mask & branchOps_branchMask; // @[utils.scala 92:27]
  wire  _T_5 = |_T_4; // @[utils.scala 92:51]
  wire [4:0] _toResponse_request_branch_mask_T = memoryResponseBuffer_branch_mask ^ branchOps_branchMask; // @[utils.scala 93:42]
  wire [4:0] _GEN_15 = |_T_4 ? _toResponse_request_branch_mask_T : memoryResponseBuffer_branch_mask; // @[utils.scala 92:56 93:27 96:27]
  wire [4:0] _GEN_16 = _T_5 ? 5'h0 : memoryResponseBuffer_branch_mask; // @[utils.scala 101:56 102:27 106:27]
  wire  _GEN_17 = _T_5 ? 1'h0 : memoryResponseBuffer_branch_valid; // @[utils.scala 101:56 103:28 107:28]
  wire [4:0] _GEN_18 = branchOps_passed ? _GEN_15 : _GEN_16; // @[utils.scala 90:30]
  wire  _GEN_19 = branchOps_passed ? memoryResponseBuffer_branch_valid : _GEN_17; // @[utils.scala 90:30 98:26]
  wire [4:0] _GEN_20 = branchOps_valid ? _GEN_18 : memoryResponseBuffer_branch_mask; // @[utils.scala 111:23 89:27]
  wire  _GEN_21 = branchOps_valid ? _GEN_19 : memoryResponseBuffer_branch_valid; // @[utils.scala 112:24 89:27]
  wire  _GEN_34 = memoryResponseBuffer_valid ? 1'h0 : memoryResponseBuffer_valid; // @[cacheLookupUnit.scala 166:35 167:32 160:37]
  reg  coherencyResponseBuffer_valid; // @[cacheLookupUnit.scala 170:40]
  reg [1:0] coherencyResponseBuffer_response; // @[cacheLookupUnit.scala 170:40]
  reg [511:0] coherencyResponseBuffer_cacheLine; // @[cacheLookupUnit.scala 170:40]
  reg  coherencyResponseBuffer_dataValid; // @[cacheLookupUnit.scala 170:40]
  wire  _GEN_40 = toCoherency_ready ? 1'h0 : coherencyResponseBuffer_valid; // @[cacheLookupUnit.scala 172:26 174:35 170:40]
  reg  writeBackBuffer_valid; // @[cacheLookupUnit.scala 177:32]
  reg [31:0] writeBackBuffer_address; // @[cacheLookupUnit.scala 177:32]
  reg [511:0] writeBackBuffer_data; // @[cacheLookupUnit.scala 177:32]
  wire  _GEN_44 = toWriteBack_ready ? 1'h0 : writeBackBuffer_valid; // @[cacheLookupUnit.scala 179:26 181:27 177:32]
  reg  writeCommitInstructionBuffer; // @[cacheLookupUnit.scala 184:45]
  wire  _GEN_45 = writeInstructionCommit_fired ? 1'h0 : writeCommitInstructionBuffer; // @[cacheLookupUnit.scala 186:37 187:34 184:45]
  wire  _request_holdInOrder_T = lastMissRecordRegister_valid & lastMissRecordRegister_branch_valid; // @[cacheLookupUnit.scala 194:55]
  wire  _GEN_51 = request_request_valid & request_request_branch_valid & request_request_valid; // @[cacheLookupUnit.scala 203:62 207:16 210:22]
  wire  _GEN_56 = request_request_valid & request_request_branch_valid ? request_request_branch_valid :
    readBuffer_branch_valid; // @[cacheLookupUnit.scala 203:62 207:16 146:27]
  wire [4:0] _GEN_57 = request_request_valid & request_request_branch_valid ? request_request_branch_mask :
    readBuffer_branch_mask; // @[cacheLookupUnit.scala 203:62 207:16 146:27]
  wire  isReadWire = readBuffer_core_instruction[6:0] == 7'h3; // @[cacheLookupUnit.scala 214:67]
  wire  isWriteWire = readBuffer_core_instruction[6:0] == 7'h23; // @[cacheLookupUnit.scala 215:68]
  wire  isCoherentWire = requestType == 2'h3; // @[cacheLookupUnit.scala 216:50]
  wire  isAtomicsWire = readBuffer_core_instruction[6:0] == 7'h2f; // @[cacheLookupUnit.scala 217:71]
  wire  isLRWire = readBuffer_core_instruction[31:27] == 5'h2 & isAtomicsWire; // @[cacheLookupUnit.scala 218:82]
  wire  isSCWire = readBuffer_core_instruction[31:27] == 5'h3 & isAtomicsWire; // @[cacheLookupUnit.scala 219:82]
  wire  _isAtmoicReadWire_T = ~readBuffer_writeData_valid; // @[cacheLookupUnit.scala 220:57]
  wire  _isAtmoicReadWire_T_3 = ~(isSCWire | isLRWire); // @[cacheLookupUnit.scala 220:88]
  wire  isAtmoicReadWire = isAtomicsWire & ~readBuffer_writeData_valid & ~(isSCWire | isLRWire); // @[cacheLookupUnit.scala 220:85]
  wire  isAtmoicWriteWire = isAtomicsWire & readBuffer_writeData_valid & _isAtmoicReadWire_T_3; // @[cacheLookupUnit.scala 221:85]
  wire  isLRReadWire = isLRWire & _isAtmoicReadWire_T; // @[cacheLookupUnit.scala 222:45]
  wire  isLRWriteWire = isLRWire & readBuffer_writeData_valid; // @[cacheLookupUnit.scala 223:46]
  wire  isSCReadWire = isSCWire & _isAtmoicReadWire_T; // @[cacheLookupUnit.scala 224:45]
  wire  isSCWriteWire = isSCWire & readBuffer_writeData_valid; // @[cacheLookupUnit.scala 225:46]
  wire [22:0] tagChunks_0 = tagBRAM_rdData[22:0]; // @[cacheLookupUnit.scala 230:21]
  wire [22:0] tagChunks_1 = tagBRAM_rdData[45:23]; // @[cacheLookupUnit.scala 230:21]
  wire [22:0] tagChunks_2 = tagBRAM_rdData[68:46]; // @[cacheLookupUnit.scala 230:21]
  wire [22:0] tagChunks_3 = tagBRAM_rdData[91:69]; // @[cacheLookupUnit.scala 230:21]
  wire  matchFoundVec_0 = tagChunks_0[18:0] == readBuffer_address[31:13]; // @[cacheLookupUnit.scala 236:25]
  wire  matchFoundVec_1 = tagChunks_1[18:0] == readBuffer_address[31:13]; // @[cacheLookupUnit.scala 236:25]
  wire  matchFoundVec_2 = tagChunks_2[18:0] == readBuffer_address[31:13]; // @[cacheLookupUnit.scala 236:25]
  wire  matchFoundVec_3 = tagChunks_3[18:0] == readBuffer_address[31:13]; // @[cacheLookupUnit.scala 236:25]
  wire [1:0] _hitTagWire_T = matchFoundVec_2 ? 2'h2 : 2'h3; // @[Mux.scala 47:70]
  wire [1:0] _hitTagWire_T_1 = matchFoundVec_1 ? 2'h1 : _hitTagWire_T; // @[Mux.scala 47:70]
  wire [1:0] hitTagWire = matchFoundVec_0 ? 2'h0 : _hitTagWire_T_1; // @[Mux.scala 47:70]
  wire [22:0] _GEN_65 = 2'h1 == hitTagWire ? tagChunks_1 : tagChunks_0; // @[cacheLookupUnit.scala 239:{57,57}]
  wire [22:0] _GEN_66 = 2'h2 == hitTagWire ? tagChunks_2 : _GEN_65; // @[cacheLookupUnit.scala 239:{57,57}]
  wire [22:0] _GEN_67 = 2'h3 == hitTagWire ? tagChunks_3 : _GEN_66; // @[cacheLookupUnit.scala 239:{57,57}]
  wire  validBitWire = _GEN_67[19]; // @[cacheLookupUnit.scala 239:57]
  wire  shareBitWire = _GEN_67[21]; // @[cacheLookupUnit.scala 240:57]
  wire  dirtyBitWire = _GEN_67[20]; // @[cacheLookupUnit.scala 241:57]
  wire  isDirtyWire = dirtyBitWire & validBitWire; // @[cacheLookupUnit.scala 244:48]
  wire  isSharedWire = shareBitWire & validBitWire; // @[cacheLookupUnit.scala 245:49]
  wire  isDataMissWire = ~((matchFoundVec_0 | matchFoundVec_1 | matchFoundVec_2 | matchFoundVec_3) & validBitWire); // @[cacheLookupUnit.scala 246:38]
  wire  _isPermissionMiss_T = ~isDataMissWire; // @[cacheLookupUnit.scala 247:40]
  wire  isPermissionMiss = ~isDataMissWire & isSharedWire; // @[cacheLookupUnit.scala 247:56]
  wire  isReplayValidWire = requestType == 2'h2; // @[cacheLookupUnit.scala 248:53]
  wire  _cacheLineChoosen_T = isDataMissWire & isReplayValidWire; // @[cacheLookupUnit.scala 261:47]
  wire [511:0] dataBRAMVec_0_rdData = dataBRAM_0_rdData; // @[cacheLookupUnit.scala 75:28 93:16]
  wire [511:0] dataBRAMVec_1_rdData = dataBRAM_1_rdData; // @[cacheLookupUnit.scala 75:28 93:16]
  wire [511:0] _GEN_101 = 2'h1 == hitTagWire ? dataBRAMVec_1_rdData : dataBRAMVec_0_rdData; // @[cacheLookupUnit.scala 261:{31,31}]
  wire [511:0] dataBRAMVec_2_rdData = dataBRAM_2_rdData; // @[cacheLookupUnit.scala 75:28 93:16]
  wire [511:0] _GEN_102 = 2'h2 == hitTagWire ? dataBRAMVec_2_rdData : _GEN_101; // @[cacheLookupUnit.scala 261:{31,31}]
  wire [511:0] dataBRAMVec_3_rdData = dataBRAM_3_rdData; // @[cacheLookupUnit.scala 75:28 93:16]
  wire [511:0] _GEN_103 = 2'h3 == hitTagWire ? dataBRAMVec_3_rdData : _GEN_102; // @[cacheLookupUnit.scala 261:{31,31}]
  wire [511:0] cacheLineChoosen = isDataMissWire & isReplayValidWire ? readBuffer_cacheLine_cacheLine : _GEN_103; // @[cacheLookupUnit.scala 261:31]
  wire [3:0] _doubleWordWrite_T_1 = {readBuffer_address[5:3],1'h1}; // @[cacheLookupUnit.scala 269:68]
  wire [3:0] _doubleWordWrite_T_3 = {readBuffer_address[5:3],1'h0}; // @[cacheLookupUnit.scala 269:114]
  wire  _T_14 = isWriteWire | isAtmoicWriteWire; // @[cacheLookupUnit.scala 313:22]
  wire  _T_18 = ~isPermissionMiss & _isPermissionMiss_T; // @[cacheLookupUnit.scala 314:30]
  wire  _T_10 = isLRReadWire | isAtmoicReadWire; // @[cacheLookupUnit.scala 295:23]
  wire [31:0] _GEN_145 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[31:0] : cacheLineChoosen[31:0]; // @[cacheLookupUnit.scala 284:37 291:26 262:30]
  wire [31:0] _GEN_166 = _isPermissionMiss_T ? cacheLineChoosen[31:0] : _GEN_145; // @[cacheLookupUnit.scala 282:28 262:30]
  wire [31:0] _GEN_187 = isReadWire ? _GEN_166 : cacheLineChoosen[31:0]; // @[cacheLookupUnit.scala 281:21 262:30]
  wire [31:0] _GEN_208 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[31:0] : _GEN_187; // @[cacheLookupUnit.scala 298:37 305:26]
  wire [31:0] _GEN_229 = _T_18 ? _GEN_187 : _GEN_208; // @[cacheLookupUnit.scala 296:49]
  wire [31:0] _GEN_250 = isLRReadWire | isAtmoicReadWire ? _GEN_229 : _GEN_187; // @[cacheLookupUnit.scala 295:43]
  wire [31:0] _GEN_274 = isReplayValidWire & isDataMissWire ? readBuffer_cacheLine_cacheLine[31:0] : _GEN_250; // @[cacheLookupUnit.scala 317:55 324:26]
  wire [31:0] _GEN_295 = ~isPermissionMiss & _isPermissionMiss_T ? _GEN_250 : _GEN_274; // @[cacheLookupUnit.scala 314:49]
  wire [31:0] writeChunks_0 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_295 : _GEN_250; // @[cacheLookupUnit.scala 313:61]
  wire [31:0] _GEN_146 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[63:32] : cacheLineChoosen[63:32]; // @[cacheLookupUnit.scala 284:37 291:26 262:30]
  wire [31:0] _GEN_167 = _isPermissionMiss_T ? cacheLineChoosen[63:32] : _GEN_146; // @[cacheLookupUnit.scala 282:28 262:30]
  wire [31:0] _GEN_188 = isReadWire ? _GEN_167 : cacheLineChoosen[63:32]; // @[cacheLookupUnit.scala 281:21 262:30]
  wire [31:0] _GEN_209 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[63:32] : _GEN_188; // @[cacheLookupUnit.scala 298:37 305:26]
  wire [31:0] _GEN_230 = _T_18 ? _GEN_188 : _GEN_209; // @[cacheLookupUnit.scala 296:49]
  wire [31:0] _GEN_251 = isLRReadWire | isAtmoicReadWire ? _GEN_230 : _GEN_188; // @[cacheLookupUnit.scala 295:43]
  wire [31:0] _GEN_275 = isReplayValidWire & isDataMissWire ? readBuffer_cacheLine_cacheLine[63:32] : _GEN_251; // @[cacheLookupUnit.scala 317:55 324:26]
  wire [31:0] _GEN_296 = ~isPermissionMiss & _isPermissionMiss_T ? _GEN_251 : _GEN_275; // @[cacheLookupUnit.scala 314:49]
  wire [31:0] writeChunks_1 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_296 : _GEN_251; // @[cacheLookupUnit.scala 313:61]
  wire [31:0] _GEN_105 = 4'h1 == _doubleWordWrite_T_1 ? writeChunks_1 : writeChunks_0; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_147 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[95:64] : cacheLineChoosen[95:64]; // @[cacheLookupUnit.scala 284:37 291:26 262:30]
  wire [31:0] _GEN_168 = _isPermissionMiss_T ? cacheLineChoosen[95:64] : _GEN_147; // @[cacheLookupUnit.scala 282:28 262:30]
  wire [31:0] _GEN_189 = isReadWire ? _GEN_168 : cacheLineChoosen[95:64]; // @[cacheLookupUnit.scala 281:21 262:30]
  wire [31:0] _GEN_210 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[95:64] : _GEN_189; // @[cacheLookupUnit.scala 298:37 305:26]
  wire [31:0] _GEN_231 = _T_18 ? _GEN_189 : _GEN_210; // @[cacheLookupUnit.scala 296:49]
  wire [31:0] _GEN_252 = isLRReadWire | isAtmoicReadWire ? _GEN_231 : _GEN_189; // @[cacheLookupUnit.scala 295:43]
  wire [31:0] _GEN_276 = isReplayValidWire & isDataMissWire ? readBuffer_cacheLine_cacheLine[95:64] : _GEN_252; // @[cacheLookupUnit.scala 317:55 324:26]
  wire [31:0] _GEN_297 = ~isPermissionMiss & _isPermissionMiss_T ? _GEN_252 : _GEN_276; // @[cacheLookupUnit.scala 314:49]
  wire [31:0] writeChunks_2 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_297 : _GEN_252; // @[cacheLookupUnit.scala 313:61]
  wire [31:0] _GEN_106 = 4'h2 == _doubleWordWrite_T_1 ? writeChunks_2 : _GEN_105; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_148 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[127:96] : cacheLineChoosen[127:96]; // @[cacheLookupUnit.scala 284:37 291:26 262:30]
  wire [31:0] _GEN_169 = _isPermissionMiss_T ? cacheLineChoosen[127:96] : _GEN_148; // @[cacheLookupUnit.scala 282:28 262:30]
  wire [31:0] _GEN_190 = isReadWire ? _GEN_169 : cacheLineChoosen[127:96]; // @[cacheLookupUnit.scala 281:21 262:30]
  wire [31:0] _GEN_211 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[127:96] : _GEN_190; // @[cacheLookupUnit.scala 298:37 305:26]
  wire [31:0] _GEN_232 = _T_18 ? _GEN_190 : _GEN_211; // @[cacheLookupUnit.scala 296:49]
  wire [31:0] _GEN_253 = isLRReadWire | isAtmoicReadWire ? _GEN_232 : _GEN_190; // @[cacheLookupUnit.scala 295:43]
  wire [31:0] _GEN_277 = isReplayValidWire & isDataMissWire ? readBuffer_cacheLine_cacheLine[127:96] : _GEN_253; // @[cacheLookupUnit.scala 317:55 324:26]
  wire [31:0] _GEN_298 = ~isPermissionMiss & _isPermissionMiss_T ? _GEN_253 : _GEN_277; // @[cacheLookupUnit.scala 314:49]
  wire [31:0] writeChunks_3 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_298 : _GEN_253; // @[cacheLookupUnit.scala 313:61]
  wire [31:0] _GEN_107 = 4'h3 == _doubleWordWrite_T_1 ? writeChunks_3 : _GEN_106; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_149 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[159:128] : cacheLineChoosen[159:128]; // @[cacheLookupUnit.scala 284:37 291:26 262:30]
  wire [31:0] _GEN_170 = _isPermissionMiss_T ? cacheLineChoosen[159:128] : _GEN_149; // @[cacheLookupUnit.scala 282:28 262:30]
  wire [31:0] _GEN_191 = isReadWire ? _GEN_170 : cacheLineChoosen[159:128]; // @[cacheLookupUnit.scala 281:21 262:30]
  wire [31:0] _GEN_212 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[159:128] : _GEN_191; // @[cacheLookupUnit.scala 298:37 305:26]
  wire [31:0] _GEN_233 = _T_18 ? _GEN_191 : _GEN_212; // @[cacheLookupUnit.scala 296:49]
  wire [31:0] _GEN_254 = isLRReadWire | isAtmoicReadWire ? _GEN_233 : _GEN_191; // @[cacheLookupUnit.scala 295:43]
  wire [31:0] _GEN_278 = isReplayValidWire & isDataMissWire ? readBuffer_cacheLine_cacheLine[159:128] : _GEN_254; // @[cacheLookupUnit.scala 317:55 324:26]
  wire [31:0] _GEN_299 = ~isPermissionMiss & _isPermissionMiss_T ? _GEN_254 : _GEN_278; // @[cacheLookupUnit.scala 314:49]
  wire [31:0] writeChunks_4 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_299 : _GEN_254; // @[cacheLookupUnit.scala 313:61]
  wire [31:0] _GEN_108 = 4'h4 == _doubleWordWrite_T_1 ? writeChunks_4 : _GEN_107; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_150 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[191:160] : cacheLineChoosen[191:160]; // @[cacheLookupUnit.scala 284:37 291:26 262:30]
  wire [31:0] _GEN_171 = _isPermissionMiss_T ? cacheLineChoosen[191:160] : _GEN_150; // @[cacheLookupUnit.scala 282:28 262:30]
  wire [31:0] _GEN_192 = isReadWire ? _GEN_171 : cacheLineChoosen[191:160]; // @[cacheLookupUnit.scala 281:21 262:30]
  wire [31:0] _GEN_213 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[191:160] : _GEN_192; // @[cacheLookupUnit.scala 298:37 305:26]
  wire [31:0] _GEN_234 = _T_18 ? _GEN_192 : _GEN_213; // @[cacheLookupUnit.scala 296:49]
  wire [31:0] _GEN_255 = isLRReadWire | isAtmoicReadWire ? _GEN_234 : _GEN_192; // @[cacheLookupUnit.scala 295:43]
  wire [31:0] _GEN_279 = isReplayValidWire & isDataMissWire ? readBuffer_cacheLine_cacheLine[191:160] : _GEN_255; // @[cacheLookupUnit.scala 317:55 324:26]
  wire [31:0] _GEN_300 = ~isPermissionMiss & _isPermissionMiss_T ? _GEN_255 : _GEN_279; // @[cacheLookupUnit.scala 314:49]
  wire [31:0] writeChunks_5 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_300 : _GEN_255; // @[cacheLookupUnit.scala 313:61]
  wire [31:0] _GEN_109 = 4'h5 == _doubleWordWrite_T_1 ? writeChunks_5 : _GEN_108; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_151 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[223:192] : cacheLineChoosen[223:192]; // @[cacheLookupUnit.scala 284:37 291:26 262:30]
  wire [31:0] _GEN_172 = _isPermissionMiss_T ? cacheLineChoosen[223:192] : _GEN_151; // @[cacheLookupUnit.scala 282:28 262:30]
  wire [31:0] _GEN_193 = isReadWire ? _GEN_172 : cacheLineChoosen[223:192]; // @[cacheLookupUnit.scala 281:21 262:30]
  wire [31:0] _GEN_214 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[223:192] : _GEN_193; // @[cacheLookupUnit.scala 298:37 305:26]
  wire [31:0] _GEN_235 = _T_18 ? _GEN_193 : _GEN_214; // @[cacheLookupUnit.scala 296:49]
  wire [31:0] _GEN_256 = isLRReadWire | isAtmoicReadWire ? _GEN_235 : _GEN_193; // @[cacheLookupUnit.scala 295:43]
  wire [31:0] _GEN_280 = isReplayValidWire & isDataMissWire ? readBuffer_cacheLine_cacheLine[223:192] : _GEN_256; // @[cacheLookupUnit.scala 317:55 324:26]
  wire [31:0] _GEN_301 = ~isPermissionMiss & _isPermissionMiss_T ? _GEN_256 : _GEN_280; // @[cacheLookupUnit.scala 314:49]
  wire [31:0] writeChunks_6 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_301 : _GEN_256; // @[cacheLookupUnit.scala 313:61]
  wire [31:0] _GEN_110 = 4'h6 == _doubleWordWrite_T_1 ? writeChunks_6 : _GEN_109; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_152 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[255:224] : cacheLineChoosen[255:224]; // @[cacheLookupUnit.scala 284:37 291:26 262:30]
  wire [31:0] _GEN_173 = _isPermissionMiss_T ? cacheLineChoosen[255:224] : _GEN_152; // @[cacheLookupUnit.scala 282:28 262:30]
  wire [31:0] _GEN_194 = isReadWire ? _GEN_173 : cacheLineChoosen[255:224]; // @[cacheLookupUnit.scala 281:21 262:30]
  wire [31:0] _GEN_215 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[255:224] : _GEN_194; // @[cacheLookupUnit.scala 298:37 305:26]
  wire [31:0] _GEN_236 = _T_18 ? _GEN_194 : _GEN_215; // @[cacheLookupUnit.scala 296:49]
  wire [31:0] _GEN_257 = isLRReadWire | isAtmoicReadWire ? _GEN_236 : _GEN_194; // @[cacheLookupUnit.scala 295:43]
  wire [31:0] _GEN_281 = isReplayValidWire & isDataMissWire ? readBuffer_cacheLine_cacheLine[255:224] : _GEN_257; // @[cacheLookupUnit.scala 317:55 324:26]
  wire [31:0] _GEN_302 = ~isPermissionMiss & _isPermissionMiss_T ? _GEN_257 : _GEN_281; // @[cacheLookupUnit.scala 314:49]
  wire [31:0] writeChunks_7 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_302 : _GEN_257; // @[cacheLookupUnit.scala 313:61]
  wire [31:0] _GEN_111 = 4'h7 == _doubleWordWrite_T_1 ? writeChunks_7 : _GEN_110; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_153 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[287:256] : cacheLineChoosen[287:256]; // @[cacheLookupUnit.scala 284:37 291:26 262:30]
  wire [31:0] _GEN_174 = _isPermissionMiss_T ? cacheLineChoosen[287:256] : _GEN_153; // @[cacheLookupUnit.scala 282:28 262:30]
  wire [31:0] _GEN_195 = isReadWire ? _GEN_174 : cacheLineChoosen[287:256]; // @[cacheLookupUnit.scala 281:21 262:30]
  wire [31:0] _GEN_216 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[287:256] : _GEN_195; // @[cacheLookupUnit.scala 298:37 305:26]
  wire [31:0] _GEN_237 = _T_18 ? _GEN_195 : _GEN_216; // @[cacheLookupUnit.scala 296:49]
  wire [31:0] _GEN_258 = isLRReadWire | isAtmoicReadWire ? _GEN_237 : _GEN_195; // @[cacheLookupUnit.scala 295:43]
  wire [31:0] _GEN_282 = isReplayValidWire & isDataMissWire ? readBuffer_cacheLine_cacheLine[287:256] : _GEN_258; // @[cacheLookupUnit.scala 317:55 324:26]
  wire [31:0] _GEN_303 = ~isPermissionMiss & _isPermissionMiss_T ? _GEN_258 : _GEN_282; // @[cacheLookupUnit.scala 314:49]
  wire [31:0] writeChunks_8 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_303 : _GEN_258; // @[cacheLookupUnit.scala 313:61]
  wire [31:0] _GEN_112 = 4'h8 == _doubleWordWrite_T_1 ? writeChunks_8 : _GEN_111; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_154 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[319:288] : cacheLineChoosen[319:288]; // @[cacheLookupUnit.scala 284:37 291:26 262:30]
  wire [31:0] _GEN_175 = _isPermissionMiss_T ? cacheLineChoosen[319:288] : _GEN_154; // @[cacheLookupUnit.scala 282:28 262:30]
  wire [31:0] _GEN_196 = isReadWire ? _GEN_175 : cacheLineChoosen[319:288]; // @[cacheLookupUnit.scala 281:21 262:30]
  wire [31:0] _GEN_217 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[319:288] : _GEN_196; // @[cacheLookupUnit.scala 298:37 305:26]
  wire [31:0] _GEN_238 = _T_18 ? _GEN_196 : _GEN_217; // @[cacheLookupUnit.scala 296:49]
  wire [31:0] _GEN_259 = isLRReadWire | isAtmoicReadWire ? _GEN_238 : _GEN_196; // @[cacheLookupUnit.scala 295:43]
  wire [31:0] _GEN_283 = isReplayValidWire & isDataMissWire ? readBuffer_cacheLine_cacheLine[319:288] : _GEN_259; // @[cacheLookupUnit.scala 317:55 324:26]
  wire [31:0] _GEN_304 = ~isPermissionMiss & _isPermissionMiss_T ? _GEN_259 : _GEN_283; // @[cacheLookupUnit.scala 314:49]
  wire [31:0] writeChunks_9 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_304 : _GEN_259; // @[cacheLookupUnit.scala 313:61]
  wire [31:0] _GEN_113 = 4'h9 == _doubleWordWrite_T_1 ? writeChunks_9 : _GEN_112; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_155 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[351:320] : cacheLineChoosen[351:320]; // @[cacheLookupUnit.scala 284:37 291:26 262:30]
  wire [31:0] _GEN_176 = _isPermissionMiss_T ? cacheLineChoosen[351:320] : _GEN_155; // @[cacheLookupUnit.scala 282:28 262:30]
  wire [31:0] _GEN_197 = isReadWire ? _GEN_176 : cacheLineChoosen[351:320]; // @[cacheLookupUnit.scala 281:21 262:30]
  wire [31:0] _GEN_218 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[351:320] : _GEN_197; // @[cacheLookupUnit.scala 298:37 305:26]
  wire [31:0] _GEN_239 = _T_18 ? _GEN_197 : _GEN_218; // @[cacheLookupUnit.scala 296:49]
  wire [31:0] _GEN_260 = isLRReadWire | isAtmoicReadWire ? _GEN_239 : _GEN_197; // @[cacheLookupUnit.scala 295:43]
  wire [31:0] _GEN_284 = isReplayValidWire & isDataMissWire ? readBuffer_cacheLine_cacheLine[351:320] : _GEN_260; // @[cacheLookupUnit.scala 317:55 324:26]
  wire [31:0] _GEN_305 = ~isPermissionMiss & _isPermissionMiss_T ? _GEN_260 : _GEN_284; // @[cacheLookupUnit.scala 314:49]
  wire [31:0] writeChunks_10 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_305 : _GEN_260; // @[cacheLookupUnit.scala 313:61]
  wire [31:0] _GEN_114 = 4'ha == _doubleWordWrite_T_1 ? writeChunks_10 : _GEN_113; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_156 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[383:352] : cacheLineChoosen[383:352]; // @[cacheLookupUnit.scala 284:37 291:26 262:30]
  wire [31:0] _GEN_177 = _isPermissionMiss_T ? cacheLineChoosen[383:352] : _GEN_156; // @[cacheLookupUnit.scala 282:28 262:30]
  wire [31:0] _GEN_198 = isReadWire ? _GEN_177 : cacheLineChoosen[383:352]; // @[cacheLookupUnit.scala 281:21 262:30]
  wire [31:0] _GEN_219 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[383:352] : _GEN_198; // @[cacheLookupUnit.scala 298:37 305:26]
  wire [31:0] _GEN_240 = _T_18 ? _GEN_198 : _GEN_219; // @[cacheLookupUnit.scala 296:49]
  wire [31:0] _GEN_261 = isLRReadWire | isAtmoicReadWire ? _GEN_240 : _GEN_198; // @[cacheLookupUnit.scala 295:43]
  wire [31:0] _GEN_285 = isReplayValidWire & isDataMissWire ? readBuffer_cacheLine_cacheLine[383:352] : _GEN_261; // @[cacheLookupUnit.scala 317:55 324:26]
  wire [31:0] _GEN_306 = ~isPermissionMiss & _isPermissionMiss_T ? _GEN_261 : _GEN_285; // @[cacheLookupUnit.scala 314:49]
  wire [31:0] writeChunks_11 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_306 : _GEN_261; // @[cacheLookupUnit.scala 313:61]
  wire [31:0] _GEN_115 = 4'hb == _doubleWordWrite_T_1 ? writeChunks_11 : _GEN_114; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_157 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[415:384] : cacheLineChoosen[415:384]; // @[cacheLookupUnit.scala 284:37 291:26 262:30]
  wire [31:0] _GEN_178 = _isPermissionMiss_T ? cacheLineChoosen[415:384] : _GEN_157; // @[cacheLookupUnit.scala 282:28 262:30]
  wire [31:0] _GEN_199 = isReadWire ? _GEN_178 : cacheLineChoosen[415:384]; // @[cacheLookupUnit.scala 281:21 262:30]
  wire [31:0] _GEN_220 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[415:384] : _GEN_199; // @[cacheLookupUnit.scala 298:37 305:26]
  wire [31:0] _GEN_241 = _T_18 ? _GEN_199 : _GEN_220; // @[cacheLookupUnit.scala 296:49]
  wire [31:0] _GEN_262 = isLRReadWire | isAtmoicReadWire ? _GEN_241 : _GEN_199; // @[cacheLookupUnit.scala 295:43]
  wire [31:0] _GEN_286 = isReplayValidWire & isDataMissWire ? readBuffer_cacheLine_cacheLine[415:384] : _GEN_262; // @[cacheLookupUnit.scala 317:55 324:26]
  wire [31:0] _GEN_307 = ~isPermissionMiss & _isPermissionMiss_T ? _GEN_262 : _GEN_286; // @[cacheLookupUnit.scala 314:49]
  wire [31:0] writeChunks_12 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_307 : _GEN_262; // @[cacheLookupUnit.scala 313:61]
  wire [31:0] _GEN_116 = 4'hc == _doubleWordWrite_T_1 ? writeChunks_12 : _GEN_115; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_158 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[447:416] : cacheLineChoosen[447:416]; // @[cacheLookupUnit.scala 284:37 291:26 262:30]
  wire [31:0] _GEN_179 = _isPermissionMiss_T ? cacheLineChoosen[447:416] : _GEN_158; // @[cacheLookupUnit.scala 282:28 262:30]
  wire [31:0] _GEN_200 = isReadWire ? _GEN_179 : cacheLineChoosen[447:416]; // @[cacheLookupUnit.scala 281:21 262:30]
  wire [31:0] _GEN_221 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[447:416] : _GEN_200; // @[cacheLookupUnit.scala 298:37 305:26]
  wire [31:0] _GEN_242 = _T_18 ? _GEN_200 : _GEN_221; // @[cacheLookupUnit.scala 296:49]
  wire [31:0] _GEN_263 = isLRReadWire | isAtmoicReadWire ? _GEN_242 : _GEN_200; // @[cacheLookupUnit.scala 295:43]
  wire [31:0] _GEN_287 = isReplayValidWire & isDataMissWire ? readBuffer_cacheLine_cacheLine[447:416] : _GEN_263; // @[cacheLookupUnit.scala 317:55 324:26]
  wire [31:0] _GEN_308 = ~isPermissionMiss & _isPermissionMiss_T ? _GEN_263 : _GEN_287; // @[cacheLookupUnit.scala 314:49]
  wire [31:0] writeChunks_13 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_308 : _GEN_263; // @[cacheLookupUnit.scala 313:61]
  wire [31:0] _GEN_117 = 4'hd == _doubleWordWrite_T_1 ? writeChunks_13 : _GEN_116; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_159 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[479:448] : cacheLineChoosen[479:448]; // @[cacheLookupUnit.scala 284:37 291:26 262:30]
  wire [31:0] _GEN_180 = _isPermissionMiss_T ? cacheLineChoosen[479:448] : _GEN_159; // @[cacheLookupUnit.scala 282:28 262:30]
  wire [31:0] _GEN_201 = isReadWire ? _GEN_180 : cacheLineChoosen[479:448]; // @[cacheLookupUnit.scala 281:21 262:30]
  wire [31:0] _GEN_222 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[479:448] : _GEN_201; // @[cacheLookupUnit.scala 298:37 305:26]
  wire [31:0] _GEN_243 = _T_18 ? _GEN_201 : _GEN_222; // @[cacheLookupUnit.scala 296:49]
  wire [31:0] _GEN_264 = isLRReadWire | isAtmoicReadWire ? _GEN_243 : _GEN_201; // @[cacheLookupUnit.scala 295:43]
  wire [31:0] _GEN_288 = isReplayValidWire & isDataMissWire ? readBuffer_cacheLine_cacheLine[479:448] : _GEN_264; // @[cacheLookupUnit.scala 317:55 324:26]
  wire [31:0] _GEN_309 = ~isPermissionMiss & _isPermissionMiss_T ? _GEN_264 : _GEN_288; // @[cacheLookupUnit.scala 314:49]
  wire [31:0] writeChunks_14 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_309 : _GEN_264; // @[cacheLookupUnit.scala 313:61]
  wire [31:0] _GEN_118 = 4'he == _doubleWordWrite_T_1 ? writeChunks_14 : _GEN_117; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_160 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[511:480] : cacheLineChoosen[511:480]; // @[cacheLookupUnit.scala 284:37 291:26 262:30]
  wire [31:0] _GEN_181 = _isPermissionMiss_T ? cacheLineChoosen[511:480] : _GEN_160; // @[cacheLookupUnit.scala 282:28 262:30]
  wire [31:0] _GEN_202 = isReadWire ? _GEN_181 : cacheLineChoosen[511:480]; // @[cacheLookupUnit.scala 281:21 262:30]
  wire [31:0] _GEN_223 = isReplayValidWire ? readBuffer_cacheLine_cacheLine[511:480] : _GEN_202; // @[cacheLookupUnit.scala 298:37 305:26]
  wire [31:0] _GEN_244 = _T_18 ? _GEN_202 : _GEN_223; // @[cacheLookupUnit.scala 296:49]
  wire [31:0] _GEN_265 = isLRReadWire | isAtmoicReadWire ? _GEN_244 : _GEN_202; // @[cacheLookupUnit.scala 295:43]
  wire [31:0] _GEN_289 = isReplayValidWire & isDataMissWire ? readBuffer_cacheLine_cacheLine[511:480] : _GEN_265; // @[cacheLookupUnit.scala 317:55 324:26]
  wire [31:0] _GEN_310 = ~isPermissionMiss & _isPermissionMiss_T ? _GEN_265 : _GEN_289; // @[cacheLookupUnit.scala 314:49]
  wire [31:0] writeChunks_15 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_310 : _GEN_265; // @[cacheLookupUnit.scala 313:61]
  wire [31:0] _GEN_119 = 4'hf == _doubleWordWrite_T_1 ? writeChunks_15 : _GEN_118; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_121 = 4'h1 == _doubleWordWrite_T_3 ? writeChunks_1 : writeChunks_0; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_122 = 4'h2 == _doubleWordWrite_T_3 ? writeChunks_2 : _GEN_121; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_123 = 4'h3 == _doubleWordWrite_T_3 ? writeChunks_3 : _GEN_122; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_124 = 4'h4 == _doubleWordWrite_T_3 ? writeChunks_4 : _GEN_123; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_125 = 4'h5 == _doubleWordWrite_T_3 ? writeChunks_5 : _GEN_124; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_126 = 4'h6 == _doubleWordWrite_T_3 ? writeChunks_6 : _GEN_125; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_127 = 4'h7 == _doubleWordWrite_T_3 ? writeChunks_7 : _GEN_126; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_128 = 4'h8 == _doubleWordWrite_T_3 ? writeChunks_8 : _GEN_127; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_129 = 4'h9 == _doubleWordWrite_T_3 ? writeChunks_9 : _GEN_128; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_130 = 4'ha == _doubleWordWrite_T_3 ? writeChunks_10 : _GEN_129; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_131 = 4'hb == _doubleWordWrite_T_3 ? writeChunks_11 : _GEN_130; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_132 = 4'hc == _doubleWordWrite_T_3 ? writeChunks_12 : _GEN_131; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_133 = 4'hd == _doubleWordWrite_T_3 ? writeChunks_13 : _GEN_132; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_134 = 4'he == _doubleWordWrite_T_3 ? writeChunks_14 : _GEN_133; // @[Cat.scala 33:{92,92}]
  wire [31:0] _GEN_135 = 4'hf == _doubleWordWrite_T_3 ? writeChunks_15 : _GEN_134; // @[Cat.scala 33:{92,92}]
  wire [63:0] doubleWordWrite = {_GEN_119,_GEN_135}; // @[Cat.scala 33:92]
  wire  PLRUSetWire_0 = tagChunks_0[22]; // @[cacheLookupUnit.scala 273:71]
  wire  PLRUSetWire_1 = tagChunks_1[22]; // @[cacheLookupUnit.scala 273:71]
  wire  PLRUSetWire_2 = tagChunks_2[22]; // @[cacheLookupUnit.scala 273:71]
  wire  PLRUSetWire_3 = tagChunks_3[22]; // @[cacheLookupUnit.scala 273:71]
  wire  flippedPLRUSetWire_0 = ~PLRUSetWire_0; // @[cacheLookupUnit.scala 274:73]
  wire  flippedPLRUSetWire_1 = ~PLRUSetWire_1; // @[cacheLookupUnit.scala 274:73]
  wire  flippedPLRUSetWire_2 = ~PLRUSetWire_2; // @[cacheLookupUnit.scala 274:73]
  wire [1:0] _replacingset_T = flippedPLRUSetWire_2 ? 2'h2 : 2'h3; // @[Mux.scala 47:70]
  wire [1:0] _replacingset_T_1 = flippedPLRUSetWire_1 ? 2'h1 : _replacingset_T; // @[Mux.scala 47:70]
  wire [1:0] replacingset = flippedPLRUSetWire_0 ? 2'h0 : _replacingset_T_1; // @[Mux.scala 47:70]
  wire [22:0] _GEN_137 = 2'h1 == replacingset ? tagChunks_1 : tagChunks_0; // @[cacheLookupUnit.scala 277:{64,64}]
  wire [22:0] _GEN_138 = 2'h2 == replacingset ? tagChunks_2 : _GEN_137; // @[cacheLookupUnit.scala 277:{64,64}]
  wire [22:0] _GEN_139 = 2'h3 == replacingset ? tagChunks_3 : _GEN_138; // @[cacheLookupUnit.scala 277:{64,64}]
  wire  isUpdateValidWire = _GEN_139[19]; // @[cacheLookupUnit.scala 277:64]
  wire  isUpdateDirtyWire = _GEN_139[20]; // @[cacheLookupUnit.scala 278:64]
  wire  _newPLRUBitWire_T_5 = PLRUSetWire_0 & PLRUSetWire_1 & PLRUSetWire_2 & PLRUSetWire_3; // @[cacheLookupUnit.scala 283:52]
  wire  _newPLRUBitWire_T_6 = PLRUSetWire_0 & PLRUSetWire_1 & PLRUSetWire_2 & PLRUSetWire_3 ? 1'h0 : 1'h1; // @[cacheLookupUnit.scala 283:30]
  wire  _GEN_140 = isReplayValidWire ? _newPLRUBitWire_T_6 : _GEN_67[22]; // @[cacheLookupUnit.scala 284:37 285:24]
  wire  _GEN_141 = isReplayValidWire | validBitWire; // @[cacheLookupUnit.scala 284:37 286:25]
  wire  _GEN_142 = isReplayValidWire ? readBuffer_cacheLine_response[1] : shareBitWire; // @[cacheLookupUnit.scala 284:37 287:25]
  wire  _GEN_143 = isReplayValidWire ? readBuffer_cacheLine_response[0] : dirtyBitWire; // @[cacheLookupUnit.scala 284:37 288:25]
  wire [18:0] _GEN_144 = isReplayValidWire ? readBuffer_address[31:13] : _GEN_67[18:0]; // @[cacheLookupUnit.scala 284:37 289:21]
  wire  _GEN_161 = _isPermissionMiss_T ? _newPLRUBitWire_T_6 : _GEN_140; // @[cacheLookupUnit.scala 282:28 283:24]
  wire  _GEN_162 = _isPermissionMiss_T ? validBitWire : _GEN_141; // @[cacheLookupUnit.scala 282:28]
  wire  _GEN_163 = _isPermissionMiss_T ? shareBitWire : _GEN_142; // @[cacheLookupUnit.scala 282:28]
  wire  _GEN_164 = _isPermissionMiss_T ? dirtyBitWire : _GEN_143; // @[cacheLookupUnit.scala 282:28]
  wire [18:0] _GEN_165 = _isPermissionMiss_T ? _GEN_67[18:0] : _GEN_144; // @[cacheLookupUnit.scala 282:28]
  wire  _GEN_182 = isReadWire ? _GEN_161 : _GEN_67[22]; // @[cacheLookupUnit.scala 281:21]
  wire  _GEN_183 = isReadWire ? _GEN_162 : validBitWire; // @[cacheLookupUnit.scala 281:21]
  wire  _GEN_184 = isReadWire ? _GEN_163 : shareBitWire; // @[cacheLookupUnit.scala 281:21]
  wire  _GEN_185 = isReadWire ? _GEN_164 : dirtyBitWire; // @[cacheLookupUnit.scala 281:21]
  wire [18:0] _GEN_186 = isReadWire ? _GEN_165 : _GEN_67[18:0]; // @[cacheLookupUnit.scala 281:21]
  wire  _GEN_203 = isReplayValidWire ? _newPLRUBitWire_T_6 : _GEN_182; // @[cacheLookupUnit.scala 298:37 299:24]
  wire  _GEN_204 = isReplayValidWire | _GEN_183; // @[cacheLookupUnit.scala 298:37 300:25]
  wire  _GEN_205 = isReplayValidWire ? readBuffer_cacheLine_response[1] : _GEN_184; // @[cacheLookupUnit.scala 298:37 301:25]
  wire  _GEN_206 = isReplayValidWire ? readBuffer_cacheLine_response[0] : _GEN_185; // @[cacheLookupUnit.scala 298:37 302:25]
  wire [18:0] _GEN_207 = isReplayValidWire ? readBuffer_address[31:13] : _GEN_186; // @[cacheLookupUnit.scala 298:37 303:21]
  wire  _GEN_224 = _T_18 ? _newPLRUBitWire_T_6 : _GEN_203; // @[cacheLookupUnit.scala 296:49 297:24]
  wire  _GEN_225 = _T_18 ? _GEN_183 : _GEN_204; // @[cacheLookupUnit.scala 296:49]
  wire  _GEN_226 = _T_18 ? _GEN_184 : _GEN_205; // @[cacheLookupUnit.scala 296:49]
  wire  _GEN_227 = _T_18 ? _GEN_185 : _GEN_206; // @[cacheLookupUnit.scala 296:49]
  wire [18:0] _GEN_228 = _T_18 ? _GEN_186 : _GEN_207; // @[cacheLookupUnit.scala 296:49]
  wire  _GEN_245 = isLRReadWire | isAtmoicReadWire ? _GEN_224 : _GEN_182; // @[cacheLookupUnit.scala 295:43]
  wire  _GEN_246 = isLRReadWire | isAtmoicReadWire ? _GEN_225 : _GEN_183; // @[cacheLookupUnit.scala 295:43]
  wire  _GEN_247 = isLRReadWire | isAtmoicReadWire ? _GEN_226 : _GEN_184; // @[cacheLookupUnit.scala 295:43]
  wire  _GEN_248 = isLRReadWire | isAtmoicReadWire ? _GEN_227 : _GEN_185; // @[cacheLookupUnit.scala 295:43]
  wire [18:0] _GEN_249 = isLRReadWire | isAtmoicReadWire ? _GEN_228 : _GEN_186; // @[cacheLookupUnit.scala 295:43]
  wire  _GEN_266 = isReplayValidWire & isPermissionMiss | _GEN_246; // @[cacheLookupUnit.scala 327:57 328:25]
  wire  _GEN_267 = isReplayValidWire & isPermissionMiss ? readBuffer_cacheLine_response[1] : _GEN_247; // @[cacheLookupUnit.scala 327:57 329:25]
  wire [18:0] _GEN_268 = isReplayValidWire & isPermissionMiss ? readBuffer_address[31:13] : _GEN_249; // @[cacheLookupUnit.scala 327:57 330:21]
  wire  _GEN_269 = isReplayValidWire & isDataMissWire | _GEN_266; // @[cacheLookupUnit.scala 317:55 318:25]
  wire  _GEN_270 = isReplayValidWire & isDataMissWire | _GEN_248; // @[cacheLookupUnit.scala 317:55 319:25]
  wire  _GEN_271 = isReplayValidWire & isDataMissWire ? readBuffer_cacheLine_response[1] : _GEN_267; // @[cacheLookupUnit.scala 317:55 320:25]
  wire  _GEN_272 = isReplayValidWire & isDataMissWire ? _newPLRUBitWire_T_6 : _GEN_245; // @[cacheLookupUnit.scala 317:55 321:24]
  wire [18:0] _GEN_273 = isReplayValidWire & isDataMissWire ? readBuffer_address[31:13] : _GEN_268; // @[cacheLookupUnit.scala 317:55 322:21]
  wire  _GEN_290 = ~isPermissionMiss & _isPermissionMiss_T | _GEN_270; // @[cacheLookupUnit.scala 314:49 315:25]
  wire  _GEN_291 = ~isPermissionMiss & _isPermissionMiss_T ? _newPLRUBitWire_T_6 : _GEN_272; // @[cacheLookupUnit.scala 314:49 316:24]
  wire  _GEN_292 = ~isPermissionMiss & _isPermissionMiss_T ? _GEN_246 : _GEN_269; // @[cacheLookupUnit.scala 314:49]
  wire  _GEN_293 = ~isPermissionMiss & _isPermissionMiss_T ? _GEN_247 : _GEN_271; // @[cacheLookupUnit.scala 314:49]
  wire [18:0] _GEN_294 = ~isPermissionMiss & _isPermissionMiss_T ? _GEN_249 : _GEN_273; // @[cacheLookupUnit.scala 314:49]
  wire  _T_24 = 5'h1 == readBuffer_core_instruction[31:27]; // @[cacheLookupUnit.scala 334:53]
  wire  _T_25 = 5'h0 == readBuffer_core_instruction[31:27]; // @[cacheLookupUnit.scala 334:53]
  wire [31:0] _GEN_312 = 4'h1 == readBuffer_address[5:2] ? writeChunks_1 : writeChunks_0; // @[cacheLookupUnit.scala 336:{50,50}]
  wire [31:0] _GEN_313 = 4'h2 == readBuffer_address[5:2] ? writeChunks_2 : _GEN_312; // @[cacheLookupUnit.scala 336:{50,50}]
  wire [31:0] _GEN_314 = 4'h3 == readBuffer_address[5:2] ? writeChunks_3 : _GEN_313; // @[cacheLookupUnit.scala 336:{50,50}]
  wire [31:0] _GEN_315 = 4'h4 == readBuffer_address[5:2] ? writeChunks_4 : _GEN_314; // @[cacheLookupUnit.scala 336:{50,50}]
  wire [31:0] _GEN_316 = 4'h5 == readBuffer_address[5:2] ? writeChunks_5 : _GEN_315; // @[cacheLookupUnit.scala 336:{50,50}]
  wire [31:0] _GEN_317 = 4'h6 == readBuffer_address[5:2] ? writeChunks_6 : _GEN_316; // @[cacheLookupUnit.scala 336:{50,50}]
  wire [31:0] _GEN_318 = 4'h7 == readBuffer_address[5:2] ? writeChunks_7 : _GEN_317; // @[cacheLookupUnit.scala 336:{50,50}]
  wire [31:0] _GEN_319 = 4'h8 == readBuffer_address[5:2] ? writeChunks_8 : _GEN_318; // @[cacheLookupUnit.scala 336:{50,50}]
  wire [31:0] _GEN_320 = 4'h9 == readBuffer_address[5:2] ? writeChunks_9 : _GEN_319; // @[cacheLookupUnit.scala 336:{50,50}]
  wire [31:0] _GEN_321 = 4'ha == readBuffer_address[5:2] ? writeChunks_10 : _GEN_320; // @[cacheLookupUnit.scala 336:{50,50}]
  wire [31:0] _GEN_322 = 4'hb == readBuffer_address[5:2] ? writeChunks_11 : _GEN_321; // @[cacheLookupUnit.scala 336:{50,50}]
  wire [31:0] _GEN_323 = 4'hc == readBuffer_address[5:2] ? writeChunks_12 : _GEN_322; // @[cacheLookupUnit.scala 336:{50,50}]
  wire [31:0] _GEN_324 = 4'hd == readBuffer_address[5:2] ? writeChunks_13 : _GEN_323; // @[cacheLookupUnit.scala 336:{50,50}]
  wire [31:0] _GEN_325 = 4'he == readBuffer_address[5:2] ? writeChunks_14 : _GEN_324; // @[cacheLookupUnit.scala 336:{50,50}]
  wire [31:0] _GEN_326 = 4'hf == readBuffer_address[5:2] ? writeChunks_15 : _GEN_325; // @[cacheLookupUnit.scala 336:{50,50}]
  wire [31:0] _result32_T_3 = _GEN_326 + readBuffer_writeData_data[31:0]; // @[cacheLookupUnit.scala 336:50]
  wire  _T_26 = 5'h4 == readBuffer_core_instruction[31:27]; // @[cacheLookupUnit.scala 334:53]
  wire [31:0] _result32_T_5 = _GEN_326 ^ readBuffer_writeData_data[31:0]; // @[cacheLookupUnit.scala 337:50]
  wire  _T_27 = 5'hc == readBuffer_core_instruction[31:27]; // @[cacheLookupUnit.scala 334:53]
  wire [31:0] _result32_T_7 = _GEN_326 & readBuffer_writeData_data[31:0]; // @[cacheLookupUnit.scala 338:50]
  wire  _T_28 = 5'h8 == readBuffer_core_instruction[31:27]; // @[cacheLookupUnit.scala 334:53]
  wire [31:0] _result32_T_9 = _GEN_326 | readBuffer_writeData_data[31:0]; // @[cacheLookupUnit.scala 339:50]
  wire  _T_29 = 5'h10 == readBuffer_core_instruction[31:27]; // @[cacheLookupUnit.scala 334:53]
  wire [31:0] _result32_T_10 = 4'hf == readBuffer_address[5:2] ? writeChunks_15 : _GEN_325; // @[cacheLookupUnit.scala 340:54]
  wire [31:0] _result32_T_12 = readBuffer_writeData_data[31:0]; // @[cacheLookupUnit.scala 340:95]
  wire [31:0] _result32_T_15 = $signed(_result32_T_10) < $signed(_result32_T_12) ? _GEN_326 : readBuffer_writeData_data[
    31:0]; // @[cacheLookupUnit.scala 340:43]
  wire  _T_30 = 5'h14 == readBuffer_core_instruction[31:27]; // @[cacheLookupUnit.scala 334:53]
  wire [31:0] _result32_T_21 = $signed(_result32_T_10) > $signed(_result32_T_12) ? _GEN_326 : readBuffer_writeData_data[
    31:0]; // @[cacheLookupUnit.scala 341:43]
  wire  _T_31 = 5'h18 == readBuffer_core_instruction[31:27]; // @[cacheLookupUnit.scala 334:53]
  wire [31:0] _result32_T_25 = _GEN_326 < readBuffer_writeData_data[31:0] ? _GEN_326 : readBuffer_writeData_data[31:0]; // @[cacheLookupUnit.scala 342:43]
  wire  _T_32 = 5'h1c == readBuffer_core_instruction[31:27]; // @[cacheLookupUnit.scala 334:53]
  wire [31:0] _result32_T_29 = _GEN_326 > readBuffer_writeData_data[31:0] ? _GEN_326 : readBuffer_writeData_data[31:0]; // @[cacheLookupUnit.scala 343:43]
  wire [31:0] _GEN_327 = 5'h1c == readBuffer_core_instruction[31:27] ? _result32_T_29 : 32'h0; // @[cacheLookupUnit.scala 334:53 343:37]
  wire [31:0] _GEN_328 = 5'h18 == readBuffer_core_instruction[31:27] ? _result32_T_25 : _GEN_327; // @[cacheLookupUnit.scala 334:53 342:37]
  wire [31:0] _GEN_329 = 5'h14 == readBuffer_core_instruction[31:27] ? _result32_T_21 : _GEN_328; // @[cacheLookupUnit.scala 334:53 341:37]
  wire [31:0] _GEN_330 = 5'h10 == readBuffer_core_instruction[31:27] ? _result32_T_15 : _GEN_329; // @[cacheLookupUnit.scala 334:53 340:37]
  wire [31:0] _GEN_331 = 5'h8 == readBuffer_core_instruction[31:27] ? _result32_T_9 : _GEN_330; // @[cacheLookupUnit.scala 334:53 339:37]
  wire [31:0] _GEN_332 = 5'hc == readBuffer_core_instruction[31:27] ? _result32_T_7 : _GEN_331; // @[cacheLookupUnit.scala 334:53 338:37]
  wire [31:0] _GEN_333 = 5'h4 == readBuffer_core_instruction[31:27] ? _result32_T_5 : _GEN_332; // @[cacheLookupUnit.scala 334:53 337:37]
  wire [31:0] _GEN_334 = 5'h0 == readBuffer_core_instruction[31:27] ? _result32_T_3 : _GEN_333; // @[cacheLookupUnit.scala 334:53 336:37]
  wire [31:0] _GEN_335 = 5'h1 == readBuffer_core_instruction[31:27] ? readBuffer_writeData_data[31:0] : _GEN_334; // @[cacheLookupUnit.scala 334:53 335:37]
  wire [31:0] _GEN_352 = readBuffer_core_instruction[14:12] == 3'h2 ? _GEN_335 : 32'h0; // @[cacheLookupUnit.scala 333:62]
  wire [31:0] _GEN_547 = isAtmoicWriteWire ? _GEN_352 : 32'h0; // @[cacheLookupUnit.scala 332:30]
  wire [31:0] result32 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_547 : 32'h0; // @[cacheLookupUnit.scala 313:61]
  wire [31:0] _GEN_336 = 4'h0 == readBuffer_address[5:2] ? result32 : cacheLineChoosen[31:0]; // @[cacheLookupUnit.scala 265:33 345:{51,51}]
  wire [31:0] _GEN_337 = 4'h1 == readBuffer_address[5:2] ? result32 : cacheLineChoosen[63:32]; // @[cacheLookupUnit.scala 265:33 345:{51,51}]
  wire [31:0] _GEN_338 = 4'h2 == readBuffer_address[5:2] ? result32 : cacheLineChoosen[95:64]; // @[cacheLookupUnit.scala 265:33 345:{51,51}]
  wire [31:0] _GEN_339 = 4'h3 == readBuffer_address[5:2] ? result32 : cacheLineChoosen[127:96]; // @[cacheLookupUnit.scala 265:33 345:{51,51}]
  wire [31:0] _GEN_340 = 4'h4 == readBuffer_address[5:2] ? result32 : cacheLineChoosen[159:128]; // @[cacheLookupUnit.scala 265:33 345:{51,51}]
  wire [31:0] _GEN_341 = 4'h5 == readBuffer_address[5:2] ? result32 : cacheLineChoosen[191:160]; // @[cacheLookupUnit.scala 265:33 345:{51,51}]
  wire [31:0] _GEN_342 = 4'h6 == readBuffer_address[5:2] ? result32 : cacheLineChoosen[223:192]; // @[cacheLookupUnit.scala 265:33 345:{51,51}]
  wire [31:0] _GEN_343 = 4'h7 == readBuffer_address[5:2] ? result32 : cacheLineChoosen[255:224]; // @[cacheLookupUnit.scala 265:33 345:{51,51}]
  wire [31:0] _GEN_344 = 4'h8 == readBuffer_address[5:2] ? result32 : cacheLineChoosen[287:256]; // @[cacheLookupUnit.scala 265:33 345:{51,51}]
  wire [31:0] _GEN_345 = 4'h9 == readBuffer_address[5:2] ? result32 : cacheLineChoosen[319:288]; // @[cacheLookupUnit.scala 265:33 345:{51,51}]
  wire [31:0] _GEN_346 = 4'ha == readBuffer_address[5:2] ? result32 : cacheLineChoosen[351:320]; // @[cacheLookupUnit.scala 265:33 345:{51,51}]
  wire [31:0] _GEN_347 = 4'hb == readBuffer_address[5:2] ? result32 : cacheLineChoosen[383:352]; // @[cacheLookupUnit.scala 265:33 345:{51,51}]
  wire [31:0] _GEN_348 = 4'hc == readBuffer_address[5:2] ? result32 : cacheLineChoosen[415:384]; // @[cacheLookupUnit.scala 265:33 345:{51,51}]
  wire [31:0] _GEN_349 = 4'hd == readBuffer_address[5:2] ? result32 : cacheLineChoosen[447:416]; // @[cacheLookupUnit.scala 265:33 345:{51,51}]
  wire [31:0] _GEN_350 = 4'he == readBuffer_address[5:2] ? result32 : cacheLineChoosen[479:448]; // @[cacheLookupUnit.scala 265:33 345:{51,51}]
  wire [31:0] _GEN_351 = 4'hf == readBuffer_address[5:2] ? result32 : cacheLineChoosen[511:480]; // @[cacheLookupUnit.scala 265:33 345:{51,51}]
  wire [31:0] _GEN_353 = readBuffer_core_instruction[14:12] == 3'h2 ? _GEN_336 : cacheLineChoosen[31:0]; // @[cacheLookupUnit.scala 265:33 333:62]
  wire [31:0] _GEN_354 = readBuffer_core_instruction[14:12] == 3'h2 ? _GEN_337 : cacheLineChoosen[63:32]; // @[cacheLookupUnit.scala 265:33 333:62]
  wire [31:0] _GEN_355 = readBuffer_core_instruction[14:12] == 3'h2 ? _GEN_338 : cacheLineChoosen[95:64]; // @[cacheLookupUnit.scala 265:33 333:62]
  wire [31:0] _GEN_356 = readBuffer_core_instruction[14:12] == 3'h2 ? _GEN_339 : cacheLineChoosen[127:96]; // @[cacheLookupUnit.scala 265:33 333:62]
  wire [31:0] _GEN_357 = readBuffer_core_instruction[14:12] == 3'h2 ? _GEN_340 : cacheLineChoosen[159:128]; // @[cacheLookupUnit.scala 265:33 333:62]
  wire [31:0] _GEN_358 = readBuffer_core_instruction[14:12] == 3'h2 ? _GEN_341 : cacheLineChoosen[191:160]; // @[cacheLookupUnit.scala 265:33 333:62]
  wire [31:0] _GEN_359 = readBuffer_core_instruction[14:12] == 3'h2 ? _GEN_342 : cacheLineChoosen[223:192]; // @[cacheLookupUnit.scala 265:33 333:62]
  wire [31:0] _GEN_360 = readBuffer_core_instruction[14:12] == 3'h2 ? _GEN_343 : cacheLineChoosen[255:224]; // @[cacheLookupUnit.scala 265:33 333:62]
  wire [31:0] _GEN_361 = readBuffer_core_instruction[14:12] == 3'h2 ? _GEN_344 : cacheLineChoosen[287:256]; // @[cacheLookupUnit.scala 265:33 333:62]
  wire [31:0] _GEN_362 = readBuffer_core_instruction[14:12] == 3'h2 ? _GEN_345 : cacheLineChoosen[319:288]; // @[cacheLookupUnit.scala 265:33 333:62]
  wire [31:0] _GEN_363 = readBuffer_core_instruction[14:12] == 3'h2 ? _GEN_346 : cacheLineChoosen[351:320]; // @[cacheLookupUnit.scala 265:33 333:62]
  wire [31:0] _GEN_364 = readBuffer_core_instruction[14:12] == 3'h2 ? _GEN_347 : cacheLineChoosen[383:352]; // @[cacheLookupUnit.scala 265:33 333:62]
  wire [31:0] _GEN_365 = readBuffer_core_instruction[14:12] == 3'h2 ? _GEN_348 : cacheLineChoosen[415:384]; // @[cacheLookupUnit.scala 265:33 333:62]
  wire [31:0] _GEN_366 = readBuffer_core_instruction[14:12] == 3'h2 ? _GEN_349 : cacheLineChoosen[447:416]; // @[cacheLookupUnit.scala 265:33 333:62]
  wire [31:0] _GEN_367 = readBuffer_core_instruction[14:12] == 3'h2 ? _GEN_350 : cacheLineChoosen[479:448]; // @[cacheLookupUnit.scala 265:33 333:62]
  wire [31:0] _GEN_368 = readBuffer_core_instruction[14:12] == 3'h2 ? _GEN_351 : cacheLineChoosen[511:480]; // @[cacheLookupUnit.scala 265:33 333:62]
  wire [63:0] _result64_T_1 = doubleWordWrite + readBuffer_writeData_data; // @[cacheLookupUnit.scala 350:56]
  wire [63:0] _result64_T_2 = doubleWordWrite ^ readBuffer_writeData_data; // @[cacheLookupUnit.scala 351:56]
  wire [63:0] _result64_T_3 = doubleWordWrite & readBuffer_writeData_data; // @[cacheLookupUnit.scala 352:56]
  wire [63:0] _result64_T_4 = doubleWordWrite | readBuffer_writeData_data; // @[cacheLookupUnit.scala 353:56]
  wire [63:0] _result64_T_5 = {_GEN_119,_GEN_135}; // @[cacheLookupUnit.scala 354:60]
  wire [63:0] _result64_T_8 = $signed(_result64_T_5) < $signed(readBuffer_writeData_data) ? doubleWordWrite :
    readBuffer_writeData_data; // @[cacheLookupUnit.scala 354:43]
  wire [63:0] _result64_T_12 = $signed(_result64_T_5) > $signed(readBuffer_writeData_data) ? doubleWordWrite :
    readBuffer_writeData_data; // @[cacheLookupUnit.scala 355:43]
  wire [63:0] _result64_T_14 = doubleWordWrite < readBuffer_writeData_data ? doubleWordWrite : readBuffer_writeData_data
    ; // @[cacheLookupUnit.scala 356:43]
  wire [63:0] _result64_T_16 = doubleWordWrite > readBuffer_writeData_data ? doubleWordWrite : readBuffer_writeData_data
    ; // @[cacheLookupUnit.scala 357:43]
  wire [63:0] _GEN_369 = _T_32 ? _result64_T_16 : 64'h0; // @[cacheLookupUnit.scala 348:53 357:37]
  wire [63:0] _GEN_370 = _T_31 ? _result64_T_14 : _GEN_369; // @[cacheLookupUnit.scala 348:53 356:37]
  wire [63:0] _GEN_371 = _T_30 ? _result64_T_12 : _GEN_370; // @[cacheLookupUnit.scala 348:53 355:37]
  wire [63:0] _GEN_372 = _T_29 ? _result64_T_8 : _GEN_371; // @[cacheLookupUnit.scala 348:53 354:37]
  wire [63:0] _GEN_373 = _T_28 ? _result64_T_4 : _GEN_372; // @[cacheLookupUnit.scala 348:53 353:37]
  wire [63:0] _GEN_374 = _T_27 ? _result64_T_3 : _GEN_373; // @[cacheLookupUnit.scala 348:53 352:37]
  wire [63:0] _GEN_375 = _T_26 ? _result64_T_2 : _GEN_374; // @[cacheLookupUnit.scala 348:53 351:37]
  wire [63:0] _GEN_376 = _T_25 ? _result64_T_1 : _GEN_375; // @[cacheLookupUnit.scala 348:53 350:37]
  wire [63:0] _GEN_377 = _T_24 ? readBuffer_writeData_data : _GEN_376; // @[cacheLookupUnit.scala 348:53 349:37]
  wire [63:0] _GEN_410 = readBuffer_core_instruction[14:12] == 3'h3 ? _GEN_377 : 64'h0; // @[cacheLookupUnit.scala 347:62]
  wire [63:0] _GEN_564 = isAtmoicWriteWire ? _GEN_410 : 64'h0; // @[cacheLookupUnit.scala 332:30]
  wire [63:0] result64 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_564 : 64'h0; // @[cacheLookupUnit.scala 313:61]
  wire [31:0] _GEN_378 = 4'h0 == readBuffer_address[5:2] ? result64[31:0] : _GEN_353; // @[cacheLookupUnit.scala 359:{51,51}]
  wire [31:0] _GEN_379 = 4'h1 == readBuffer_address[5:2] ? result64[31:0] : _GEN_354; // @[cacheLookupUnit.scala 359:{51,51}]
  wire [31:0] _GEN_380 = 4'h2 == readBuffer_address[5:2] ? result64[31:0] : _GEN_355; // @[cacheLookupUnit.scala 359:{51,51}]
  wire [31:0] _GEN_381 = 4'h3 == readBuffer_address[5:2] ? result64[31:0] : _GEN_356; // @[cacheLookupUnit.scala 359:{51,51}]
  wire [31:0] _GEN_382 = 4'h4 == readBuffer_address[5:2] ? result64[31:0] : _GEN_357; // @[cacheLookupUnit.scala 359:{51,51}]
  wire [31:0] _GEN_383 = 4'h5 == readBuffer_address[5:2] ? result64[31:0] : _GEN_358; // @[cacheLookupUnit.scala 359:{51,51}]
  wire [31:0] _GEN_384 = 4'h6 == readBuffer_address[5:2] ? result64[31:0] : _GEN_359; // @[cacheLookupUnit.scala 359:{51,51}]
  wire [31:0] _GEN_385 = 4'h7 == readBuffer_address[5:2] ? result64[31:0] : _GEN_360; // @[cacheLookupUnit.scala 359:{51,51}]
  wire [31:0] _GEN_386 = 4'h8 == readBuffer_address[5:2] ? result64[31:0] : _GEN_361; // @[cacheLookupUnit.scala 359:{51,51}]
  wire [31:0] _GEN_387 = 4'h9 == readBuffer_address[5:2] ? result64[31:0] : _GEN_362; // @[cacheLookupUnit.scala 359:{51,51}]
  wire [31:0] _GEN_388 = 4'ha == readBuffer_address[5:2] ? result64[31:0] : _GEN_363; // @[cacheLookupUnit.scala 359:{51,51}]
  wire [31:0] _GEN_389 = 4'hb == readBuffer_address[5:2] ? result64[31:0] : _GEN_364; // @[cacheLookupUnit.scala 359:{51,51}]
  wire [31:0] _GEN_390 = 4'hc == readBuffer_address[5:2] ? result64[31:0] : _GEN_365; // @[cacheLookupUnit.scala 359:{51,51}]
  wire [31:0] _GEN_391 = 4'hd == readBuffer_address[5:2] ? result64[31:0] : _GEN_366; // @[cacheLookupUnit.scala 359:{51,51}]
  wire [31:0] _GEN_392 = 4'he == readBuffer_address[5:2] ? result64[31:0] : _GEN_367; // @[cacheLookupUnit.scala 359:{51,51}]
  wire [31:0] _GEN_393 = 4'hf == readBuffer_address[5:2] ? result64[31:0] : _GEN_368; // @[cacheLookupUnit.scala 359:{51,51}]
  wire [3:0] _T_49 = readBuffer_address[5:2] + 4'h1; // @[cacheLookupUnit.scala 360:50]
  wire [31:0] _GEN_394 = 4'h0 == _T_49 ? result64[63:32] : _GEN_378; // @[cacheLookupUnit.scala 360:{57,57}]
  wire [31:0] _GEN_395 = 4'h1 == _T_49 ? result64[63:32] : _GEN_379; // @[cacheLookupUnit.scala 360:{57,57}]
  wire [31:0] _GEN_396 = 4'h2 == _T_49 ? result64[63:32] : _GEN_380; // @[cacheLookupUnit.scala 360:{57,57}]
  wire [31:0] _GEN_397 = 4'h3 == _T_49 ? result64[63:32] : _GEN_381; // @[cacheLookupUnit.scala 360:{57,57}]
  wire [31:0] _GEN_398 = 4'h4 == _T_49 ? result64[63:32] : _GEN_382; // @[cacheLookupUnit.scala 360:{57,57}]
  wire [31:0] _GEN_399 = 4'h5 == _T_49 ? result64[63:32] : _GEN_383; // @[cacheLookupUnit.scala 360:{57,57}]
  wire [31:0] _GEN_400 = 4'h6 == _T_49 ? result64[63:32] : _GEN_384; // @[cacheLookupUnit.scala 360:{57,57}]
  wire [31:0] _GEN_401 = 4'h7 == _T_49 ? result64[63:32] : _GEN_385; // @[cacheLookupUnit.scala 360:{57,57}]
  wire [31:0] _GEN_402 = 4'h8 == _T_49 ? result64[63:32] : _GEN_386; // @[cacheLookupUnit.scala 360:{57,57}]
  wire [31:0] _GEN_403 = 4'h9 == _T_49 ? result64[63:32] : _GEN_387; // @[cacheLookupUnit.scala 360:{57,57}]
  wire [31:0] _GEN_404 = 4'ha == _T_49 ? result64[63:32] : _GEN_388; // @[cacheLookupUnit.scala 360:{57,57}]
  wire [31:0] _GEN_405 = 4'hb == _T_49 ? result64[63:32] : _GEN_389; // @[cacheLookupUnit.scala 360:{57,57}]
  wire [31:0] _GEN_406 = 4'hc == _T_49 ? result64[63:32] : _GEN_390; // @[cacheLookupUnit.scala 360:{57,57}]
  wire [31:0] _GEN_407 = 4'hd == _T_49 ? result64[63:32] : _GEN_391; // @[cacheLookupUnit.scala 360:{57,57}]
  wire [31:0] _GEN_408 = 4'he == _T_49 ? result64[63:32] : _GEN_392; // @[cacheLookupUnit.scala 360:{57,57}]
  wire [31:0] _GEN_409 = 4'hf == _T_49 ? result64[63:32] : _GEN_393; // @[cacheLookupUnit.scala 360:{57,57}]
  wire [31:0] _GEN_411 = readBuffer_core_instruction[14:12] == 3'h3 ? _GEN_394 : _GEN_353; // @[cacheLookupUnit.scala 347:62]
  wire [31:0] _GEN_412 = readBuffer_core_instruction[14:12] == 3'h3 ? _GEN_395 : _GEN_354; // @[cacheLookupUnit.scala 347:62]
  wire [31:0] _GEN_413 = readBuffer_core_instruction[14:12] == 3'h3 ? _GEN_396 : _GEN_355; // @[cacheLookupUnit.scala 347:62]
  wire [31:0] _GEN_414 = readBuffer_core_instruction[14:12] == 3'h3 ? _GEN_397 : _GEN_356; // @[cacheLookupUnit.scala 347:62]
  wire [31:0] _GEN_415 = readBuffer_core_instruction[14:12] == 3'h3 ? _GEN_398 : _GEN_357; // @[cacheLookupUnit.scala 347:62]
  wire [31:0] _GEN_416 = readBuffer_core_instruction[14:12] == 3'h3 ? _GEN_399 : _GEN_358; // @[cacheLookupUnit.scala 347:62]
  wire [31:0] _GEN_417 = readBuffer_core_instruction[14:12] == 3'h3 ? _GEN_400 : _GEN_359; // @[cacheLookupUnit.scala 347:62]
  wire [31:0] _GEN_418 = readBuffer_core_instruction[14:12] == 3'h3 ? _GEN_401 : _GEN_360; // @[cacheLookupUnit.scala 347:62]
  wire [31:0] _GEN_419 = readBuffer_core_instruction[14:12] == 3'h3 ? _GEN_402 : _GEN_361; // @[cacheLookupUnit.scala 347:62]
  wire [31:0] _GEN_420 = readBuffer_core_instruction[14:12] == 3'h3 ? _GEN_403 : _GEN_362; // @[cacheLookupUnit.scala 347:62]
  wire [31:0] _GEN_421 = readBuffer_core_instruction[14:12] == 3'h3 ? _GEN_404 : _GEN_363; // @[cacheLookupUnit.scala 347:62]
  wire [31:0] _GEN_422 = readBuffer_core_instruction[14:12] == 3'h3 ? _GEN_405 : _GEN_364; // @[cacheLookupUnit.scala 347:62]
  wire [31:0] _GEN_423 = readBuffer_core_instruction[14:12] == 3'h3 ? _GEN_406 : _GEN_365; // @[cacheLookupUnit.scala 347:62]
  wire [31:0] _GEN_424 = readBuffer_core_instruction[14:12] == 3'h3 ? _GEN_407 : _GEN_366; // @[cacheLookupUnit.scala 347:62]
  wire [31:0] _GEN_425 = readBuffer_core_instruction[14:12] == 3'h3 ? _GEN_408 : _GEN_367; // @[cacheLookupUnit.scala 347:62]
  wire [31:0] _GEN_426 = readBuffer_core_instruction[14:12] == 3'h3 ? _GEN_409 : _GEN_368; // @[cacheLookupUnit.scala 347:62]
  wire  _T_51 = 2'h0 == readBuffer_core_instruction[13:12]; // @[cacheLookupUnit.scala 363:53]
  wire [3:0] _T_53 = {{1'd0}, readBuffer_address[2:0]}; // @[cacheLookupUnit.scala 364:88]
  wire [7:0] _GEN_427 = 3'h0 == _T_53[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[7:0]; // @[cacheLookupUnit.scala 270:46 364:{95,95}]
  wire [7:0] _GEN_428 = 3'h1 == _T_53[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[15:8]; // @[cacheLookupUnit.scala 270:46 364:{95,95}]
  wire [7:0] _GEN_429 = 3'h2 == _T_53[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[23:16]; // @[cacheLookupUnit.scala 270:46 364:{95,95}]
  wire [7:0] _GEN_430 = 3'h3 == _T_53[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[31:24]; // @[cacheLookupUnit.scala 270:46 364:{95,95}]
  wire [7:0] _GEN_431 = 3'h4 == _T_53[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[39:32]; // @[cacheLookupUnit.scala 270:46 364:{95,95}]
  wire [7:0] _GEN_432 = 3'h5 == _T_53[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[47:40]; // @[cacheLookupUnit.scala 270:46 364:{95,95}]
  wire [7:0] _GEN_433 = 3'h6 == _T_53[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[55:48]; // @[cacheLookupUnit.scala 270:46 364:{95,95}]
  wire [7:0] _GEN_434 = 3'h7 == _T_53[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[63:56]; // @[cacheLookupUnit.scala 270:46 364:{95,95}]
  wire  _T_55 = 2'h1 == readBuffer_core_instruction[13:12]; // @[cacheLookupUnit.scala 363:53]
  wire [3:0] _T_57 = readBuffer_address[2:1] * 2'h2; // @[cacheLookupUnit.scala 365:87]
  wire [4:0] _T_58 = {{1'd0}, _T_57}; // @[cacheLookupUnit.scala 365:92]
  wire [7:0] _GEN_435 = 3'h0 == _T_58[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[7:0]; // @[cacheLookupUnit.scala 270:46 365:{99,99}]
  wire [7:0] _GEN_436 = 3'h1 == _T_58[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[15:8]; // @[cacheLookupUnit.scala 270:46 365:{99,99}]
  wire [7:0] _GEN_437 = 3'h2 == _T_58[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[23:16]; // @[cacheLookupUnit.scala 270:46 365:{99,99}]
  wire [7:0] _GEN_438 = 3'h3 == _T_58[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[31:24]; // @[cacheLookupUnit.scala 270:46 365:{99,99}]
  wire [7:0] _GEN_439 = 3'h4 == _T_58[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[39:32]; // @[cacheLookupUnit.scala 270:46 365:{99,99}]
  wire [7:0] _GEN_440 = 3'h5 == _T_58[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[47:40]; // @[cacheLookupUnit.scala 270:46 365:{99,99}]
  wire [7:0] _GEN_441 = 3'h6 == _T_58[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[55:48]; // @[cacheLookupUnit.scala 270:46 365:{99,99}]
  wire [7:0] _GEN_442 = 3'h7 == _T_58[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[63:56]; // @[cacheLookupUnit.scala 270:46 365:{99,99}]
  wire [3:0] _T_64 = _T_57 + 4'h1; // @[cacheLookupUnit.scala 365:92]
  wire [7:0] _GEN_443 = 3'h0 == _T_64[2:0] ? readBuffer_writeData_data[15:8] : _GEN_435; // @[cacheLookupUnit.scala 365:{99,99}]
  wire [7:0] _GEN_444 = 3'h1 == _T_64[2:0] ? readBuffer_writeData_data[15:8] : _GEN_436; // @[cacheLookupUnit.scala 365:{99,99}]
  wire [7:0] _GEN_445 = 3'h2 == _T_64[2:0] ? readBuffer_writeData_data[15:8] : _GEN_437; // @[cacheLookupUnit.scala 365:{99,99}]
  wire [7:0] _GEN_446 = 3'h3 == _T_64[2:0] ? readBuffer_writeData_data[15:8] : _GEN_438; // @[cacheLookupUnit.scala 365:{99,99}]
  wire [7:0] _GEN_447 = 3'h4 == _T_64[2:0] ? readBuffer_writeData_data[15:8] : _GEN_439; // @[cacheLookupUnit.scala 365:{99,99}]
  wire [7:0] _GEN_448 = 3'h5 == _T_64[2:0] ? readBuffer_writeData_data[15:8] : _GEN_440; // @[cacheLookupUnit.scala 365:{99,99}]
  wire [7:0] _GEN_449 = 3'h6 == _T_64[2:0] ? readBuffer_writeData_data[15:8] : _GEN_441; // @[cacheLookupUnit.scala 365:{99,99}]
  wire [7:0] _GEN_450 = 3'h7 == _T_64[2:0] ? readBuffer_writeData_data[15:8] : _GEN_442; // @[cacheLookupUnit.scala 365:{99,99}]
  wire  _T_66 = 2'h2 == readBuffer_core_instruction[13:12]; // @[cacheLookupUnit.scala 363:53]
  wire [3:0] _T_68 = readBuffer_address[2] * 3'h4; // @[cacheLookupUnit.scala 366:84]
  wire [4:0] _T_69 = {{1'd0}, _T_68}; // @[cacheLookupUnit.scala 366:89]
  wire [7:0] _GEN_451 = 3'h0 == _T_69[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[7:0]; // @[cacheLookupUnit.scala 270:46 366:{96,96}]
  wire [7:0] _GEN_452 = 3'h1 == _T_69[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[15:8]; // @[cacheLookupUnit.scala 270:46 366:{96,96}]
  wire [7:0] _GEN_453 = 3'h2 == _T_69[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[23:16]; // @[cacheLookupUnit.scala 270:46 366:{96,96}]
  wire [7:0] _GEN_454 = 3'h3 == _T_69[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[31:24]; // @[cacheLookupUnit.scala 270:46 366:{96,96}]
  wire [7:0] _GEN_455 = 3'h4 == _T_69[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[39:32]; // @[cacheLookupUnit.scala 270:46 366:{96,96}]
  wire [7:0] _GEN_456 = 3'h5 == _T_69[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[47:40]; // @[cacheLookupUnit.scala 270:46 366:{96,96}]
  wire [7:0] _GEN_457 = 3'h6 == _T_69[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[55:48]; // @[cacheLookupUnit.scala 270:46 366:{96,96}]
  wire [7:0] _GEN_458 = 3'h7 == _T_69[2:0] ? readBuffer_writeData_data[7:0] : doubleWordWrite[63:56]; // @[cacheLookupUnit.scala 270:46 366:{96,96}]
  wire [3:0] _T_75 = _T_68 + 4'h1; // @[cacheLookupUnit.scala 366:89]
  wire [7:0] _GEN_459 = 3'h0 == _T_75[2:0] ? readBuffer_writeData_data[15:8] : _GEN_451; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_460 = 3'h1 == _T_75[2:0] ? readBuffer_writeData_data[15:8] : _GEN_452; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_461 = 3'h2 == _T_75[2:0] ? readBuffer_writeData_data[15:8] : _GEN_453; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_462 = 3'h3 == _T_75[2:0] ? readBuffer_writeData_data[15:8] : _GEN_454; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_463 = 3'h4 == _T_75[2:0] ? readBuffer_writeData_data[15:8] : _GEN_455; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_464 = 3'h5 == _T_75[2:0] ? readBuffer_writeData_data[15:8] : _GEN_456; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_465 = 3'h6 == _T_75[2:0] ? readBuffer_writeData_data[15:8] : _GEN_457; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_466 = 3'h7 == _T_75[2:0] ? readBuffer_writeData_data[15:8] : _GEN_458; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [3:0] _T_80 = _T_68 + 4'h2; // @[cacheLookupUnit.scala 366:89]
  wire [7:0] _GEN_467 = 3'h0 == _T_80[2:0] ? readBuffer_writeData_data[23:16] : _GEN_459; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_468 = 3'h1 == _T_80[2:0] ? readBuffer_writeData_data[23:16] : _GEN_460; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_469 = 3'h2 == _T_80[2:0] ? readBuffer_writeData_data[23:16] : _GEN_461; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_470 = 3'h3 == _T_80[2:0] ? readBuffer_writeData_data[23:16] : _GEN_462; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_471 = 3'h4 == _T_80[2:0] ? readBuffer_writeData_data[23:16] : _GEN_463; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_472 = 3'h5 == _T_80[2:0] ? readBuffer_writeData_data[23:16] : _GEN_464; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_473 = 3'h6 == _T_80[2:0] ? readBuffer_writeData_data[23:16] : _GEN_465; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_474 = 3'h7 == _T_80[2:0] ? readBuffer_writeData_data[23:16] : _GEN_466; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [3:0] _T_85 = _T_68 + 4'h3; // @[cacheLookupUnit.scala 366:89]
  wire [7:0] _GEN_475 = 3'h0 == _T_85[2:0] ? readBuffer_writeData_data[31:24] : _GEN_467; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_476 = 3'h1 == _T_85[2:0] ? readBuffer_writeData_data[31:24] : _GEN_468; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_477 = 3'h2 == _T_85[2:0] ? readBuffer_writeData_data[31:24] : _GEN_469; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_478 = 3'h3 == _T_85[2:0] ? readBuffer_writeData_data[31:24] : _GEN_470; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_479 = 3'h4 == _T_85[2:0] ? readBuffer_writeData_data[31:24] : _GEN_471; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_480 = 3'h5 == _T_85[2:0] ? readBuffer_writeData_data[31:24] : _GEN_472; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_481 = 3'h6 == _T_85[2:0] ? readBuffer_writeData_data[31:24] : _GEN_473; // @[cacheLookupUnit.scala 366:{96,96}]
  wire [7:0] _GEN_482 = 3'h7 == _T_85[2:0] ? readBuffer_writeData_data[31:24] : _GEN_474; // @[cacheLookupUnit.scala 366:{96,96}]
  wire  _T_87 = 2'h3 == readBuffer_core_instruction[13:12]; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_483 = 2'h3 == readBuffer_core_instruction[13:12] ? readBuffer_writeData_data[7:0] : doubleWordWrite[7:
    0]; // @[cacheLookupUnit.scala 270:46 363:53 367:68]
  wire [7:0] _GEN_484 = 2'h3 == readBuffer_core_instruction[13:12] ? readBuffer_writeData_data[15:8] : doubleWordWrite[
    15:8]; // @[cacheLookupUnit.scala 270:46 363:53 367:68]
  wire [7:0] _GEN_485 = 2'h3 == readBuffer_core_instruction[13:12] ? readBuffer_writeData_data[23:16] : doubleWordWrite[
    23:16]; // @[cacheLookupUnit.scala 270:46 363:53 367:68]
  wire [7:0] _GEN_486 = 2'h3 == readBuffer_core_instruction[13:12] ? readBuffer_writeData_data[31:24] : doubleWordWrite[
    31:24]; // @[cacheLookupUnit.scala 270:46 363:53 367:68]
  wire [7:0] _GEN_487 = 2'h3 == readBuffer_core_instruction[13:12] ? readBuffer_writeData_data[39:32] : doubleWordWrite[
    39:32]; // @[cacheLookupUnit.scala 270:46 363:53 367:68]
  wire [7:0] _GEN_488 = 2'h3 == readBuffer_core_instruction[13:12] ? readBuffer_writeData_data[47:40] : doubleWordWrite[
    47:40]; // @[cacheLookupUnit.scala 270:46 363:53 367:68]
  wire [7:0] _GEN_489 = 2'h3 == readBuffer_core_instruction[13:12] ? readBuffer_writeData_data[55:48] : doubleWordWrite[
    55:48]; // @[cacheLookupUnit.scala 270:46 363:53 367:68]
  wire [7:0] _GEN_490 = 2'h3 == readBuffer_core_instruction[13:12] ? readBuffer_writeData_data[63:56] : doubleWordWrite[
    63:56]; // @[cacheLookupUnit.scala 270:46 363:53 367:68]
  wire [7:0] _GEN_491 = 2'h2 == readBuffer_core_instruction[13:12] ? _GEN_475 : _GEN_483; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_492 = 2'h2 == readBuffer_core_instruction[13:12] ? _GEN_476 : _GEN_484; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_493 = 2'h2 == readBuffer_core_instruction[13:12] ? _GEN_477 : _GEN_485; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_494 = 2'h2 == readBuffer_core_instruction[13:12] ? _GEN_478 : _GEN_486; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_495 = 2'h2 == readBuffer_core_instruction[13:12] ? _GEN_479 : _GEN_487; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_496 = 2'h2 == readBuffer_core_instruction[13:12] ? _GEN_480 : _GEN_488; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_497 = 2'h2 == readBuffer_core_instruction[13:12] ? _GEN_481 : _GEN_489; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_498 = 2'h2 == readBuffer_core_instruction[13:12] ? _GEN_482 : _GEN_490; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_499 = 2'h1 == readBuffer_core_instruction[13:12] ? _GEN_443 : _GEN_491; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_500 = 2'h1 == readBuffer_core_instruction[13:12] ? _GEN_444 : _GEN_492; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_501 = 2'h1 == readBuffer_core_instruction[13:12] ? _GEN_445 : _GEN_493; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_502 = 2'h1 == readBuffer_core_instruction[13:12] ? _GEN_446 : _GEN_494; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_503 = 2'h1 == readBuffer_core_instruction[13:12] ? _GEN_447 : _GEN_495; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_504 = 2'h1 == readBuffer_core_instruction[13:12] ? _GEN_448 : _GEN_496; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_505 = 2'h1 == readBuffer_core_instruction[13:12] ? _GEN_449 : _GEN_497; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_506 = 2'h1 == readBuffer_core_instruction[13:12] ? _GEN_450 : _GEN_498; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_507 = 2'h0 == readBuffer_core_instruction[13:12] ? _GEN_427 : _GEN_499; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_508 = 2'h0 == readBuffer_core_instruction[13:12] ? _GEN_428 : _GEN_500; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_509 = 2'h0 == readBuffer_core_instruction[13:12] ? _GEN_429 : _GEN_501; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_510 = 2'h0 == readBuffer_core_instruction[13:12] ? _GEN_430 : _GEN_502; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_511 = 2'h0 == readBuffer_core_instruction[13:12] ? _GEN_431 : _GEN_503; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_512 = 2'h0 == readBuffer_core_instruction[13:12] ? _GEN_432 : _GEN_504; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_513 = 2'h0 == readBuffer_core_instruction[13:12] ? _GEN_433 : _GEN_505; // @[cacheLookupUnit.scala 363:53]
  wire [7:0] _GEN_514 = 2'h0 == readBuffer_core_instruction[13:12] ? _GEN_434 : _GEN_506; // @[cacheLookupUnit.scala 363:53]
  wire [4:0] _T_89 = readBuffer_address[5:3] * 2'h2; // @[cacheLookupUnit.scala 369:50]
  wire [7:0] _GEN_566 = isAtmoicWriteWire ? doubleWordWrite[15:8] : _GEN_508; // @[cacheLookupUnit.scala 332:30 270:46]
  wire [7:0] writeByteChunks_1 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_566 : doubleWordWrite[15:8]; // @[cacheLookupUnit.scala 270:46 313:61]
  wire [7:0] _GEN_565 = isAtmoicWriteWire ? doubleWordWrite[7:0] : _GEN_507; // @[cacheLookupUnit.scala 332:30 270:46]
  wire [7:0] writeByteChunks_0 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_565 : doubleWordWrite[7:0]; // @[cacheLookupUnit.scala 270:46 313:61]
  wire [7:0] _GEN_568 = isAtmoicWriteWire ? doubleWordWrite[31:24] : _GEN_510; // @[cacheLookupUnit.scala 332:30 270:46]
  wire [7:0] writeByteChunks_3 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_568 : doubleWordWrite[31:24]; // @[cacheLookupUnit.scala 270:46 313:61]
  wire [7:0] _GEN_567 = isAtmoicWriteWire ? doubleWordWrite[23:16] : _GEN_509; // @[cacheLookupUnit.scala 332:30 270:46]
  wire [7:0] writeByteChunks_2 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_567 : doubleWordWrite[23:16]; // @[cacheLookupUnit.scala 270:46 313:61]
  wire [31:0] _newWriteChunks_T_18 = {writeByteChunks_3,writeByteChunks_2,writeByteChunks_1,writeByteChunks_0}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_515 = 4'h0 == _T_89[3:0] ? _newWriteChunks_T_18 : cacheLineChoosen[31:0]; // @[cacheLookupUnit.scala 265:33 369:{56,56}]
  wire [31:0] _GEN_516 = 4'h1 == _T_89[3:0] ? _newWriteChunks_T_18 : cacheLineChoosen[63:32]; // @[cacheLookupUnit.scala 265:33 369:{56,56}]
  wire [31:0] _GEN_517 = 4'h2 == _T_89[3:0] ? _newWriteChunks_T_18 : cacheLineChoosen[95:64]; // @[cacheLookupUnit.scala 265:33 369:{56,56}]
  wire [31:0] _GEN_518 = 4'h3 == _T_89[3:0] ? _newWriteChunks_T_18 : cacheLineChoosen[127:96]; // @[cacheLookupUnit.scala 265:33 369:{56,56}]
  wire [31:0] _GEN_519 = 4'h4 == _T_89[3:0] ? _newWriteChunks_T_18 : cacheLineChoosen[159:128]; // @[cacheLookupUnit.scala 265:33 369:{56,56}]
  wire [31:0] _GEN_520 = 4'h5 == _T_89[3:0] ? _newWriteChunks_T_18 : cacheLineChoosen[191:160]; // @[cacheLookupUnit.scala 265:33 369:{56,56}]
  wire [31:0] _GEN_521 = 4'h6 == _T_89[3:0] ? _newWriteChunks_T_18 : cacheLineChoosen[223:192]; // @[cacheLookupUnit.scala 265:33 369:{56,56}]
  wire [31:0] _GEN_522 = 4'h7 == _T_89[3:0] ? _newWriteChunks_T_18 : cacheLineChoosen[255:224]; // @[cacheLookupUnit.scala 265:33 369:{56,56}]
  wire [31:0] _GEN_523 = 4'h8 == _T_89[3:0] ? _newWriteChunks_T_18 : cacheLineChoosen[287:256]; // @[cacheLookupUnit.scala 265:33 369:{56,56}]
  wire [31:0] _GEN_524 = 4'h9 == _T_89[3:0] ? _newWriteChunks_T_18 : cacheLineChoosen[319:288]; // @[cacheLookupUnit.scala 265:33 369:{56,56}]
  wire [31:0] _GEN_525 = 4'ha == _T_89[3:0] ? _newWriteChunks_T_18 : cacheLineChoosen[351:320]; // @[cacheLookupUnit.scala 265:33 369:{56,56}]
  wire [31:0] _GEN_526 = 4'hb == _T_89[3:0] ? _newWriteChunks_T_18 : cacheLineChoosen[383:352]; // @[cacheLookupUnit.scala 265:33 369:{56,56}]
  wire [31:0] _GEN_527 = 4'hc == _T_89[3:0] ? _newWriteChunks_T_18 : cacheLineChoosen[415:384]; // @[cacheLookupUnit.scala 265:33 369:{56,56}]
  wire [31:0] _GEN_528 = 4'hd == _T_89[3:0] ? _newWriteChunks_T_18 : cacheLineChoosen[447:416]; // @[cacheLookupUnit.scala 265:33 369:{56,56}]
  wire [31:0] _GEN_529 = 4'he == _T_89[3:0] ? _newWriteChunks_T_18 : cacheLineChoosen[479:448]; // @[cacheLookupUnit.scala 265:33 369:{56,56}]
  wire [31:0] _GEN_530 = 4'hf == _T_89[3:0] ? _newWriteChunks_T_18 : cacheLineChoosen[511:480]; // @[cacheLookupUnit.scala 265:33 369:{56,56}]
  wire [4:0] _T_94 = _T_89 + 5'h1; // @[cacheLookupUnit.scala 370:55]
  wire [7:0] _GEN_570 = isAtmoicWriteWire ? doubleWordWrite[47:40] : _GEN_512; // @[cacheLookupUnit.scala 332:30 270:46]
  wire [7:0] writeByteChunks_5 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_570 : doubleWordWrite[47:40]; // @[cacheLookupUnit.scala 270:46 313:61]
  wire [7:0] _GEN_569 = isAtmoicWriteWire ? doubleWordWrite[39:32] : _GEN_511; // @[cacheLookupUnit.scala 332:30 270:46]
  wire [7:0] writeByteChunks_4 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_569 : doubleWordWrite[39:32]; // @[cacheLookupUnit.scala 270:46 313:61]
  wire [7:0] _GEN_572 = isAtmoicWriteWire ? doubleWordWrite[63:56] : _GEN_514; // @[cacheLookupUnit.scala 332:30 270:46]
  wire [7:0] writeByteChunks_7 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_572 : doubleWordWrite[63:56]; // @[cacheLookupUnit.scala 270:46 313:61]
  wire [7:0] _GEN_571 = isAtmoicWriteWire ? doubleWordWrite[55:48] : _GEN_513; // @[cacheLookupUnit.scala 332:30 270:46]
  wire [7:0] writeByteChunks_6 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_571 : doubleWordWrite[55:48]; // @[cacheLookupUnit.scala 270:46 313:61]
  wire [31:0] _newWriteChunks_T_19 = {writeByteChunks_7,writeByteChunks_6,writeByteChunks_5,writeByteChunks_4}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_531 = 4'h0 == _T_94[3:0] ? _newWriteChunks_T_19 : _GEN_515; // @[cacheLookupUnit.scala 370:{62,62}]
  wire [31:0] _GEN_532 = 4'h1 == _T_94[3:0] ? _newWriteChunks_T_19 : _GEN_516; // @[cacheLookupUnit.scala 370:{62,62}]
  wire [31:0] _GEN_533 = 4'h2 == _T_94[3:0] ? _newWriteChunks_T_19 : _GEN_517; // @[cacheLookupUnit.scala 370:{62,62}]
  wire [31:0] _GEN_534 = 4'h3 == _T_94[3:0] ? _newWriteChunks_T_19 : _GEN_518; // @[cacheLookupUnit.scala 370:{62,62}]
  wire [31:0] _GEN_535 = 4'h4 == _T_94[3:0] ? _newWriteChunks_T_19 : _GEN_519; // @[cacheLookupUnit.scala 370:{62,62}]
  wire [31:0] _GEN_536 = 4'h5 == _T_94[3:0] ? _newWriteChunks_T_19 : _GEN_520; // @[cacheLookupUnit.scala 370:{62,62}]
  wire [31:0] _GEN_537 = 4'h6 == _T_94[3:0] ? _newWriteChunks_T_19 : _GEN_521; // @[cacheLookupUnit.scala 370:{62,62}]
  wire [31:0] _GEN_538 = 4'h7 == _T_94[3:0] ? _newWriteChunks_T_19 : _GEN_522; // @[cacheLookupUnit.scala 370:{62,62}]
  wire [31:0] _GEN_539 = 4'h8 == _T_94[3:0] ? _newWriteChunks_T_19 : _GEN_523; // @[cacheLookupUnit.scala 370:{62,62}]
  wire [31:0] _GEN_540 = 4'h9 == _T_94[3:0] ? _newWriteChunks_T_19 : _GEN_524; // @[cacheLookupUnit.scala 370:{62,62}]
  wire [31:0] _GEN_541 = 4'ha == _T_94[3:0] ? _newWriteChunks_T_19 : _GEN_525; // @[cacheLookupUnit.scala 370:{62,62}]
  wire [31:0] _GEN_542 = 4'hb == _T_94[3:0] ? _newWriteChunks_T_19 : _GEN_526; // @[cacheLookupUnit.scala 370:{62,62}]
  wire [31:0] _GEN_543 = 4'hc == _T_94[3:0] ? _newWriteChunks_T_19 : _GEN_527; // @[cacheLookupUnit.scala 370:{62,62}]
  wire [31:0] _GEN_544 = 4'hd == _T_94[3:0] ? _newWriteChunks_T_19 : _GEN_528; // @[cacheLookupUnit.scala 370:{62,62}]
  wire [31:0] _GEN_545 = 4'he == _T_94[3:0] ? _newWriteChunks_T_19 : _GEN_529; // @[cacheLookupUnit.scala 370:{62,62}]
  wire [31:0] _GEN_546 = 4'hf == _T_94[3:0] ? _newWriteChunks_T_19 : _GEN_530; // @[cacheLookupUnit.scala 370:{62,62}]
  wire [31:0] _GEN_548 = isAtmoicWriteWire ? _GEN_411 : _GEN_531; // @[cacheLookupUnit.scala 332:30]
  wire [31:0] _GEN_549 = isAtmoicWriteWire ? _GEN_412 : _GEN_532; // @[cacheLookupUnit.scala 332:30]
  wire [31:0] _GEN_550 = isAtmoicWriteWire ? _GEN_413 : _GEN_533; // @[cacheLookupUnit.scala 332:30]
  wire [31:0] _GEN_551 = isAtmoicWriteWire ? _GEN_414 : _GEN_534; // @[cacheLookupUnit.scala 332:30]
  wire [31:0] _GEN_552 = isAtmoicWriteWire ? _GEN_415 : _GEN_535; // @[cacheLookupUnit.scala 332:30]
  wire [31:0] _GEN_553 = isAtmoicWriteWire ? _GEN_416 : _GEN_536; // @[cacheLookupUnit.scala 332:30]
  wire [31:0] _GEN_554 = isAtmoicWriteWire ? _GEN_417 : _GEN_537; // @[cacheLookupUnit.scala 332:30]
  wire [31:0] _GEN_555 = isAtmoicWriteWire ? _GEN_418 : _GEN_538; // @[cacheLookupUnit.scala 332:30]
  wire [31:0] _GEN_556 = isAtmoicWriteWire ? _GEN_419 : _GEN_539; // @[cacheLookupUnit.scala 332:30]
  wire [31:0] _GEN_557 = isAtmoicWriteWire ? _GEN_420 : _GEN_540; // @[cacheLookupUnit.scala 332:30]
  wire [31:0] _GEN_558 = isAtmoicWriteWire ? _GEN_421 : _GEN_541; // @[cacheLookupUnit.scala 332:30]
  wire [31:0] _GEN_559 = isAtmoicWriteWire ? _GEN_422 : _GEN_542; // @[cacheLookupUnit.scala 332:30]
  wire [31:0] _GEN_560 = isAtmoicWriteWire ? _GEN_423 : _GEN_543; // @[cacheLookupUnit.scala 332:30]
  wire [31:0] _GEN_561 = isAtmoicWriteWire ? _GEN_424 : _GEN_544; // @[cacheLookupUnit.scala 332:30]
  wire [31:0] _GEN_562 = isAtmoicWriteWire ? _GEN_425 : _GEN_545; // @[cacheLookupUnit.scala 332:30]
  wire [31:0] _GEN_563 = isAtmoicWriteWire ? _GEN_426 : _GEN_546; // @[cacheLookupUnit.scala 332:30]
  wire  _GEN_573 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_290 : _GEN_248; // @[cacheLookupUnit.scala 313:61]
  wire  _GEN_574 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_291 : _GEN_245; // @[cacheLookupUnit.scala 313:61]
  wire  _GEN_575 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_292 : _GEN_246; // @[cacheLookupUnit.scala 313:61]
  wire  _GEN_576 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_293 : _GEN_247; // @[cacheLookupUnit.scala 313:61]
  wire [18:0] newAddrWire = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_294 : _GEN_249; // @[cacheLookupUnit.scala 313:61]
  wire [31:0] newWriteChunks_0 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_548 : cacheLineChoosen[31:0]; // @[cacheLookupUnit.scala 265:33 313:61]
  wire [31:0] newWriteChunks_1 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_549 : cacheLineChoosen[63:32]; // @[cacheLookupUnit.scala 265:33 313:61]
  wire [31:0] newWriteChunks_2 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_550 : cacheLineChoosen[95:64]; // @[cacheLookupUnit.scala 265:33 313:61]
  wire [31:0] newWriteChunks_3 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_551 : cacheLineChoosen[127:96]; // @[cacheLookupUnit.scala 265:33 313:61]
  wire [31:0] newWriteChunks_4 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_552 : cacheLineChoosen[159:128]; // @[cacheLookupUnit.scala 265:33 313:61]
  wire [31:0] newWriteChunks_5 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_553 : cacheLineChoosen[191:160]; // @[cacheLookupUnit.scala 265:33 313:61]
  wire [31:0] newWriteChunks_6 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_554 : cacheLineChoosen[223:192]; // @[cacheLookupUnit.scala 265:33 313:61]
  wire [31:0] newWriteChunks_7 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_555 : cacheLineChoosen[255:224]; // @[cacheLookupUnit.scala 265:33 313:61]
  wire [31:0] newWriteChunks_8 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_556 : cacheLineChoosen[287:256]; // @[cacheLookupUnit.scala 265:33 313:61]
  wire [31:0] newWriteChunks_9 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_557 : cacheLineChoosen[319:288]; // @[cacheLookupUnit.scala 265:33 313:61]
  wire [31:0] newWriteChunks_10 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_558 : cacheLineChoosen[351:320]
    ; // @[cacheLookupUnit.scala 265:33 313:61]
  wire [31:0] newWriteChunks_11 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_559 : cacheLineChoosen[383:352]
    ; // @[cacheLookupUnit.scala 265:33 313:61]
  wire [31:0] newWriteChunks_12 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_560 : cacheLineChoosen[415:384]
    ; // @[cacheLookupUnit.scala 265:33 313:61]
  wire [31:0] newWriteChunks_13 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_561 : cacheLineChoosen[447:416]
    ; // @[cacheLookupUnit.scala 265:33 313:61]
  wire [31:0] newWriteChunks_14 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_562 : cacheLineChoosen[479:448]
    ; // @[cacheLookupUnit.scala 265:33 313:61]
  wire [31:0] newWriteChunks_15 = isWriteWire | isAtmoicWriteWire | isSCWriteWire ? _GEN_563 : cacheLineChoosen[511:480]
    ; // @[cacheLookupUnit.scala 265:33 313:61]
  wire  _newShareBitWire_T_9 = readBuffer_cacheLine_response[0] & _isPermissionMiss_T; // @[cacheLookupUnit.scala 380:65]
  wire  _GEN_620 = readBuffer_cacheLine_response[1] ? 1'h0 : _GEN_575; // @[cacheLookupUnit.scala 374:45 375:25]
  wire  _GEN_621 = readBuffer_cacheLine_response[1] ? 1'h0 : _GEN_574; // @[cacheLookupUnit.scala 374:45 376:24]
  wire  _GEN_622 = readBuffer_cacheLine_response[1] ? 1'h0 : readBuffer_cacheLine_response[0] & _isPermissionMiss_T |
    shareBitWire; // @[cacheLookupUnit.scala 374:45 377:25 380:25]
  wire  _GEN_623 = readBuffer_cacheLine_response[1] ? 1'h0 : _GEN_573; // @[cacheLookupUnit.scala 374:45 378:25]
  wire  newValidBitWire = isCoherentWire ? _GEN_620 : _GEN_575; // @[cacheLookupUnit.scala 373:25]
  wire  newPLRUBitWire = isCoherentWire ? _GEN_621 : _GEN_574; // @[cacheLookupUnit.scala 373:25]
  wire  newShareBitWire = isCoherentWire ? _GEN_622 : _GEN_576; // @[cacheLookupUnit.scala 373:25]
  wire  newDirtyBitWire = isCoherentWire ? _GEN_623 : _GEN_573; // @[cacheLookupUnit.scala 373:25]
  wire  isReservationMatch32 = reservationRegister_address[31:2] == readBuffer_address[31:2]; // @[cacheLookupUnit.scala 383:91]
  wire  isReservationMatch64 = reservationRegister_address[31:3] == readBuffer_address[31:3]; // @[cacheLookupUnit.scala 384:91]
  wire  isReservationMatch = reservationRegister_size ? isReservationMatch64 : isReservationMatch32; // @[cacheLookupUnit.scala 385:33]
  wire  _GEN_628 = reservationRegister_size ? ~isReservationMatch64 : reservationRegister_reserved; // @[cacheLookupUnit.scala 121:36 387:39 389:46]
  wire  _GEN_629 = ~reservationRegister_size ? ~isReservationMatch32 : _GEN_628; // @[cacheLookupUnit.scala 387:39 388:46]
  wire  _GEN_630 = reservationRegister_reserved & (isCoherentWire | isWriteWire | isAtmoicWriteWire) ? _GEN_629 :
    reservationRegister_reserved; // @[cacheLookupUnit.scala 121:36 386:96]
  wire [1:0] updatingSet = isDataMissWire ? replacingset : hitTagWire; // @[cacheLookupUnit.scala 394:26]
  wire [22:0] _newtagChunks_0_T_2 = tagChunks_0 & 23'h3fffff; // @[cacheLookupUnit.scala 397:41]
  wire [22:0] _newtagChunks_1_T_2 = tagChunks_1 & 23'h3fffff; // @[cacheLookupUnit.scala 397:41]
  wire [22:0] _newtagChunks_2_T_2 = tagChunks_2 & 23'h3fffff; // @[cacheLookupUnit.scala 397:41]
  wire [22:0] _newtagChunks_3_T_2 = tagChunks_3 & 23'h3fffff; // @[cacheLookupUnit.scala 397:41]
  wire [22:0] _GEN_631 = _newPLRUBitWire_T_5 ? _newtagChunks_0_T_2 : tagChunks_0; // @[cacheLookupUnit.scala 395:36 397:25 251:31]
  wire [22:0] _GEN_632 = _newPLRUBitWire_T_5 ? _newtagChunks_1_T_2 : tagChunks_1; // @[cacheLookupUnit.scala 395:36 397:25 251:31]
  wire [22:0] _GEN_633 = _newPLRUBitWire_T_5 ? _newtagChunks_2_T_2 : tagChunks_2; // @[cacheLookupUnit.scala 395:36 397:25 251:31]
  wire [22:0] _GEN_634 = _newPLRUBitWire_T_5 ? _newtagChunks_3_T_2 : tagChunks_3; // @[cacheLookupUnit.scala 395:36 397:25 251:31]
  wire [22:0] _newtagChunks_T_4 = {newPLRUBitWire,newShareBitWire,newDirtyBitWire,newValidBitWire,newAddrWire}; // @[Cat.scala 33:92]
  wire [22:0] newtagChunks_0 = 2'h0 == updatingSet ? _newtagChunks_T_4 : _GEN_631; // @[cacheLookupUnit.scala 400:{31,31}]
  wire [22:0] newtagChunks_1 = 2'h1 == updatingSet ? _newtagChunks_T_4 : _GEN_632; // @[cacheLookupUnit.scala 400:{31,31}]
  wire [22:0] newtagChunks_2 = 2'h2 == updatingSet ? _newtagChunks_T_4 : _GEN_633; // @[cacheLookupUnit.scala 400:{31,31}]
  wire [22:0] newtagChunks_3 = 2'h3 == updatingSet ? _newtagChunks_T_4 : _GEN_634; // @[cacheLookupUnit.scala 400:{31,31}]
  wire [91:0] _tagBRAM_wrData_T_2 = {newtagChunks_3,newtagChunks_2,newtagChunks_1,newtagChunks_0}; // @[Cat.scala 33:92]
  wire  _T_126 = reservationRegister_reserved & isReservationMatch; // @[cacheLookupUnit.scala 457:41]
  wire  _T_125 = isReplayValidWire | _T_18; // @[cacheLookupUnit.scala 443:30]
  wire  _T_115 = _cacheLineChoosen_T | _isPermissionMiss_T; // @[cacheLookupUnit.scala 414:48]
  wire  _GEN_653 = (_cacheLineChoosen_T | _isPermissionMiss_T) & _cacheLineChoosen_T; // @[cacheLookupUnit.scala 414:67 418:28]
  wire  _GEN_658 = isReadWire & _GEN_653; // @[cacheLookupUnit.scala 413:21]
  wire  _GEN_664 = _T_125 ? isReplayValidWire : _GEN_658; // @[cacheLookupUnit.scala 425:72 430:28]
  wire  _GEN_671 = _T_10 ? _GEN_664 : _GEN_658; // @[cacheLookupUnit.scala 424:43]
  wire  _GEN_680 = isReplayValidWire | _T_18 | _GEN_671; // @[cacheLookupUnit.scala 443:72 446:28]
  wire  _GEN_687 = _T_14 ? _GEN_680 : _GEN_671; // @[cacheLookupUnit.scala 442:43]
  wire  _GEN_695 = reservationRegister_reserved & isReservationMatch | _GEN_687; // @[cacheLookupUnit.scala 457:63 460:28]
  wire  dataBRAMUpdateWire = isSCWriteWire ? _GEN_695 : _GEN_687; // @[cacheLookupUnit.scala 455:24]
  wire  _GEN_639 = 2'h0 == updatingSet & dataBRAMUpdateWire; // @[cacheLookupUnit.scala 408:{36,36} 75:28]
  wire  _GEN_640 = 2'h1 == updatingSet & dataBRAMUpdateWire; // @[cacheLookupUnit.scala 408:{36,36} 75:28]
  wire  _GEN_641 = 2'h2 == updatingSet & dataBRAMUpdateWire; // @[cacheLookupUnit.scala 408:{36,36} 75:28]
  wire  _GEN_642 = 2'h3 == updatingSet & dataBRAMUpdateWire; // @[cacheLookupUnit.scala 408:{36,36} 75:28]
  wire [319:0] _dataBRAMVec_wrData_T_8 = {newWriteChunks_15,newWriteChunks_14,newWriteChunks_13,newWriteChunks_12,
    newWriteChunks_11,newWriteChunks_10,newWriteChunks_9,newWriteChunks_8,newWriteChunks_7,newWriteChunks_6}; // @[Cat.scala 33:92]
  wire [511:0] _dataBRAMVec_wrData_T_14 = {_dataBRAMVec_wrData_T_8,newWriteChunks_5,newWriteChunks_4,newWriteChunks_3,
    newWriteChunks_2,newWriteChunks_1,newWriteChunks_0}; // @[Cat.scala 33:92]
  wire [511:0] _GEN_643 = 2'h0 == updatingSet ? _dataBRAMVec_wrData_T_14 : 512'h0; // @[cacheLookupUnit.scala 409:{37,37} 75:28]
  wire [511:0] _GEN_644 = 2'h1 == updatingSet ? _dataBRAMVec_wrData_T_14 : 512'h0; // @[cacheLookupUnit.scala 409:{37,37} 75:28]
  wire [511:0] _GEN_645 = 2'h2 == updatingSet ? _dataBRAMVec_wrData_T_14 : 512'h0; // @[cacheLookupUnit.scala 409:{37,37} 75:28]
  wire [511:0] _GEN_646 = 2'h3 == updatingSet ? _dataBRAMVec_wrData_T_14 : 512'h0; // @[cacheLookupUnit.scala 409:{37,37} 75:28]
  wire [6:0] _GEN_647 = 2'h0 == updatingSet ? readBuffer_address[12:6] : 7'h0; // @[cacheLookupUnit.scala 410:{37,37} 75:28]
  wire [6:0] _GEN_648 = 2'h1 == updatingSet ? readBuffer_address[12:6] : 7'h0; // @[cacheLookupUnit.scala 410:{37,37} 75:28]
  wire [6:0] _GEN_649 = 2'h2 == updatingSet ? readBuffer_address[12:6] : 7'h0; // @[cacheLookupUnit.scala 410:{37,37} 75:28]
  wire [6:0] _GEN_650 = 2'h3 == updatingSet ? readBuffer_address[12:6] : 7'h0; // @[cacheLookupUnit.scala 410:{37,37} 75:28]
  wire  _toWriteBackValidWire_T_1 = isUpdateDirtyWire & isUpdateValidWire & isReplayValidWire; // @[cacheLookupUnit.scala 417:74]
  wire  _GEN_652 = (_cacheLineChoosen_T | _isPermissionMiss_T) & (isUpdateDirtyWire & isUpdateValidWire &
    isReplayValidWire & isDataMissWire); // @[cacheLookupUnit.scala 414:67 417:30]
  wire  _GEN_654 = _cacheLineChoosen_T | _isPermissionMiss_T ? 1'h0 : 1'h1; // @[cacheLookupUnit.scala 414:67 420:27]
  wire  _GEN_656 = isReadWire & _T_115; // @[cacheLookupUnit.scala 413:21]
  wire  _GEN_657 = isReadWire & _GEN_652; // @[cacheLookupUnit.scala 413:21]
  wire  _GEN_659 = isReadWire & _GEN_654; // @[cacheLookupUnit.scala 413:21]
  wire  _GEN_661 = _T_125 | _GEN_656; // @[cacheLookupUnit.scala 425:72 426:35]
  wire  _GEN_663 = _T_125 ? _toWriteBackValidWire_T_1 : _GEN_657; // @[cacheLookupUnit.scala 425:72 429:30]
  wire  _GEN_665 = _T_125 ? _GEN_659 : 1'h1; // @[cacheLookupUnit.scala 425:72 432:27]
  wire [1:0] _GEN_666 = _T_125 ? 2'h0 : 2'h1; // @[cacheLookupUnit.scala 425:72 433:30]
  wire  _GEN_667 = _T_125 ? 1'h0 : 1'h1; // @[cacheLookupUnit.scala 425:72 434:34]
  wire  _GEN_668 = _T_10 ? _GEN_661 : _GEN_656; // @[cacheLookupUnit.scala 424:43]
  wire  _GEN_669 = _T_10 & _T_125; // @[cacheLookupUnit.scala 424:43]
  wire  _GEN_670 = _T_10 ? _GEN_663 : _GEN_657; // @[cacheLookupUnit.scala 424:43]
  wire  _GEN_672 = _T_10 ? _GEN_665 : _GEN_659; // @[cacheLookupUnit.scala 424:43]
  wire [1:0] _GEN_673 = _T_10 ? _GEN_666 : 2'h0; // @[cacheLookupUnit.scala 424:43]
  wire  _GEN_674 = _T_10 & _GEN_667; // @[cacheLookupUnit.scala 424:43]
  wire  _GEN_675 = isLRWriteWire | _GEN_45; // @[cacheLookupUnit.scala 437:{24,54}]
  wire  _GEN_677 = isCoherentWire ? _isPermissionMiss_T : _GEN_668; // @[cacheLookupUnit.scala 438:25 440:24]
  wire [1:0] _requiredResponseWire_T_2 = isPermissionMiss & _isPermissionMiss_T ? 2'h3 : 2'h1; // @[cacheLookupUnit.scala 450:36]
  wire  _GEN_678 = isReplayValidWire | _T_18 ? _toWriteBackValidWire_T_1 : _GEN_670; // @[cacheLookupUnit.scala 443:72 444:30]
  wire  _GEN_679 = isReplayValidWire | _T_18 | _GEN_677; // @[cacheLookupUnit.scala 443:72 445:26]
  wire  _GEN_681 = isReplayValidWire | _T_18 | _GEN_675; // @[cacheLookupUnit.scala 443:72 447:38]
  wire  _GEN_682 = isReplayValidWire | _T_18 ? _GEN_672 : 1'h1; // @[cacheLookupUnit.scala 443:72 449:27]
  wire [1:0] _GEN_683 = isReplayValidWire | _T_18 ? _GEN_673 : _requiredResponseWire_T_2; // @[cacheLookupUnit.scala 443:72 450:30]
  wire  _GEN_684 = isReplayValidWire | _T_18 ? _GEN_674 : 1'h1; // @[cacheLookupUnit.scala 443:72 451:34]
  wire  _GEN_685 = _T_14 ? _GEN_678 : _GEN_670; // @[cacheLookupUnit.scala 442:43]
  wire  _GEN_686 = _T_14 ? _GEN_679 : _GEN_677; // @[cacheLookupUnit.scala 442:43]
  wire  _GEN_688 = _T_14 ? _GEN_681 : _GEN_675; // @[cacheLookupUnit.scala 442:43]
  wire  _GEN_689 = _T_14 ? _GEN_682 : _GEN_672; // @[cacheLookupUnit.scala 442:43]
  wire  _GEN_691 = _T_14 ? _GEN_684 : _GEN_674; // @[cacheLookupUnit.scala 442:43]
  wire  _GEN_692 = isSCReadWire | _GEN_668; // @[cacheLookupUnit.scala 454:{23,50}]
  wire  _GEN_693 = reservationRegister_reserved & isReservationMatch ? isDirtyWire & isReplayValidWire & isDataMissWire
     : _GEN_685; // @[cacheLookupUnit.scala 457:63 458:30]
  wire  _GEN_694 = reservationRegister_reserved & isReservationMatch | _GEN_686; // @[cacheLookupUnit.scala 457:63 459:26]
  wire  _GEN_697 = isSCWriteWire ? _GEN_693 : _GEN_685; // @[cacheLookupUnit.scala 455:24]
  wire  tagBRAMUpdateWire = isSCWriteWire ? _GEN_694 : _GEN_686; // @[cacheLookupUnit.scala 455:24]
  wire  _GEN_700 = isSCWriteWire | _GEN_688; // @[cacheLookupUnit.scala 455:24 462:36]
  wire [63:0] doubleWordChunks_0 = cacheLineChoosen[63:0]; // @[cacheLookupUnit.scala 470:23]
  wire [63:0] doubleWordChunks_1 = cacheLineChoosen[127:64]; // @[cacheLookupUnit.scala 470:23]
  wire [63:0] doubleWordChunks_2 = cacheLineChoosen[191:128]; // @[cacheLookupUnit.scala 470:23]
  wire [63:0] doubleWordChunks_3 = cacheLineChoosen[255:192]; // @[cacheLookupUnit.scala 470:23]
  wire [63:0] doubleWordChunks_4 = cacheLineChoosen[319:256]; // @[cacheLookupUnit.scala 470:23]
  wire [63:0] doubleWordChunks_5 = cacheLineChoosen[383:320]; // @[cacheLookupUnit.scala 470:23]
  wire [63:0] doubleWordChunks_6 = cacheLineChoosen[447:384]; // @[cacheLookupUnit.scala 470:23]
  wire [63:0] doubleWordChunks_7 = cacheLineChoosen[511:448]; // @[cacheLookupUnit.scala 470:23]
  wire [63:0] _GEN_702 = 3'h1 == readBuffer_address[5:3] ? doubleWordChunks_1 : doubleWordChunks_0; // @[cacheLookupUnit.scala 476:{24,24}]
  wire [63:0] _GEN_703 = 3'h2 == readBuffer_address[5:3] ? doubleWordChunks_2 : _GEN_702; // @[cacheLookupUnit.scala 476:{24,24}]
  wire [63:0] _GEN_704 = 3'h3 == readBuffer_address[5:3] ? doubleWordChunks_3 : _GEN_703; // @[cacheLookupUnit.scala 476:{24,24}]
  wire [63:0] _GEN_705 = 3'h4 == readBuffer_address[5:3] ? doubleWordChunks_4 : _GEN_704; // @[cacheLookupUnit.scala 476:{24,24}]
  wire [63:0] _GEN_706 = 3'h5 == readBuffer_address[5:3] ? doubleWordChunks_5 : _GEN_705; // @[cacheLookupUnit.scala 476:{24,24}]
  wire [63:0] _GEN_707 = 3'h6 == readBuffer_address[5:3] ? doubleWordChunks_6 : _GEN_706; // @[cacheLookupUnit.scala 476:{24,24}]
  wire [63:0] _GEN_708 = 3'h7 == readBuffer_address[5:3] ? doubleWordChunks_7 : _GEN_707; // @[cacheLookupUnit.scala 476:{24,24}]
  wire [7:0] byteChunks_0 = _GEN_708[7:0]; // @[cacheLookupUnit.scala 476:24]
  wire [7:0] byteChunks_1 = _GEN_708[15:8]; // @[cacheLookupUnit.scala 476:24]
  wire [7:0] byteChunks_2 = _GEN_708[23:16]; // @[cacheLookupUnit.scala 476:24]
  wire [7:0] byteChunks_3 = _GEN_708[31:24]; // @[cacheLookupUnit.scala 476:24]
  wire [7:0] byteChunks_4 = _GEN_708[39:32]; // @[cacheLookupUnit.scala 476:24]
  wire [7:0] byteChunks_5 = _GEN_708[47:40]; // @[cacheLookupUnit.scala 476:24]
  wire [7:0] byteChunks_6 = _GEN_708[55:48]; // @[cacheLookupUnit.scala 476:24]
  wire [7:0] byteChunks_7 = _GEN_708[63:56]; // @[cacheLookupUnit.scala 476:24]
  wire [3:0] _halfwordChoosed_T_1 = 2'h2 * readBuffer_address[2:1]; // @[cacheLookupUnit.scala 479:46]
  wire [3:0] _halfwordChoosed_T_3 = _halfwordChoosed_T_1 + 4'h1; // @[cacheLookupUnit.scala 479:72]
  wire [7:0] _GEN_710 = 3'h1 == _halfwordChoosed_T_3[2:0] ? byteChunks_1 : byteChunks_0; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_711 = 3'h2 == _halfwordChoosed_T_3[2:0] ? byteChunks_2 : _GEN_710; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_712 = 3'h3 == _halfwordChoosed_T_3[2:0] ? byteChunks_3 : _GEN_711; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_713 = 3'h4 == _halfwordChoosed_T_3[2:0] ? byteChunks_4 : _GEN_712; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_714 = 3'h5 == _halfwordChoosed_T_3[2:0] ? byteChunks_5 : _GEN_713; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_715 = 3'h6 == _halfwordChoosed_T_3[2:0] ? byteChunks_6 : _GEN_714; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_716 = 3'h7 == _halfwordChoosed_T_3[2:0] ? byteChunks_7 : _GEN_715; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_718 = 3'h1 == _halfwordChoosed_T_1[2:0] ? byteChunks_1 : byteChunks_0; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_719 = 3'h2 == _halfwordChoosed_T_1[2:0] ? byteChunks_2 : _GEN_718; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_720 = 3'h3 == _halfwordChoosed_T_1[2:0] ? byteChunks_3 : _GEN_719; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_721 = 3'h4 == _halfwordChoosed_T_1[2:0] ? byteChunks_4 : _GEN_720; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_722 = 3'h5 == _halfwordChoosed_T_1[2:0] ? byteChunks_5 : _GEN_721; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_723 = 3'h6 == _halfwordChoosed_T_1[2:0] ? byteChunks_6 : _GEN_722; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_724 = 3'h7 == _halfwordChoosed_T_1[2:0] ? byteChunks_7 : _GEN_723; // @[Cat.scala 33:{92,92}]
  wire [15:0] halfwordChoosed = {_GEN_716,_GEN_724}; // @[Cat.scala 33:92]
  wire [3:0] _wordChoosed_T_1 = 3'h4 * readBuffer_address[2]; // @[cacheLookupUnit.scala 480:46]
  wire [3:0] _wordChoosed_T_3 = _wordChoosed_T_1 + 4'h3; // @[cacheLookupUnit.scala 480:70]
  wire [3:0] _wordChoosed_T_8 = _wordChoosed_T_1 + 4'h2; // @[cacheLookupUnit.scala 480:116]
  wire [3:0] _wordChoosed_T_13 = _wordChoosed_T_1 + 4'h1; // @[cacheLookupUnit.scala 481:70]
  wire [7:0] _GEN_726 = 3'h1 == _wordChoosed_T_13[2:0] ? byteChunks_1 : byteChunks_0; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_727 = 3'h2 == _wordChoosed_T_13[2:0] ? byteChunks_2 : _GEN_726; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_728 = 3'h3 == _wordChoosed_T_13[2:0] ? byteChunks_3 : _GEN_727; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_729 = 3'h4 == _wordChoosed_T_13[2:0] ? byteChunks_4 : _GEN_728; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_730 = 3'h5 == _wordChoosed_T_13[2:0] ? byteChunks_5 : _GEN_729; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_731 = 3'h6 == _wordChoosed_T_13[2:0] ? byteChunks_6 : _GEN_730; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_732 = 3'h7 == _wordChoosed_T_13[2:0] ? byteChunks_7 : _GEN_731; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_734 = 3'h1 == _wordChoosed_T_1[2:0] ? byteChunks_1 : byteChunks_0; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_735 = 3'h2 == _wordChoosed_T_1[2:0] ? byteChunks_2 : _GEN_734; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_736 = 3'h3 == _wordChoosed_T_1[2:0] ? byteChunks_3 : _GEN_735; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_737 = 3'h4 == _wordChoosed_T_1[2:0] ? byteChunks_4 : _GEN_736; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_738 = 3'h5 == _wordChoosed_T_1[2:0] ? byteChunks_5 : _GEN_737; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_739 = 3'h6 == _wordChoosed_T_1[2:0] ? byteChunks_6 : _GEN_738; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_740 = 3'h7 == _wordChoosed_T_1[2:0] ? byteChunks_7 : _GEN_739; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_742 = 3'h1 == _wordChoosed_T_3[2:0] ? byteChunks_1 : byteChunks_0; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_743 = 3'h2 == _wordChoosed_T_3[2:0] ? byteChunks_2 : _GEN_742; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_744 = 3'h3 == _wordChoosed_T_3[2:0] ? byteChunks_3 : _GEN_743; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_745 = 3'h4 == _wordChoosed_T_3[2:0] ? byteChunks_4 : _GEN_744; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_746 = 3'h5 == _wordChoosed_T_3[2:0] ? byteChunks_5 : _GEN_745; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_747 = 3'h6 == _wordChoosed_T_3[2:0] ? byteChunks_6 : _GEN_746; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_748 = 3'h7 == _wordChoosed_T_3[2:0] ? byteChunks_7 : _GEN_747; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_750 = 3'h1 == _wordChoosed_T_8[2:0] ? byteChunks_1 : byteChunks_0; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_751 = 3'h2 == _wordChoosed_T_8[2:0] ? byteChunks_2 : _GEN_750; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_752 = 3'h3 == _wordChoosed_T_8[2:0] ? byteChunks_3 : _GEN_751; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_753 = 3'h4 == _wordChoosed_T_8[2:0] ? byteChunks_4 : _GEN_752; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_754 = 3'h5 == _wordChoosed_T_8[2:0] ? byteChunks_5 : _GEN_753; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_755 = 3'h6 == _wordChoosed_T_8[2:0] ? byteChunks_6 : _GEN_754; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_756 = 3'h7 == _wordChoosed_T_8[2:0] ? byteChunks_7 : _GEN_755; // @[Cat.scala 33:{92,92}]
  wire [31:0] wordChoosed = {_GEN_748,_GEN_756,_GEN_732,_GEN_740}; // @[Cat.scala 33:92]
  wire [7:0] _GEN_758 = 3'h1 == readBuffer_address[2:0] ? byteChunks_1 : byteChunks_0; // @[cacheLookupUnit.scala 485:{73,73}]
  wire [7:0] _GEN_759 = 3'h2 == readBuffer_address[2:0] ? byteChunks_2 : _GEN_758; // @[cacheLookupUnit.scala 485:{73,73}]
  wire [7:0] _GEN_760 = 3'h3 == readBuffer_address[2:0] ? byteChunks_3 : _GEN_759; // @[cacheLookupUnit.scala 485:{73,73}]
  wire [7:0] _GEN_761 = 3'h4 == readBuffer_address[2:0] ? byteChunks_4 : _GEN_760; // @[cacheLookupUnit.scala 485:{73,73}]
  wire [7:0] _GEN_762 = 3'h5 == readBuffer_address[2:0] ? byteChunks_5 : _GEN_761; // @[cacheLookupUnit.scala 485:{73,73}]
  wire [7:0] _GEN_763 = 3'h6 == readBuffer_address[2:0] ? byteChunks_6 : _GEN_762; // @[cacheLookupUnit.scala 485:{73,73}]
  wire [7:0] _GEN_764 = 3'h7 == readBuffer_address[2:0] ? byteChunks_7 : _GEN_763; // @[cacheLookupUnit.scala 485:{73,73}]
  wire [55:0] _responseResultWire_T_3 = _GEN_764[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _responseResultWire_T_4 = {_responseResultWire_T_3,_GEN_764}; // @[Cat.scala 33:92]
  wire [63:0] _responseResultWire_T_5 = readBuffer_core_instruction[14] ? {{56'd0}, _GEN_764} : _responseResultWire_T_4; // @[cacheLookupUnit.scala 484:44]
  wire [47:0] _responseResultWire_T_9 = halfwordChoosed[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _responseResultWire_T_10 = {_responseResultWire_T_9,_GEN_716,_GEN_724}; // @[Cat.scala 33:92]
  wire [63:0] _responseResultWire_T_11 = readBuffer_core_instruction[14] ? {{48'd0}, halfwordChoosed} :
    _responseResultWire_T_10; // @[cacheLookupUnit.scala 486:44]
  wire [31:0] _responseResultWire_T_15 = wordChoosed[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _responseResultWire_T_16 = {_responseResultWire_T_15,_GEN_748,_GEN_756,_GEN_732,_GEN_740}; // @[Cat.scala 33:92]
  wire [63:0] _responseResultWire_T_17 = readBuffer_core_instruction[14] ? {{32'd0}, wordChoosed} :
    _responseResultWire_T_16; // @[cacheLookupUnit.scala 488:44]
  wire [63:0] _responseResultWire_T_19 = readBuffer_core_instruction[14] ? 64'h0 : _GEN_708; // @[cacheLookupUnit.scala 490:44]
  wire [63:0] _GEN_765 = _T_87 ? _responseResultWire_T_19 : 64'h0; // @[cacheLookupUnit.scala 483:48 490:38]
  wire [63:0] _GEN_766 = _T_66 ? _responseResultWire_T_17 : _GEN_765; // @[cacheLookupUnit.scala 483:48 488:38]
  wire [63:0] _GEN_767 = _T_55 ? _responseResultWire_T_11 : _GEN_766; // @[cacheLookupUnit.scala 483:48 486:38]
  wire [63:0] _GEN_768 = _T_51 ? _responseResultWire_T_5 : _GEN_767; // @[cacheLookupUnit.scala 483:48 484:38]
  wire  _responseResultWire_T_21 = _T_126 ? 1'h0 : 1'h1; // @[cacheLookupUnit.scala 494:32]
  wire  toReplayValidWire = operationValid & _GEN_689; // @[cacheLookupUnit.scala 212:23]
  wire  _GEN_775 = toReplayValidWire & readBuffer_branch_valid ? readBuffer_branch_valid : replayBuffer_branch_valid; // @[cacheLookupUnit.scala 499:55 500:20 153:29]
  wire [4:0] _GEN_776 = toReplayValidWire & readBuffer_branch_valid ? readBuffer_branch_mask : replayBuffer_branch_mask; // @[cacheLookupUnit.scala 499:55 500:20 153:29]
  wire  toMemoryResponseValidWire = operationValid & _GEN_692; // @[cacheLookupUnit.scala 212:23]
  wire  _GEN_787 = toMemoryResponseValidWire & readBuffer_branch_valid ? readBuffer_branch_valid :
    memoryResponseBuffer_branch_valid; // @[cacheLookupUnit.scala 506:63 507:28 160:37]
  wire [4:0] _GEN_788 = toMemoryResponseValidWire & readBuffer_branch_valid ? readBuffer_branch_mask :
    memoryResponseBuffer_branch_mask; // @[cacheLookupUnit.scala 506:63 507:28 160:37]
  wire [511:0] _coherencyResponseBuffer_cacheLine_T_3 = _isPermissionMiss_T ? _GEN_103 : 512'h0; // @[cacheLookupUnit.scala 515:49]
  wire  _coherencyResponseBuffer_response_T_2 = readBuffer_cacheLine_response[1] ? ~isDirtyWire : 1'h1; // @[cacheLookupUnit.scala 517:67]
  wire [1:0] _coherencyResponseBuffer_response_T_3 = {newShareBitWire,_coherencyResponseBuffer_response_T_2}; // @[cacheLookupUnit.scala 517:61]
  wire  toCoherencyResponseValidWire = operationValid & isCoherentWire; // @[cacheLookupUnit.scala 212:23]
  wire [22:0] _GEN_806 = 2'h1 == updatingSet ? tagChunks_1 : tagChunks_0; // @[Cat.scala 33:{92,92}]
  wire [22:0] _GEN_807 = 2'h2 == updatingSet ? tagChunks_2 : _GEN_806; // @[Cat.scala 33:{92,92}]
  wire [22:0] _GEN_808 = 2'h3 == updatingSet ? tagChunks_3 : _GEN_807; // @[Cat.scala 33:{92,92}]
  wire [35:0] _writeBackBuffer_address_T_3 = {_GEN_808,readBuffer_address[12:6],6'h0}; // @[Cat.scala 33:92]
  wire [511:0] _GEN_810 = 2'h1 == updatingSet ? dataBRAMVec_1_rdData : dataBRAMVec_0_rdData; // @[cacheLookupUnit.scala 528:{28,28}]
  wire [511:0] _GEN_811 = 2'h2 == updatingSet ? dataBRAMVec_2_rdData : _GEN_810; // @[cacheLookupUnit.scala 528:{28,28}]
  wire  toWriteBackValidWire = operationValid & _GEN_697; // @[cacheLookupUnit.scala 212:23]
  wire [35:0] _GEN_814 = toWriteBackValidWire ? _writeBackBuffer_address_T_3 : {{4'd0}, writeBackBuffer_address}; // @[cacheLookupUnit.scala 525:31 527:31 177:32]
  wire  toLastMissRecordRegister = operationValid & _GEN_691; // @[cacheLookupUnit.scala 212:23]
  wire  _GEN_821 = toLastMissRecordRegister & readBuffer_branch_valid ? readBuffer_branch_valid :
    lastMissRecordRegister_branch_valid; // @[cacheLookupUnit.scala 532:62 533:30 130:39]
  wire [4:0] _GEN_822 = toLastMissRecordRegister & readBuffer_branch_valid ? readBuffer_branch_mask :
    lastMissRecordRegister_branch_mask; // @[cacheLookupUnit.scala 532:62 533:30 130:39]
  wire  toReservationRegisterWire = operationValid & _GEN_669; // @[cacheLookupUnit.scala 212:23]
  wire  _GEN_859 = operationValid ? _GEN_775 : replayBuffer_branch_valid; // @[cacheLookupUnit.scala 212:23 153:29]
  wire [4:0] _GEN_860 = operationValid ? _GEN_776 : replayBuffer_branch_mask; // @[cacheLookupUnit.scala 212:23 153:29]
  wire  _GEN_871 = operationValid ? _GEN_787 : memoryResponseBuffer_branch_valid; // @[cacheLookupUnit.scala 212:23 160:37]
  wire [4:0] _GEN_872 = operationValid ? _GEN_788 : memoryResponseBuffer_branch_mask; // @[cacheLookupUnit.scala 212:23 160:37]
  wire [35:0] _GEN_883 = operationValid ? _GEN_814 : {{4'd0}, writeBackBuffer_address}; // @[cacheLookupUnit.scala 212:23 177:32]
  wire  _GEN_890 = operationValid ? _GEN_821 : lastMissRecordRegister_branch_valid; // @[cacheLookupUnit.scala 212:23 130:39]
  wire [4:0] _GEN_891 = operationValid ? _GEN_822 : lastMissRecordRegister_branch_mask; // @[cacheLookupUnit.scala 212:23 130:39]
  wire [4:0] _T_136 = readBuffer_branch_mask & branchOps_branchMask; // @[utils.scala 92:27]
  wire  _T_137 = |_T_136; // @[utils.scala 92:51]
  wire [4:0] _replayBuffer_branch_mask_T = readBuffer_branch_mask ^ branchOps_branchMask; // @[utils.scala 93:42]
  wire [4:0] _GEN_899 = |_T_136 ? _replayBuffer_branch_mask_T : readBuffer_branch_mask; // @[utils.scala 92:56 93:27 96:27]
  wire [4:0] _GEN_900 = _T_137 ? 5'h0 : readBuffer_branch_mask; // @[utils.scala 101:56 102:27 106:27]
  wire  _GEN_901 = _T_137 ? 1'h0 : readBuffer_branch_valid; // @[utils.scala 101:56 103:28 107:28]
  wire [4:0] _GEN_902 = branchOps_passed ? _GEN_899 : _GEN_900; // @[utils.scala 90:30]
  wire  _GEN_903 = branchOps_passed ? readBuffer_branch_valid : _GEN_901; // @[utils.scala 90:30 98:26]
  wire [4:0] _T_146 = replayBuffer_branch_mask & branchOps_branchMask; // @[utils.scala 122:29]
  wire  _T_147 = |_T_146; // @[utils.scala 122:53]
  wire [4:0] _replayBuffer_branch_mask_T_1 = replayBuffer_branch_mask ^ branchOps_branchMask; // @[utils.scala 123:40]
  wire [4:0] _GEN_917 = |_T_146 ? _replayBuffer_branch_mask_T_1 : _GEN_860; // @[utils.scala 122:58 123:25]
  wire  _GEN_918 = _T_147 ? 1'h0 : _GEN_859; // @[utils.scala 127:58 128:26]
  wire [4:0] _GEN_919 = _T_147 ? 5'h0 : _GEN_860; // @[utils.scala 127:58 129:25]
  wire [4:0] _GEN_920 = branchOps_passed ? _GEN_917 : _GEN_919; // @[utils.scala 121:32]
  wire  _GEN_921 = branchOps_passed ? replayBuffer_branch_valid : _GEN_918; // @[utils.scala 121:32 125:24]
  wire [4:0] _GEN_922 = branchOps_valid ? _GEN_920 : _GEN_860; // @[utils.scala 120:29]
  wire  _GEN_923 = branchOps_valid ? _GEN_921 : _GEN_859; // @[utils.scala 120:29]
  wire [4:0] _GEN_928 = _T_137 ? _replayBuffer_branch_mask_T : _GEN_57; // @[utils.scala 122:58 123:25]
  wire  _GEN_929 = _T_137 ? 1'h0 : _GEN_56; // @[utils.scala 127:58 128:26]
  wire [4:0] _GEN_930 = _T_137 ? 5'h0 : _GEN_57; // @[utils.scala 127:58 129:25]
  wire [4:0] _GEN_931 = branchOps_passed ? _GEN_928 : _GEN_930; // @[utils.scala 121:32]
  wire  _GEN_932 = branchOps_passed ? readBuffer_branch_valid : _GEN_929; // @[utils.scala 121:32 125:24]
  wire [4:0] _GEN_933 = branchOps_valid ? _GEN_931 : _GEN_57; // @[utils.scala 120:29]
  wire  _GEN_934 = branchOps_valid ? _GEN_932 : _GEN_56; // @[utils.scala 120:29]
  wire [4:0] _T_156 = lastMissRecordRegister_branch_mask & branchOps_branchMask; // @[utils.scala 122:29]
  wire  _T_157 = |_T_156; // @[utils.scala 122:53]
  wire [4:0] _lastMissRecordRegister_branch_mask_T = lastMissRecordRegister_branch_mask ^ branchOps_branchMask; // @[utils.scala 123:40]
  wire [4:0] _GEN_939 = |_T_156 ? _lastMissRecordRegister_branch_mask_T : _GEN_891; // @[utils.scala 122:58 123:25]
  wire  _GEN_940 = _T_157 ? 1'h0 : _GEN_890; // @[utils.scala 127:58 128:26]
  wire [4:0] _GEN_941 = _T_157 ? 5'h0 : _GEN_891; // @[utils.scala 127:58 129:25]
  wire [4:0] _GEN_942 = branchOps_passed ? _GEN_939 : _GEN_941; // @[utils.scala 121:32]
  wire  _GEN_943 = branchOps_passed ? lastMissRecordRegister_branch_valid : _GEN_940; // @[utils.scala 121:32 125:24]
  wire [4:0] _GEN_944 = branchOps_valid ? _GEN_942 : _GEN_891; // @[utils.scala 120:29]
  wire  _GEN_945 = branchOps_valid ? _GEN_943 : _GEN_890; // @[utils.scala 120:29]
  wire [35:0] _GEN_32 = reset ? 36'h0 : _GEN_883; // @[cacheLookupUnit.scala 177:{32,32}]
  moduleForwardingMemory dataBRAM_0 ( // @[cacheLookupUnit.scala 60:39]
    .clock(dataBRAM_0_clock),
    .rdAddr(dataBRAM_0_rdAddr),
    .rdData(dataBRAM_0_rdData),
    .wrAddr(dataBRAM_0_wrAddr),
    .wrData(dataBRAM_0_wrData),
    .wrEna(dataBRAM_0_wrEna)
  );
  moduleForwardingMemory dataBRAM_1 ( // @[cacheLookupUnit.scala 60:39]
    .clock(dataBRAM_1_clock),
    .rdAddr(dataBRAM_1_rdAddr),
    .rdData(dataBRAM_1_rdData),
    .wrAddr(dataBRAM_1_wrAddr),
    .wrData(dataBRAM_1_wrData),
    .wrEna(dataBRAM_1_wrEna)
  );
  moduleForwardingMemory dataBRAM_2 ( // @[cacheLookupUnit.scala 60:39]
    .clock(dataBRAM_2_clock),
    .rdAddr(dataBRAM_2_rdAddr),
    .rdData(dataBRAM_2_rdData),
    .wrAddr(dataBRAM_2_wrAddr),
    .wrData(dataBRAM_2_wrData),
    .wrEna(dataBRAM_2_wrEna)
  );
  moduleForwardingMemory dataBRAM_3 ( // @[cacheLookupUnit.scala 60:39]
    .clock(dataBRAM_3_clock),
    .rdAddr(dataBRAM_3_rdAddr),
    .rdData(dataBRAM_3_rdData),
    .wrAddr(dataBRAM_3_wrAddr),
    .wrData(dataBRAM_3_wrData),
    .wrEna(dataBRAM_3_wrEna)
  );
  moduleForwardingMemory_4 tagBRAM ( // @[cacheLookupUnit.scala 110:23]
    .clock(tagBRAM_clock),
    .rdAddr(tagBRAM_rdAddr),
    .rdData(tagBRAM_rdData),
    .wrAddr(tagBRAM_wrAddr),
    .wrData(tagBRAM_wrData),
    .wrEna(tagBRAM_wrEna)
  );
  assign request_ready = toReplay_ready & toWriteBack_ready & toCoherency_ready; // @[cacheLookupUnit.scala 193:56]
  assign request_holdInOrder = lastMissRecordRegister_valid & lastMissRecordRegister_branch_valid & ~
    writeCommitInstructionBuffer; // @[cacheLookupUnit.scala 194:94]
  assign toReplay_request_valid = toReplay_ready & replayBuffer_valid; // @[cacheLookupUnit.scala 155:23 156:22 utils.scala 48:41]
  assign toReplay_request_address = toReplay_ready ? replayBuffer_address : 32'h0; // @[cacheLookupUnit.scala 155:23 156:22 utils.scala 49:41]
  assign toReplay_request_core_instruction = toReplay_ready ? replayBuffer_core_instruction : 32'h0; // @[cacheLookupUnit.scala 155:23 156:22 utils.scala 49:41]
  assign toReplay_request_core_robAddr = toReplay_ready ? replayBuffer_core_robAddr : 4'h0; // @[cacheLookupUnit.scala 155:23 156:22 utils.scala 49:41]
  assign toReplay_request_core_prfDest = toReplay_ready ? replayBuffer_core_prfDest : 6'h0; // @[cacheLookupUnit.scala 155:23 156:22 utils.scala 49:41]
  assign toReplay_request_branch_valid = toReplay_ready & replayBuffer_branch_valid; // @[cacheLookupUnit.scala 155:23 156:22 utils.scala 48:41]
  assign toReplay_request_branch_mask = toReplay_ready ? replayBuffer_branch_mask : 5'h0; // @[cacheLookupUnit.scala 155:23 156:22 utils.scala 49:41]
  assign toReplay_request_writeData_valid = toReplay_ready & replayBuffer_writeData_valid; // @[cacheLookupUnit.scala 155:23 156:22 utils.scala 48:41]
  assign toReplay_request_writeData_data = toReplay_ready ? replayBuffer_writeData_data : 64'h0; // @[cacheLookupUnit.scala 155:23 156:22 utils.scala 49:41]
  assign toReplay_request_cacheLine_response = toReplay_ready ? replayBuffer_cacheLine_response : 2'h0; // @[cacheLookupUnit.scala 155:23 156:22 utils.scala 49:41]
  assign toWriteBack_request_valid = toWriteBack_ready & writeBackBuffer_valid; // @[cacheLookupUnit.scala 179:26 180:25 utils.scala 48:41]
  assign toWriteBack_request_address = toWriteBack_ready ? writeBackBuffer_address : 32'h0; // @[cacheLookupUnit.scala 179:26 180:25 utils.scala 49:41]
  assign toWriteBack_request_data = toWriteBack_ready ? writeBackBuffer_data : 512'h0; // @[cacheLookupUnit.scala 179:26 180:25 utils.scala 49:41]
  assign toCoherency_request_valid = toCoherency_ready & coherencyResponseBuffer_valid; // @[cacheLookupUnit.scala 172:26 173:25 utils.scala 48:41]
  assign toCoherency_request_response = toCoherency_ready ? coherencyResponseBuffer_response : 2'h0; // @[cacheLookupUnit.scala 172:26 173:25 utils.scala 49:41]
  assign toCoherency_request_cacheLine = toCoherency_ready ? coherencyResponseBuffer_cacheLine : 512'h0; // @[cacheLookupUnit.scala 172:26 173:25 utils.scala 49:41]
  assign toCoherency_request_dataValid = toCoherency_ready & coherencyResponseBuffer_dataValid; // @[cacheLookupUnit.scala 172:26 173:25 utils.scala 48:41]
  assign toResponse_request_valid = memoryResponseBuffer_valid & memoryResponseBuffer_branch_valid &
    memoryResponseBuffer_valid; // @[cacheLookupUnit.scala 162:72 163:24 utils.scala 48:41]
  assign toResponse_request_address = memoryResponseBuffer_valid & memoryResponseBuffer_branch_valid ?
    memoryResponseBuffer_address : 32'h0; // @[cacheLookupUnit.scala 162:72 163:24 utils.scala 49:41]
  assign toResponse_request_core_instruction = memoryResponseBuffer_valid & memoryResponseBuffer_branch_valid ?
    memoryResponseBuffer_core_instruction : 32'h0; // @[cacheLookupUnit.scala 162:72 163:24 utils.scala 49:41]
  assign toResponse_request_core_robAddr = memoryResponseBuffer_valid & memoryResponseBuffer_branch_valid ?
    memoryResponseBuffer_core_robAddr : 4'h0; // @[cacheLookupUnit.scala 162:72 163:24 utils.scala 49:41]
  assign toResponse_request_core_prfDest = memoryResponseBuffer_valid & memoryResponseBuffer_branch_valid ?
    memoryResponseBuffer_core_prfDest : 6'h0; // @[cacheLookupUnit.scala 162:72 163:24 utils.scala 49:41]
  assign toResponse_request_branch_valid = memoryResponseBuffer_valid & memoryResponseBuffer_branch_valid & _GEN_21; // @[cacheLookupUnit.scala 162:72 utils.scala 48:41]
  assign toResponse_request_branch_mask = memoryResponseBuffer_valid & memoryResponseBuffer_branch_valid ? _GEN_20 : 5'h0
    ; // @[cacheLookupUnit.scala 162:72 utils.scala 49:41]
  assign toResponse_request_writeData_data = memoryResponseBuffer_valid & memoryResponseBuffer_branch_valid ?
    memoryResponseBuffer_writeData_data : 64'h0; // @[cacheLookupUnit.scala 162:72 163:24 utils.scala 49:41]
  assign writeInstructionCommit_ready = writeCommitInstructionBuffer; // @[cacheLookupUnit.scala 185:32]
  assign dataBRAM_0_clock = clock;
  assign dataBRAM_0_rdAddr = request_request_valid & request_request_branch_valid ? request_request_address[12:6] : 7'h0
    ; // @[cacheLookupUnit.scala 199:45 203:62 204:46]
  assign dataBRAM_0_wrAddr = operationValid ? _GEN_647 : 7'h0; // @[cacheLookupUnit.scala 212:23 75:28]
  assign dataBRAM_0_wrData = operationValid ? _GEN_643 : 512'h0; // @[cacheLookupUnit.scala 212:23 75:28]
  assign dataBRAM_0_wrEna = operationValid & _GEN_639; // @[cacheLookupUnit.scala 212:23 75:28]
  assign dataBRAM_1_clock = clock;
  assign dataBRAM_1_rdAddr = request_request_valid & request_request_branch_valid ? request_request_address[12:6] : 7'h0
    ; // @[cacheLookupUnit.scala 199:45 203:62 204:46]
  assign dataBRAM_1_wrAddr = operationValid ? _GEN_648 : 7'h0; // @[cacheLookupUnit.scala 212:23 75:28]
  assign dataBRAM_1_wrData = operationValid ? _GEN_644 : 512'h0; // @[cacheLookupUnit.scala 212:23 75:28]
  assign dataBRAM_1_wrEna = operationValid & _GEN_640; // @[cacheLookupUnit.scala 212:23 75:28]
  assign dataBRAM_2_clock = clock;
  assign dataBRAM_2_rdAddr = request_request_valid & request_request_branch_valid ? request_request_address[12:6] : 7'h0
    ; // @[cacheLookupUnit.scala 199:45 203:62 204:46]
  assign dataBRAM_2_wrAddr = operationValid ? _GEN_649 : 7'h0; // @[cacheLookupUnit.scala 212:23 75:28]
  assign dataBRAM_2_wrData = operationValid ? _GEN_645 : 512'h0; // @[cacheLookupUnit.scala 212:23 75:28]
  assign dataBRAM_2_wrEna = operationValid & _GEN_641; // @[cacheLookupUnit.scala 212:23 75:28]
  assign dataBRAM_3_clock = clock;
  assign dataBRAM_3_rdAddr = request_request_valid & request_request_branch_valid ? request_request_address[12:6] : 7'h0
    ; // @[cacheLookupUnit.scala 199:45 203:62 204:46]
  assign dataBRAM_3_wrAddr = operationValid ? _GEN_650 : 7'h0; // @[cacheLookupUnit.scala 212:23 75:28]
  assign dataBRAM_3_wrData = operationValid ? _GEN_646 : 512'h0; // @[cacheLookupUnit.scala 212:23 75:28]
  assign dataBRAM_3_wrEna = operationValid & _GEN_642; // @[cacheLookupUnit.scala 212:23 75:28]
  assign tagBRAM_clock = clock;
  assign tagBRAM_rdAddr = request_request_valid & request_request_branch_valid ? request_request_address[12:6] : 7'h0; // @[cacheLookupUnit.scala 200:18 203:62 205:20]
  assign tagBRAM_wrAddr = operationValid ? readBuffer_address[12:6] : 7'h0; // @[cacheLookupUnit.scala 118:18 212:23 406:20]
  assign tagBRAM_wrData = operationValid ? _tagBRAM_wrData_T_2 : 92'h0; // @[cacheLookupUnit.scala 116:18 212:23 405:20]
  assign tagBRAM_wrEna = operationValid & tagBRAMUpdateWire; // @[cacheLookupUnit.scala 117:18 212:23 404:19]
  always @(posedge clock) begin
    operationValid <= request_ready & request_request_valid & request_request_branch_valid; // @[cacheLookupUnit.scala 52:71]
    if (reset) begin // @[cacheLookupUnit.scala 121:36]
      reservationRegister_address <= 32'h0; // @[cacheLookupUnit.scala 121:36]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toReservationRegisterWire) begin // @[cacheLookupUnit.scala 537:36]
        reservationRegister_address <= readBuffer_address; // @[cacheLookupUnit.scala 539:35]
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 121:36]
      reservationRegister_reserved <= 1'h0; // @[cacheLookupUnit.scala 121:36]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toReservationRegisterWire) begin // @[cacheLookupUnit.scala 537:36]
        reservationRegister_reserved <= toReservationRegisterWire; // @[cacheLookupUnit.scala 538:36]
      end else if (isSCWriteWire) begin // @[cacheLookupUnit.scala 455:24]
        reservationRegister_reserved <= 1'h0; // @[cacheLookupUnit.scala 456:36]
      end else begin
        reservationRegister_reserved <= _GEN_630;
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 121:36]
      reservationRegister_size <= 1'h0; // @[cacheLookupUnit.scala 121:36]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toReservationRegisterWire) begin // @[cacheLookupUnit.scala 537:36]
        reservationRegister_size <= readBuffer_core_instruction[12]; // @[cacheLookupUnit.scala 540:32]
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 130:39]
      lastMissRecordRegister_valid <= 1'h0; // @[cacheLookupUnit.scala 130:39]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toLastMissRecordRegister & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 532:62]
        lastMissRecordRegister_valid <= readBuffer_valid; // @[cacheLookupUnit.scala 533:30]
      end else begin
        lastMissRecordRegister_valid <= _GEN_1;
      end
    end else begin
      lastMissRecordRegister_valid <= _GEN_1;
    end
    if (reset) begin // @[cacheLookupUnit.scala 130:39]
      lastMissRecordRegister_address <= 32'h0; // @[cacheLookupUnit.scala 130:39]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toLastMissRecordRegister & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 532:62]
        lastMissRecordRegister_address <= readBuffer_address; // @[cacheLookupUnit.scala 533:30]
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 130:39]
      lastMissRecordRegister_core_instruction <= 32'h0; // @[cacheLookupUnit.scala 130:39]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toLastMissRecordRegister & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 532:62]
        lastMissRecordRegister_core_instruction <= readBuffer_core_instruction; // @[cacheLookupUnit.scala 533:30]
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 130:39]
      lastMissRecordRegister_core_robAddr <= 4'h0; // @[cacheLookupUnit.scala 130:39]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toLastMissRecordRegister & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 532:62]
        lastMissRecordRegister_core_robAddr <= readBuffer_core_robAddr; // @[cacheLookupUnit.scala 533:30]
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 130:39]
      lastMissRecordRegister_core_prfDest <= 6'h0; // @[cacheLookupUnit.scala 130:39]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toLastMissRecordRegister & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 532:62]
        lastMissRecordRegister_core_prfDest <= readBuffer_core_prfDest; // @[cacheLookupUnit.scala 533:30]
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 130:39]
      lastMissRecordRegister_branch_valid <= 1'h0; // @[cacheLookupUnit.scala 130:39]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 545:23]
      lastMissRecordRegister_branch_valid <= _GEN_890;
    end else if (_request_holdInOrder_T) begin // @[cacheLookupUnit.scala 562:78]
      if (lastMissRecordRegister_branch_valid) begin // @[utils.scala 119:24]
        lastMissRecordRegister_branch_valid <= _GEN_945;
      end else begin
        lastMissRecordRegister_branch_valid <= _GEN_890;
      end
    end else begin
      lastMissRecordRegister_branch_valid <= _GEN_890;
    end
    if (reset) begin // @[cacheLookupUnit.scala 130:39]
      lastMissRecordRegister_branch_mask <= 5'h0; // @[cacheLookupUnit.scala 130:39]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 545:23]
      lastMissRecordRegister_branch_mask <= _GEN_891;
    end else if (_request_holdInOrder_T) begin // @[cacheLookupUnit.scala 562:78]
      if (lastMissRecordRegister_branch_valid) begin // @[utils.scala 119:24]
        lastMissRecordRegister_branch_mask <= _GEN_944;
      end else begin
        lastMissRecordRegister_branch_mask <= _GEN_891;
      end
    end else begin
      lastMissRecordRegister_branch_mask <= _GEN_891;
    end
    if (reset) begin // @[cacheLookupUnit.scala 146:27]
      readBuffer_valid <= 1'h0; // @[cacheLookupUnit.scala 146:27]
    end else begin
      readBuffer_valid <= _GEN_51;
    end
    if (reset) begin // @[cacheLookupUnit.scala 146:27]
      readBuffer_address <= 32'h0; // @[cacheLookupUnit.scala 146:27]
    end else if (request_request_valid & request_request_branch_valid) begin // @[cacheLookupUnit.scala 203:62]
      readBuffer_address <= request_request_address; // @[cacheLookupUnit.scala 207:16]
    end
    if (reset) begin // @[cacheLookupUnit.scala 146:27]
      readBuffer_core_instruction <= 32'h0; // @[cacheLookupUnit.scala 146:27]
    end else if (request_request_valid & request_request_branch_valid) begin // @[cacheLookupUnit.scala 203:62]
      readBuffer_core_instruction <= request_request_core_instruction; // @[cacheLookupUnit.scala 207:16]
    end
    if (reset) begin // @[cacheLookupUnit.scala 146:27]
      readBuffer_core_robAddr <= 4'h0; // @[cacheLookupUnit.scala 146:27]
    end else if (request_request_valid & request_request_branch_valid) begin // @[cacheLookupUnit.scala 203:62]
      readBuffer_core_robAddr <= request_request_core_robAddr; // @[cacheLookupUnit.scala 207:16]
    end
    if (reset) begin // @[cacheLookupUnit.scala 146:27]
      readBuffer_core_prfDest <= 6'h0; // @[cacheLookupUnit.scala 146:27]
    end else if (request_request_valid & request_request_branch_valid) begin // @[cacheLookupUnit.scala 203:62]
      readBuffer_core_prfDest <= request_request_core_prfDest; // @[cacheLookupUnit.scala 207:16]
    end
    if (reset) begin // @[cacheLookupUnit.scala 146:27]
      readBuffer_branch_valid <= 1'h0; // @[cacheLookupUnit.scala 146:27]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 545:23]
      readBuffer_branch_valid <= _GEN_56;
    end else if (readBuffer_valid & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 559:54]
      if (readBuffer_branch_valid) begin // @[utils.scala 119:24]
        readBuffer_branch_valid <= _GEN_934;
      end else begin
        readBuffer_branch_valid <= _GEN_56;
      end
    end else begin
      readBuffer_branch_valid <= _GEN_56;
    end
    if (reset) begin // @[cacheLookupUnit.scala 146:27]
      readBuffer_branch_mask <= 5'h0; // @[cacheLookupUnit.scala 146:27]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 545:23]
      readBuffer_branch_mask <= _GEN_57;
    end else if (readBuffer_valid & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 559:54]
      if (readBuffer_branch_valid) begin // @[utils.scala 119:24]
        readBuffer_branch_mask <= _GEN_933;
      end else begin
        readBuffer_branch_mask <= _GEN_57;
      end
    end else begin
      readBuffer_branch_mask <= _GEN_57;
    end
    if (reset) begin // @[cacheLookupUnit.scala 146:27]
      readBuffer_writeData_valid <= 1'h0; // @[cacheLookupUnit.scala 146:27]
    end else if (request_request_valid & request_request_branch_valid) begin // @[cacheLookupUnit.scala 203:62]
      readBuffer_writeData_valid <= request_request_writeData_valid; // @[cacheLookupUnit.scala 207:16]
    end
    if (reset) begin // @[cacheLookupUnit.scala 146:27]
      readBuffer_writeData_data <= 64'h0; // @[cacheLookupUnit.scala 146:27]
    end else if (request_request_valid & request_request_branch_valid) begin // @[cacheLookupUnit.scala 203:62]
      readBuffer_writeData_data <= request_request_writeData_data; // @[cacheLookupUnit.scala 207:16]
    end
    if (reset) begin // @[cacheLookupUnit.scala 146:27]
      readBuffer_cacheLine_cacheLine <= 512'h0; // @[cacheLookupUnit.scala 146:27]
    end else if (request_request_valid & request_request_branch_valid) begin // @[cacheLookupUnit.scala 203:62]
      readBuffer_cacheLine_cacheLine <= request_request_cacheLine_cacheLine; // @[cacheLookupUnit.scala 207:16]
    end
    if (reset) begin // @[cacheLookupUnit.scala 146:27]
      readBuffer_cacheLine_response <= 2'h0; // @[cacheLookupUnit.scala 146:27]
    end else if (request_request_valid & request_request_branch_valid) begin // @[cacheLookupUnit.scala 203:62]
      readBuffer_cacheLine_response <= request_request_cacheLine_response; // @[cacheLookupUnit.scala 207:16]
    end
    if (reset) begin // @[cacheLookupUnit.scala 147:28]
      requestType <= 2'h0; // @[cacheLookupUnit.scala 147:28]
    end else if (request_request_valid & request_request_branch_valid) begin // @[cacheLookupUnit.scala 203:62]
      requestType <= request_requestType; // @[cacheLookupUnit.scala 208:17]
    end
    if (reset) begin // @[cacheLookupUnit.scala 153:29]
      replayBuffer_valid <= 1'h0; // @[cacheLookupUnit.scala 153:29]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toReplayValidWire & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 499:55]
        replayBuffer_valid <= readBuffer_valid; // @[cacheLookupUnit.scala 500:20]
      end else begin
        replayBuffer_valid <= _GEN_14;
      end
    end else begin
      replayBuffer_valid <= _GEN_14;
    end
    if (reset) begin // @[cacheLookupUnit.scala 153:29]
      replayBuffer_address <= 32'h0; // @[cacheLookupUnit.scala 153:29]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toReplayValidWire & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 499:55]
        replayBuffer_address <= readBuffer_address; // @[cacheLookupUnit.scala 500:20]
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 153:29]
      replayBuffer_core_instruction <= 32'h0; // @[cacheLookupUnit.scala 153:29]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toReplayValidWire & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 499:55]
        replayBuffer_core_instruction <= readBuffer_core_instruction; // @[cacheLookupUnit.scala 500:20]
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 153:29]
      replayBuffer_core_robAddr <= 4'h0; // @[cacheLookupUnit.scala 153:29]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toReplayValidWire & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 499:55]
        replayBuffer_core_robAddr <= readBuffer_core_robAddr; // @[cacheLookupUnit.scala 500:20]
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 153:29]
      replayBuffer_core_prfDest <= 6'h0; // @[cacheLookupUnit.scala 153:29]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toReplayValidWire & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 499:55]
        replayBuffer_core_prfDest <= readBuffer_core_prfDest; // @[cacheLookupUnit.scala 500:20]
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 153:29]
      replayBuffer_branch_valid <= 1'h0; // @[cacheLookupUnit.scala 153:29]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 545:23]
      if (toReplayValidWire) begin // @[cacheLookupUnit.scala 546:28]
        if (branchOps_valid) begin // @[utils.scala 89:27]
          replayBuffer_branch_valid <= _GEN_903;
        end else begin
          replayBuffer_branch_valid <= readBuffer_branch_valid; // @[utils.scala 112:24]
        end
      end else begin
        replayBuffer_branch_valid <= _GEN_859;
      end
    end else if (replayBuffer_valid & ~toReplay_request_valid) begin // @[cacheLookupUnit.scala 555:56]
      if (replayBuffer_branch_valid) begin // @[utils.scala 119:24]
        replayBuffer_branch_valid <= _GEN_923;
      end else begin
        replayBuffer_branch_valid <= _GEN_859;
      end
    end else begin
      replayBuffer_branch_valid <= _GEN_859;
    end
    if (reset) begin // @[cacheLookupUnit.scala 153:29]
      replayBuffer_branch_mask <= 5'h0; // @[cacheLookupUnit.scala 153:29]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 545:23]
      if (toReplayValidWire) begin // @[cacheLookupUnit.scala 546:28]
        if (branchOps_valid) begin // @[utils.scala 89:27]
          replayBuffer_branch_mask <= _GEN_902;
        end else begin
          replayBuffer_branch_mask <= readBuffer_branch_mask; // @[utils.scala 111:23]
        end
      end else begin
        replayBuffer_branch_mask <= _GEN_860;
      end
    end else if (replayBuffer_valid & ~toReplay_request_valid) begin // @[cacheLookupUnit.scala 555:56]
      if (replayBuffer_branch_valid) begin // @[utils.scala 119:24]
        replayBuffer_branch_mask <= _GEN_922;
      end else begin
        replayBuffer_branch_mask <= _GEN_860;
      end
    end else begin
      replayBuffer_branch_mask <= _GEN_860;
    end
    if (reset) begin // @[cacheLookupUnit.scala 153:29]
      replayBuffer_writeData_valid <= 1'h0; // @[cacheLookupUnit.scala 153:29]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toReplayValidWire & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 499:55]
        replayBuffer_writeData_valid <= readBuffer_writeData_valid; // @[cacheLookupUnit.scala 500:20]
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 153:29]
      replayBuffer_writeData_data <= 64'h0; // @[cacheLookupUnit.scala 153:29]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toReplayValidWire & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 499:55]
        replayBuffer_writeData_data <= readBuffer_writeData_data; // @[cacheLookupUnit.scala 500:20]
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 153:29]
      replayBuffer_cacheLine_response <= 2'h0; // @[cacheLookupUnit.scala 153:29]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toReplayValidWire & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 499:55]
        if (_T_14) begin // @[cacheLookupUnit.scala 442:43]
          replayBuffer_cacheLine_response <= _GEN_683;
        end else begin
          replayBuffer_cacheLine_response <= _GEN_673;
        end
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 160:37]
      memoryResponseBuffer_valid <= 1'h0; // @[cacheLookupUnit.scala 160:37]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toMemoryResponseValidWire & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 506:63]
        memoryResponseBuffer_valid <= readBuffer_valid; // @[cacheLookupUnit.scala 507:28]
      end else begin
        memoryResponseBuffer_valid <= _GEN_34;
      end
    end else begin
      memoryResponseBuffer_valid <= _GEN_34;
    end
    if (reset) begin // @[cacheLookupUnit.scala 160:37]
      memoryResponseBuffer_address <= 32'h0; // @[cacheLookupUnit.scala 160:37]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toMemoryResponseValidWire & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 506:63]
        memoryResponseBuffer_address <= readBuffer_address; // @[cacheLookupUnit.scala 507:28]
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 160:37]
      memoryResponseBuffer_core_instruction <= 32'h0; // @[cacheLookupUnit.scala 160:37]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toMemoryResponseValidWire & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 506:63]
        memoryResponseBuffer_core_instruction <= readBuffer_core_instruction; // @[cacheLookupUnit.scala 507:28]
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 160:37]
      memoryResponseBuffer_core_robAddr <= 4'h0; // @[cacheLookupUnit.scala 160:37]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toMemoryResponseValidWire & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 506:63]
        memoryResponseBuffer_core_robAddr <= readBuffer_core_robAddr; // @[cacheLookupUnit.scala 507:28]
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 160:37]
      memoryResponseBuffer_core_prfDest <= 6'h0; // @[cacheLookupUnit.scala 160:37]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toMemoryResponseValidWire & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 506:63]
        memoryResponseBuffer_core_prfDest <= readBuffer_core_prfDest; // @[cacheLookupUnit.scala 507:28]
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 160:37]
      memoryResponseBuffer_branch_valid <= 1'h0; // @[cacheLookupUnit.scala 160:37]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 545:23]
      if (toMemoryResponseValidWire) begin // @[cacheLookupUnit.scala 549:36]
        if (branchOps_valid) begin // @[utils.scala 89:27]
          memoryResponseBuffer_branch_valid <= _GEN_903;
        end else begin
          memoryResponseBuffer_branch_valid <= readBuffer_branch_valid; // @[utils.scala 112:24]
        end
      end else begin
        memoryResponseBuffer_branch_valid <= _GEN_871;
      end
    end else begin
      memoryResponseBuffer_branch_valid <= _GEN_871;
    end
    if (reset) begin // @[cacheLookupUnit.scala 160:37]
      memoryResponseBuffer_branch_mask <= 5'h0; // @[cacheLookupUnit.scala 160:37]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 545:23]
      if (toMemoryResponseValidWire) begin // @[cacheLookupUnit.scala 549:36]
        if (branchOps_valid) begin // @[utils.scala 89:27]
          memoryResponseBuffer_branch_mask <= _GEN_902;
        end else begin
          memoryResponseBuffer_branch_mask <= readBuffer_branch_mask; // @[utils.scala 111:23]
        end
      end else begin
        memoryResponseBuffer_branch_mask <= _GEN_872;
      end
    end else begin
      memoryResponseBuffer_branch_mask <= _GEN_872;
    end
    if (reset) begin // @[cacheLookupUnit.scala 160:37]
      memoryResponseBuffer_writeData_data <= 64'h0; // @[cacheLookupUnit.scala 160:37]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toMemoryResponseValidWire & readBuffer_branch_valid) begin // @[cacheLookupUnit.scala 506:63]
        if (isSCReadWire) begin // @[cacheLookupUnit.scala 493:23]
          memoryResponseBuffer_writeData_data <= {{63'd0}, _responseResultWire_T_21}; // @[cacheLookupUnit.scala 494:26]
        end else begin
          memoryResponseBuffer_writeData_data <= _GEN_768;
        end
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 170:40]
      coherencyResponseBuffer_valid <= 1'h0; // @[cacheLookupUnit.scala 170:40]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toCoherencyResponseValidWire) begin // @[cacheLookupUnit.scala 512:39]
        coherencyResponseBuffer_valid <= toCoherencyResponseValidWire; // @[cacheLookupUnit.scala 513:37]
      end else begin
        coherencyResponseBuffer_valid <= _GEN_40;
      end
    end else begin
      coherencyResponseBuffer_valid <= _GEN_40;
    end
    if (reset) begin // @[cacheLookupUnit.scala 170:40]
      coherencyResponseBuffer_response <= 2'h0; // @[cacheLookupUnit.scala 170:40]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toCoherencyResponseValidWire) begin // @[cacheLookupUnit.scala 512:39]
        if (readBuffer_cacheLine_response[0]) begin // @[cacheLookupUnit.scala 514:45]
          coherencyResponseBuffer_response <= _coherencyResponseBuffer_response_T_3; // @[cacheLookupUnit.scala 517:42]
        end
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 170:40]
      coherencyResponseBuffer_cacheLine <= 512'h0; // @[cacheLookupUnit.scala 170:40]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toCoherencyResponseValidWire) begin // @[cacheLookupUnit.scala 512:39]
        if (readBuffer_cacheLine_response[0]) begin // @[cacheLookupUnit.scala 514:45]
          coherencyResponseBuffer_cacheLine <= _coherencyResponseBuffer_cacheLine_T_3; // @[cacheLookupUnit.scala 515:43]
        end else begin
          coherencyResponseBuffer_cacheLine <= 512'h0; // @[cacheLookupUnit.scala 519:43]
        end
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 170:40]
      coherencyResponseBuffer_dataValid <= 1'h0; // @[cacheLookupUnit.scala 170:40]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toCoherencyResponseValidWire) begin // @[cacheLookupUnit.scala 512:39]
        coherencyResponseBuffer_dataValid <= _newShareBitWire_T_9;
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 177:32]
      writeBackBuffer_valid <= 1'h0; // @[cacheLookupUnit.scala 177:32]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toWriteBackValidWire) begin // @[cacheLookupUnit.scala 525:31]
        writeBackBuffer_valid <= toWriteBackValidWire; // @[cacheLookupUnit.scala 526:29]
      end else begin
        writeBackBuffer_valid <= _GEN_44;
      end
    end else begin
      writeBackBuffer_valid <= _GEN_44;
    end
    writeBackBuffer_address <= _GEN_32[31:0]; // @[cacheLookupUnit.scala 177:{32,32}]
    if (reset) begin // @[cacheLookupUnit.scala 177:32]
      writeBackBuffer_data <= 512'h0; // @[cacheLookupUnit.scala 177:32]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      if (toWriteBackValidWire) begin // @[cacheLookupUnit.scala 525:31]
        if (2'h3 == updatingSet) begin // @[cacheLookupUnit.scala 528:28]
          writeBackBuffer_data <= dataBRAMVec_3_rdData; // @[cacheLookupUnit.scala 528:28]
        end else begin
          writeBackBuffer_data <= _GEN_811;
        end
      end
    end
    if (reset) begin // @[cacheLookupUnit.scala 184:45]
      writeCommitInstructionBuffer <= 1'h0; // @[cacheLookupUnit.scala 184:45]
    end else if (operationValid) begin // @[cacheLookupUnit.scala 212:23]
      writeCommitInstructionBuffer <= _GEN_700;
    end else if (writeInstructionCommit_fired) begin // @[cacheLookupUnit.scala 186:37]
      writeCommitInstructionBuffer <= 1'h0; // @[cacheLookupUnit.scala 187:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  operationValid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reservationRegister_address = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reservationRegister_reserved = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  reservationRegister_size = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  lastMissRecordRegister_valid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lastMissRecordRegister_address = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  lastMissRecordRegister_core_instruction = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  lastMissRecordRegister_core_robAddr = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  lastMissRecordRegister_core_prfDest = _RAND_8[5:0];
  _RAND_9 = {1{`RANDOM}};
  lastMissRecordRegister_branch_valid = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  lastMissRecordRegister_branch_mask = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  readBuffer_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  readBuffer_address = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  readBuffer_core_instruction = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  readBuffer_core_robAddr = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  readBuffer_core_prfDest = _RAND_15[5:0];
  _RAND_16 = {1{`RANDOM}};
  readBuffer_branch_valid = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  readBuffer_branch_mask = _RAND_17[4:0];
  _RAND_18 = {1{`RANDOM}};
  readBuffer_writeData_valid = _RAND_18[0:0];
  _RAND_19 = {2{`RANDOM}};
  readBuffer_writeData_data = _RAND_19[63:0];
  _RAND_20 = {16{`RANDOM}};
  readBuffer_cacheLine_cacheLine = _RAND_20[511:0];
  _RAND_21 = {1{`RANDOM}};
  readBuffer_cacheLine_response = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  requestType = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  replayBuffer_valid = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  replayBuffer_address = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  replayBuffer_core_instruction = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  replayBuffer_core_robAddr = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  replayBuffer_core_prfDest = _RAND_27[5:0];
  _RAND_28 = {1{`RANDOM}};
  replayBuffer_branch_valid = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  replayBuffer_branch_mask = _RAND_29[4:0];
  _RAND_30 = {1{`RANDOM}};
  replayBuffer_writeData_valid = _RAND_30[0:0];
  _RAND_31 = {2{`RANDOM}};
  replayBuffer_writeData_data = _RAND_31[63:0];
  _RAND_32 = {1{`RANDOM}};
  replayBuffer_cacheLine_response = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  memoryResponseBuffer_valid = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  memoryResponseBuffer_address = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  memoryResponseBuffer_core_instruction = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  memoryResponseBuffer_core_robAddr = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  memoryResponseBuffer_core_prfDest = _RAND_37[5:0];
  _RAND_38 = {1{`RANDOM}};
  memoryResponseBuffer_branch_valid = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  memoryResponseBuffer_branch_mask = _RAND_39[4:0];
  _RAND_40 = {2{`RANDOM}};
  memoryResponseBuffer_writeData_data = _RAND_40[63:0];
  _RAND_41 = {1{`RANDOM}};
  coherencyResponseBuffer_valid = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  coherencyResponseBuffer_response = _RAND_42[1:0];
  _RAND_43 = {16{`RANDOM}};
  coherencyResponseBuffer_cacheLine = _RAND_43[511:0];
  _RAND_44 = {1{`RANDOM}};
  coherencyResponseBuffer_dataValid = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  writeBackBuffer_valid = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  writeBackBuffer_address = _RAND_46[31:0];
  _RAND_47 = {16{`RANDOM}};
  writeBackBuffer_data = _RAND_47[511:0];
  _RAND_48 = {1{`RANDOM}};
  writeCommitInstructionBuffer = _RAND_48[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module fifoBypassModule(
  input          clock,
  input          reset,
  output         write_ready,
  input          write_data_valid,
  input  [31:0]  write_data_address,
  input  [511:0] write_data_data,
  input          read_ready,
  output         read_data_valid,
  output [31:0]  read_data_address,
  output [511:0] read_data_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [511:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [511:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [511:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [511:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [511:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [511:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [511:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [511:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [511:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [511:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [511:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [511:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [511:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [511:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [511:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [511:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] memReg_0_address; // @[fifo.scala 179:33]
  reg [511:0] memReg_0_data; // @[fifo.scala 179:33]
  reg [31:0] memReg_1_address; // @[fifo.scala 179:33]
  reg [511:0] memReg_1_data; // @[fifo.scala 179:33]
  reg [31:0] memReg_2_address; // @[fifo.scala 179:33]
  reg [511:0] memReg_2_data; // @[fifo.scala 179:33]
  reg [31:0] memReg_3_address; // @[fifo.scala 179:33]
  reg [511:0] memReg_3_data; // @[fifo.scala 179:33]
  reg [31:0] memReg_4_address; // @[fifo.scala 179:33]
  reg [511:0] memReg_4_data; // @[fifo.scala 179:33]
  reg [31:0] memReg_5_address; // @[fifo.scala 179:33]
  reg [511:0] memReg_5_data; // @[fifo.scala 179:33]
  reg [31:0] memReg_6_address; // @[fifo.scala 179:33]
  reg [511:0] memReg_6_data; // @[fifo.scala 179:33]
  reg [31:0] memReg_7_address; // @[fifo.scala 179:33]
  reg [511:0] memReg_7_data; // @[fifo.scala 179:33]
  reg [31:0] memReg_8_address; // @[fifo.scala 179:33]
  reg [511:0] memReg_8_data; // @[fifo.scala 179:33]
  reg [31:0] memReg_9_address; // @[fifo.scala 179:33]
  reg [511:0] memReg_9_data; // @[fifo.scala 179:33]
  reg [31:0] memReg_10_address; // @[fifo.scala 179:33]
  reg [511:0] memReg_10_data; // @[fifo.scala 179:33]
  reg [31:0] memReg_11_address; // @[fifo.scala 179:33]
  reg [511:0] memReg_11_data; // @[fifo.scala 179:33]
  reg [31:0] memReg_12_address; // @[fifo.scala 179:33]
  reg [511:0] memReg_12_data; // @[fifo.scala 179:33]
  reg [31:0] memReg_13_address; // @[fifo.scala 179:33]
  reg [511:0] memReg_13_data; // @[fifo.scala 179:33]
  reg [31:0] memReg_14_address; // @[fifo.scala 179:33]
  reg [511:0] memReg_14_data; // @[fifo.scala 179:33]
  reg [31:0] memReg_15_address; // @[fifo.scala 179:33]
  reg [511:0] memReg_15_data; // @[fifo.scala 179:33]
  reg [3:0] readPtr; // @[fifo.scala 185:25]
  wire [3:0] _nextVal_T_2 = readPtr + 4'h1; // @[fifo.scala 186:60]
  wire [3:0] nextRead = readPtr == 4'hf ? 4'h0 : _nextVal_T_2; // @[fifo.scala 186:22]
  reg  emptyReg; // @[fifo.scala 194:25]
  wire [1:0] op = {write_data_valid,read_ready}; // @[fifo.scala 197:29]
  wire  bypass = emptyReg & op == 2'h3; // @[fifo.scala 198:25]
  wire  _T_2 = ~emptyReg; // @[fifo.scala 204:12]
  wire  _GEN_21 = 2'h2 == op ? 1'h0 : 2'h3 == op & _T_2; // @[fifo.scala 201:14]
  wire  _GEN_24 = 2'h1 == op ? _T_2 : _GEN_21; // @[fifo.scala 201:14]
  wire  _GEN_28 = 2'h0 == op ? 1'h0 : _GEN_24; // @[fifo.scala 201:14]
  wire  incrRead = bypass ? 1'h0 : _GEN_28; // @[fifo.scala 234:16 236:14]
  reg [3:0] writePtr; // @[fifo.scala 185:25]
  wire [3:0] _nextVal_T_5 = writePtr + 4'h1; // @[fifo.scala 186:60]
  wire [3:0] nextWrite = writePtr == 4'hf ? 4'h0 : _nextVal_T_5; // @[fifo.scala 186:22]
  reg  fullReg; // @[fifo.scala 195:34]
  wire  _T_4 = ~fullReg; // @[fifo.scala 211:12]
  wire  _GEN_18 = 2'h2 == op ? _T_4 : 2'h3 == op & _T_4; // @[fifo.scala 201:14]
  wire  _GEN_25 = 2'h1 == op ? 1'h0 : _GEN_18; // @[fifo.scala 201:14]
  wire  _GEN_29 = 2'h0 == op ? 1'h0 : _GEN_25; // @[fifo.scala 201:14]
  wire  incrWrite = bypass ? 1'h0 : _GEN_29; // @[fifo.scala 234:16 235:13]
  wire  _GEN_2 = ~emptyReg ? 1'h0 : fullReg; // @[fifo.scala 204:23 205:17 195:34]
  wire  _GEN_3 = ~emptyReg ? nextRead == writePtr : emptyReg; // @[fifo.scala 204:23 206:18 194:25]
  wire  _GEN_6 = ~fullReg ? 1'h0 : emptyReg; // @[fifo.scala 211:22 213:18 194:25]
  wire  _GEN_7 = ~fullReg ? nextWrite == readPtr : fullReg; // @[fifo.scala 211:22 214:17 195:34]
  wire  _fullReg_T_2 = emptyReg ? 1'h0 : nextWrite == nextRead; // @[fifo.scala 222:23]
  wire  _GEN_10 = _T_4 ? _fullReg_T_2 : fullReg; // @[fifo.scala 219:22 222:17 195:34]
  wire  _emptyReg_T_2 = fullReg ? 1'h0 : nextRead == nextWrite; // @[fifo.scala 227:24]
  wire  _GEN_11 = _T_2 ? 1'h0 : _GEN_10; // @[fifo.scala 225:23 226:17]
  wire  _GEN_12 = _T_2 ? _emptyReg_T_2 : _GEN_6; // @[fifo.scala 225:23 227:18]
  wire  _GEN_15 = 2'h3 == op ? _GEN_12 : emptyReg; // @[fifo.scala 201:14 194:25]
  wire  _GEN_16 = 2'h3 == op ? _GEN_11 : fullReg; // @[fifo.scala 201:14 195:34]
  wire  _GEN_19 = 2'h2 == op ? _GEN_6 : _GEN_15; // @[fifo.scala 201:14]
  wire  _GEN_20 = 2'h2 == op ? _GEN_7 : _GEN_16; // @[fifo.scala 201:14]
  wire  _GEN_23 = 2'h1 == op ? _GEN_3 : _GEN_19; // @[fifo.scala 201:14]
  wire  _GEN_27 = 2'h0 == op ? emptyReg : _GEN_23; // @[fifo.scala 201:14 194:25]
  wire  _GEN_32 = bypass | _GEN_27; // @[fifo.scala 234:16 238:14]
  wire [31:0] _GEN_134 = 4'h1 == readPtr ? memReg_1_address : memReg_0_address; // @[fifo.scala 247:{19,19}]
  wire [511:0] _GEN_135 = 4'h1 == readPtr ? memReg_1_data : memReg_0_data; // @[fifo.scala 247:{19,19}]
  wire [31:0] _GEN_137 = 4'h2 == readPtr ? memReg_2_address : _GEN_134; // @[fifo.scala 247:{19,19}]
  wire [511:0] _GEN_138 = 4'h2 == readPtr ? memReg_2_data : _GEN_135; // @[fifo.scala 247:{19,19}]
  wire [31:0] _GEN_140 = 4'h3 == readPtr ? memReg_3_address : _GEN_137; // @[fifo.scala 247:{19,19}]
  wire [511:0] _GEN_141 = 4'h3 == readPtr ? memReg_3_data : _GEN_138; // @[fifo.scala 247:{19,19}]
  wire [31:0] _GEN_143 = 4'h4 == readPtr ? memReg_4_address : _GEN_140; // @[fifo.scala 247:{19,19}]
  wire [511:0] _GEN_144 = 4'h4 == readPtr ? memReg_4_data : _GEN_141; // @[fifo.scala 247:{19,19}]
  wire [31:0] _GEN_146 = 4'h5 == readPtr ? memReg_5_address : _GEN_143; // @[fifo.scala 247:{19,19}]
  wire [511:0] _GEN_147 = 4'h5 == readPtr ? memReg_5_data : _GEN_144; // @[fifo.scala 247:{19,19}]
  wire [31:0] _GEN_149 = 4'h6 == readPtr ? memReg_6_address : _GEN_146; // @[fifo.scala 247:{19,19}]
  wire [511:0] _GEN_150 = 4'h6 == readPtr ? memReg_6_data : _GEN_147; // @[fifo.scala 247:{19,19}]
  wire [31:0] _GEN_152 = 4'h7 == readPtr ? memReg_7_address : _GEN_149; // @[fifo.scala 247:{19,19}]
  wire [511:0] _GEN_153 = 4'h7 == readPtr ? memReg_7_data : _GEN_150; // @[fifo.scala 247:{19,19}]
  wire [31:0] _GEN_155 = 4'h8 == readPtr ? memReg_8_address : _GEN_152; // @[fifo.scala 247:{19,19}]
  wire [511:0] _GEN_156 = 4'h8 == readPtr ? memReg_8_data : _GEN_153; // @[fifo.scala 247:{19,19}]
  wire [31:0] _GEN_158 = 4'h9 == readPtr ? memReg_9_address : _GEN_155; // @[fifo.scala 247:{19,19}]
  wire [511:0] _GEN_159 = 4'h9 == readPtr ? memReg_9_data : _GEN_156; // @[fifo.scala 247:{19,19}]
  wire [31:0] _GEN_161 = 4'ha == readPtr ? memReg_10_address : _GEN_158; // @[fifo.scala 247:{19,19}]
  wire [511:0] _GEN_162 = 4'ha == readPtr ? memReg_10_data : _GEN_159; // @[fifo.scala 247:{19,19}]
  wire [31:0] _GEN_164 = 4'hb == readPtr ? memReg_11_address : _GEN_161; // @[fifo.scala 247:{19,19}]
  wire [511:0] _GEN_165 = 4'hb == readPtr ? memReg_11_data : _GEN_162; // @[fifo.scala 247:{19,19}]
  wire [31:0] _GEN_167 = 4'hc == readPtr ? memReg_12_address : _GEN_164; // @[fifo.scala 247:{19,19}]
  wire [511:0] _GEN_168 = 4'hc == readPtr ? memReg_12_data : _GEN_165; // @[fifo.scala 247:{19,19}]
  wire [31:0] _GEN_170 = 4'hd == readPtr ? memReg_13_address : _GEN_167; // @[fifo.scala 247:{19,19}]
  wire [511:0] _GEN_171 = 4'hd == readPtr ? memReg_13_data : _GEN_168; // @[fifo.scala 247:{19,19}]
  wire [31:0] _GEN_173 = 4'he == readPtr ? memReg_14_address : _GEN_170; // @[fifo.scala 247:{19,19}]
  wire [511:0] _GEN_174 = 4'he == readPtr ? memReg_14_data : _GEN_171; // @[fifo.scala 247:{19,19}]
  wire [31:0] _GEN_176 = 4'hf == readPtr ? memReg_15_address : _GEN_173; // @[fifo.scala 247:{19,19}]
  wire [511:0] _GEN_177 = 4'hf == readPtr ? memReg_15_data : _GEN_174; // @[fifo.scala 247:{19,19}]
  assign write_ready = ~fullReg; // @[fifo.scala 249:18]
  assign read_data_valid = bypass | _T_2; // @[fifo.scala 248:25]
  assign read_data_address = bypass ? write_data_address : _GEN_176; // @[fifo.scala 247:19]
  assign read_data_data = bypass ? write_data_data : _GEN_177; // @[fifo.scala 247:19]
  always @(posedge clock) begin
    if (reset) begin // @[fifo.scala 179:33]
      memReg_0_address <= 32'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 243:22]
        memReg_0_address <= write_data_address; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_0_data <= 512'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 243:22]
        memReg_0_data <= write_data_data; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_1_address <= 32'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 243:22]
        memReg_1_address <= write_data_address; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_1_data <= 512'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 243:22]
        memReg_1_data <= write_data_data; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_2_address <= 32'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 243:22]
        memReg_2_address <= write_data_address; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_2_data <= 512'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 243:22]
        memReg_2_data <= write_data_data; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_3_address <= 32'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 243:22]
        memReg_3_address <= write_data_address; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_3_data <= 512'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 243:22]
        memReg_3_data <= write_data_data; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_4_address <= 32'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 243:22]
        memReg_4_address <= write_data_address; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_4_data <= 512'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 243:22]
        memReg_4_data <= write_data_data; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_5_address <= 32'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 243:22]
        memReg_5_address <= write_data_address; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_5_data <= 512'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 243:22]
        memReg_5_data <= write_data_data; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_6_address <= 32'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 243:22]
        memReg_6_address <= write_data_address; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_6_data <= 512'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 243:22]
        memReg_6_data <= write_data_data; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_7_address <= 32'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 243:22]
        memReg_7_address <= write_data_address; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_7_data <= 512'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 243:22]
        memReg_7_data <= write_data_data; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_8_address <= 32'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 243:22]
        memReg_8_address <= write_data_address; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_8_data <= 512'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 243:22]
        memReg_8_data <= write_data_data; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_9_address <= 32'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 243:22]
        memReg_9_address <= write_data_address; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_9_data <= 512'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 243:22]
        memReg_9_data <= write_data_data; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_10_address <= 32'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'ha == writePtr) begin // @[fifo.scala 243:22]
        memReg_10_address <= write_data_address; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_10_data <= 512'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'ha == writePtr) begin // @[fifo.scala 243:22]
        memReg_10_data <= write_data_data; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_11_address <= 32'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'hb == writePtr) begin // @[fifo.scala 243:22]
        memReg_11_address <= write_data_address; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_11_data <= 512'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'hb == writePtr) begin // @[fifo.scala 243:22]
        memReg_11_data <= write_data_data; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_12_address <= 32'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'hc == writePtr) begin // @[fifo.scala 243:22]
        memReg_12_address <= write_data_address; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_12_data <= 512'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'hc == writePtr) begin // @[fifo.scala 243:22]
        memReg_12_data <= write_data_data; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_13_address <= 32'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'hd == writePtr) begin // @[fifo.scala 243:22]
        memReg_13_address <= write_data_address; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_13_data <= 512'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'hd == writePtr) begin // @[fifo.scala 243:22]
        memReg_13_data <= write_data_data; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_14_address <= 32'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'he == writePtr) begin // @[fifo.scala 243:22]
        memReg_14_address <= write_data_address; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_14_data <= 512'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'he == writePtr) begin // @[fifo.scala 243:22]
        memReg_14_data <= write_data_data; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_15_address <= 32'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'hf == writePtr) begin // @[fifo.scala 243:22]
        memReg_15_address <= write_data_address; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 179:33]
      memReg_15_data <= 512'h0; // @[fifo.scala 179:33]
    end else if (incrWrite) begin // @[fifo.scala 242:17]
      if (4'hf == writePtr) begin // @[fifo.scala 243:22]
        memReg_15_data <= write_data_data; // @[fifo.scala 243:22]
      end
    end
    if (reset) begin // @[fifo.scala 185:25]
      readPtr <= 4'h0; // @[fifo.scala 185:25]
    end else if (incrRead) begin // @[fifo.scala 187:15]
      if (readPtr == 4'hf) begin // @[fifo.scala 186:22]
        readPtr <= 4'h0;
      end else begin
        readPtr <= _nextVal_T_2;
      end
    end
    emptyReg <= reset | _GEN_32; // @[fifo.scala 194:{25,25}]
    if (reset) begin // @[fifo.scala 185:25]
      writePtr <= 4'h0; // @[fifo.scala 185:25]
    end else if (incrWrite) begin // @[fifo.scala 187:15]
      if (writePtr == 4'hf) begin // @[fifo.scala 186:22]
        writePtr <= 4'h0;
      end else begin
        writePtr <= _nextVal_T_5;
      end
    end
    if (reset) begin // @[fifo.scala 195:34]
      fullReg <= 1'h0; // @[fifo.scala 195:34]
    end else if (bypass) begin // @[fifo.scala 234:16]
      fullReg <= 1'h0; // @[fifo.scala 239:13]
    end else if (!(2'h0 == op)) begin // @[fifo.scala 201:14]
      if (2'h1 == op) begin // @[fifo.scala 201:14]
        fullReg <= _GEN_2;
      end else begin
        fullReg <= _GEN_20;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  memReg_0_address = _RAND_0[31:0];
  _RAND_1 = {16{`RANDOM}};
  memReg_0_data = _RAND_1[511:0];
  _RAND_2 = {1{`RANDOM}};
  memReg_1_address = _RAND_2[31:0];
  _RAND_3 = {16{`RANDOM}};
  memReg_1_data = _RAND_3[511:0];
  _RAND_4 = {1{`RANDOM}};
  memReg_2_address = _RAND_4[31:0];
  _RAND_5 = {16{`RANDOM}};
  memReg_2_data = _RAND_5[511:0];
  _RAND_6 = {1{`RANDOM}};
  memReg_3_address = _RAND_6[31:0];
  _RAND_7 = {16{`RANDOM}};
  memReg_3_data = _RAND_7[511:0];
  _RAND_8 = {1{`RANDOM}};
  memReg_4_address = _RAND_8[31:0];
  _RAND_9 = {16{`RANDOM}};
  memReg_4_data = _RAND_9[511:0];
  _RAND_10 = {1{`RANDOM}};
  memReg_5_address = _RAND_10[31:0];
  _RAND_11 = {16{`RANDOM}};
  memReg_5_data = _RAND_11[511:0];
  _RAND_12 = {1{`RANDOM}};
  memReg_6_address = _RAND_12[31:0];
  _RAND_13 = {16{`RANDOM}};
  memReg_6_data = _RAND_13[511:0];
  _RAND_14 = {1{`RANDOM}};
  memReg_7_address = _RAND_14[31:0];
  _RAND_15 = {16{`RANDOM}};
  memReg_7_data = _RAND_15[511:0];
  _RAND_16 = {1{`RANDOM}};
  memReg_8_address = _RAND_16[31:0];
  _RAND_17 = {16{`RANDOM}};
  memReg_8_data = _RAND_17[511:0];
  _RAND_18 = {1{`RANDOM}};
  memReg_9_address = _RAND_18[31:0];
  _RAND_19 = {16{`RANDOM}};
  memReg_9_data = _RAND_19[511:0];
  _RAND_20 = {1{`RANDOM}};
  memReg_10_address = _RAND_20[31:0];
  _RAND_21 = {16{`RANDOM}};
  memReg_10_data = _RAND_21[511:0];
  _RAND_22 = {1{`RANDOM}};
  memReg_11_address = _RAND_22[31:0];
  _RAND_23 = {16{`RANDOM}};
  memReg_11_data = _RAND_23[511:0];
  _RAND_24 = {1{`RANDOM}};
  memReg_12_address = _RAND_24[31:0];
  _RAND_25 = {16{`RANDOM}};
  memReg_12_data = _RAND_25[511:0];
  _RAND_26 = {1{`RANDOM}};
  memReg_13_address = _RAND_26[31:0];
  _RAND_27 = {16{`RANDOM}};
  memReg_13_data = _RAND_27[511:0];
  _RAND_28 = {1{`RANDOM}};
  memReg_14_address = _RAND_28[31:0];
  _RAND_29 = {16{`RANDOM}};
  memReg_14_data = _RAND_29[511:0];
  _RAND_30 = {1{`RANDOM}};
  memReg_15_address = _RAND_30[31:0];
  _RAND_31 = {16{`RANDOM}};
  memReg_15_data = _RAND_31[511:0];
  _RAND_32 = {1{`RANDOM}};
  readPtr = _RAND_32[3:0];
  _RAND_33 = {1{`RANDOM}};
  emptyReg = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  writePtr = _RAND_34[3:0];
  _RAND_35 = {1{`RANDOM}};
  fullReg = _RAND_35[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module replayUnit(
  input          clock,
  input          reset,
  output         requestIn_ready,
  input          requestIn_request_valid,
  input  [31:0]  requestIn_request_address,
  input  [31:0]  requestIn_request_core_instruction,
  input  [3:0]   requestIn_request_core_robAddr,
  input  [5:0]   requestIn_request_core_prfDest,
  input          requestIn_request_branch_valid,
  input  [4:0]   requestIn_request_branch_mask,
  input          requestIn_request_writeData_valid,
  input  [63:0]  requestIn_request_writeData_data,
  input  [1:0]   requestIn_request_cacheLine_response,
  input          requestOut_ready,
  output         requestOut_request_valid,
  output [31:0]  requestOut_request_address,
  output [31:0]  requestOut_request_core_instruction,
  output [3:0]   requestOut_request_core_robAddr,
  output [5:0]   requestOut_request_core_prfDest,
  output         requestOut_request_branch_valid,
  output [4:0]   requestOut_request_branch_mask,
  output         requestOut_request_writeData_valid,
  output [63:0]  requestOut_request_writeData_data,
  output [1:0]   requestOut_request_cacheLine_response,
  output         responseIn_ready,
  input          responseIn_request_valid,
  input  [31:0]  responseIn_request_address,
  input  [31:0]  responseIn_request_core_instruction,
  input  [3:0]   responseIn_request_core_robAddr,
  input  [5:0]   responseIn_request_core_prfDest,
  input          responseIn_request_branch_valid,
  input  [4:0]   responseIn_request_branch_mask,
  input          responseIn_request_writeData_valid,
  input  [63:0]  responseIn_request_writeData_data,
  input  [511:0] responseIn_request_cacheLine_cacheLine,
  input  [1:0]   responseIn_request_cacheLine_response,
  input          responseOut_ready,
  output         responseOut_request_valid,
  output [31:0]  responseOut_request_address,
  output [31:0]  responseOut_request_core_instruction,
  output [3:0]   responseOut_request_core_robAddr,
  output [5:0]   responseOut_request_core_prfDest,
  output         responseOut_request_branch_valid,
  output [4:0]   responseOut_request_branch_mask,
  output         responseOut_request_writeData_valid,
  output [63:0]  responseOut_request_writeData_data,
  output [511:0] responseOut_request_cacheLine_cacheLine,
  output [1:0]   responseOut_request_cacheLine_response,
  output         writeBackIn_ready,
  input          writeBackIn_request_valid,
  input  [31:0]  writeBackIn_request_address,
  input  [511:0] writeBackIn_request_data,
  input          writeBackOut_ready,
  output         writeBackOut_request_valid,
  output [31:0]  writeBackOut_request_address,
  output [511:0] writeBackOut_request_data,
  input          branchOps_valid,
  input  [4:0]   branchOps_branchMask,
  input          branchOps_passed,
  output         fenceReady
);
  wire  requestWaitFIFO_clock; // @[replayUnit.scala 48:31]
  wire  requestWaitFIFO_reset; // @[replayUnit.scala 48:31]
  wire  requestWaitFIFO_write_ready; // @[replayUnit.scala 48:31]
  wire  requestWaitFIFO_write_data_valid; // @[replayUnit.scala 48:31]
  wire [31:0] requestWaitFIFO_write_data_address; // @[replayUnit.scala 48:31]
  wire [31:0] requestWaitFIFO_write_data_core_instruction; // @[replayUnit.scala 48:31]
  wire [3:0] requestWaitFIFO_write_data_core_robAddr; // @[replayUnit.scala 48:31]
  wire [5:0] requestWaitFIFO_write_data_core_prfDest; // @[replayUnit.scala 48:31]
  wire  requestWaitFIFO_write_data_branch_valid; // @[replayUnit.scala 48:31]
  wire [4:0] requestWaitFIFO_write_data_branch_mask; // @[replayUnit.scala 48:31]
  wire  requestWaitFIFO_write_data_writeData_valid; // @[replayUnit.scala 48:31]
  wire [63:0] requestWaitFIFO_write_data_writeData_data; // @[replayUnit.scala 48:31]
  wire [1:0] requestWaitFIFO_write_data_cacheLine_response; // @[replayUnit.scala 48:31]
  wire  requestWaitFIFO_read_ready; // @[replayUnit.scala 48:31]
  wire  requestWaitFIFO_read_data_valid; // @[replayUnit.scala 48:31]
  wire [31:0] requestWaitFIFO_read_data_address; // @[replayUnit.scala 48:31]
  wire [31:0] requestWaitFIFO_read_data_core_instruction; // @[replayUnit.scala 48:31]
  wire [3:0] requestWaitFIFO_read_data_core_robAddr; // @[replayUnit.scala 48:31]
  wire [5:0] requestWaitFIFO_read_data_core_prfDest; // @[replayUnit.scala 48:31]
  wire  requestWaitFIFO_read_data_branch_valid; // @[replayUnit.scala 48:31]
  wire [4:0] requestWaitFIFO_read_data_branch_mask; // @[replayUnit.scala 48:31]
  wire  requestWaitFIFO_read_data_writeData_valid; // @[replayUnit.scala 48:31]
  wire [63:0] requestWaitFIFO_read_data_writeData_data; // @[replayUnit.scala 48:31]
  wire [1:0] requestWaitFIFO_read_data_cacheLine_response; // @[replayUnit.scala 48:31]
  wire  requestWaitFIFO_isEmpty; // @[replayUnit.scala 48:31]
  wire  requestWaitFIFO_branchOps_valid; // @[replayUnit.scala 48:31]
  wire [4:0] requestWaitFIFO_branchOps_branchMask; // @[replayUnit.scala 48:31]
  wire  requestWaitFIFO_branchOps_passed; // @[replayUnit.scala 48:31]
  wire  writeBackFIFO_clock; // @[replayUnit.scala 56:29]
  wire  writeBackFIFO_reset; // @[replayUnit.scala 56:29]
  wire  writeBackFIFO_write_ready; // @[replayUnit.scala 56:29]
  wire  writeBackFIFO_write_data_valid; // @[replayUnit.scala 56:29]
  wire [31:0] writeBackFIFO_write_data_address; // @[replayUnit.scala 56:29]
  wire [511:0] writeBackFIFO_write_data_data; // @[replayUnit.scala 56:29]
  wire  writeBackFIFO_read_ready; // @[replayUnit.scala 56:29]
  wire  writeBackFIFO_read_data_valid; // @[replayUnit.scala 56:29]
  wire [31:0] writeBackFIFO_read_data_address; // @[replayUnit.scala 56:29]
  wire [511:0] writeBackFIFO_read_data_data; // @[replayUnit.scala 56:29]
  wire [4:0] _T_3 = requestIn_request_branch_mask & branchOps_branchMask; // @[utils.scala 62:31]
  wire  _T_4 = |_T_3; // @[utils.scala 62:55]
  wire [4:0] _requestWaitFIFO_write_data_branch_mask_T = requestIn_request_branch_mask ^ branchOps_branchMask; // @[utils.scala 63:42]
  wire [4:0] _GEN_2 = |_T_3 ? _requestWaitFIFO_write_data_branch_mask_T : requestIn_request_branch_mask; // @[utils.scala 62:60 63:23 65:23]
  wire  _GEN_3 = _T_4 ? 1'h0 : requestIn_request_branch_valid; // @[utils.scala 70:60 71:24 74:24]
  wire [4:0] _GEN_4 = _T_4 ? 5'h0 : requestIn_request_branch_mask; // @[utils.scala 70:60 72:23 75:23]
  wire [4:0] _GEN_5 = branchOps_passed ? _GEN_2 : _GEN_4; // @[utils.scala 60:30]
  wire  _GEN_6 = branchOps_passed ? requestIn_request_branch_valid : _GEN_3; // @[utils.scala 60:30 67:22]
  wire [4:0] _GEN_7 = branchOps_valid ? _GEN_5 : requestIn_request_branch_mask; // @[utils.scala 59:26 80:21]
  wire  _GEN_8 = branchOps_valid ? _GEN_6 : requestIn_request_branch_valid; // @[utils.scala 59:26 79:22]
  fifoWithBranchOps requestWaitFIFO ( // @[replayUnit.scala 48:31]
    .clock(requestWaitFIFO_clock),
    .reset(requestWaitFIFO_reset),
    .write_ready(requestWaitFIFO_write_ready),
    .write_data_valid(requestWaitFIFO_write_data_valid),
    .write_data_address(requestWaitFIFO_write_data_address),
    .write_data_core_instruction(requestWaitFIFO_write_data_core_instruction),
    .write_data_core_robAddr(requestWaitFIFO_write_data_core_robAddr),
    .write_data_core_prfDest(requestWaitFIFO_write_data_core_prfDest),
    .write_data_branch_valid(requestWaitFIFO_write_data_branch_valid),
    .write_data_branch_mask(requestWaitFIFO_write_data_branch_mask),
    .write_data_writeData_valid(requestWaitFIFO_write_data_writeData_valid),
    .write_data_writeData_data(requestWaitFIFO_write_data_writeData_data),
    .write_data_cacheLine_response(requestWaitFIFO_write_data_cacheLine_response),
    .read_ready(requestWaitFIFO_read_ready),
    .read_data_valid(requestWaitFIFO_read_data_valid),
    .read_data_address(requestWaitFIFO_read_data_address),
    .read_data_core_instruction(requestWaitFIFO_read_data_core_instruction),
    .read_data_core_robAddr(requestWaitFIFO_read_data_core_robAddr),
    .read_data_core_prfDest(requestWaitFIFO_read_data_core_prfDest),
    .read_data_branch_valid(requestWaitFIFO_read_data_branch_valid),
    .read_data_branch_mask(requestWaitFIFO_read_data_branch_mask),
    .read_data_writeData_valid(requestWaitFIFO_read_data_writeData_valid),
    .read_data_writeData_data(requestWaitFIFO_read_data_writeData_data),
    .read_data_cacheLine_response(requestWaitFIFO_read_data_cacheLine_response),
    .isEmpty(requestWaitFIFO_isEmpty),
    .branchOps_valid(requestWaitFIFO_branchOps_valid),
    .branchOps_branchMask(requestWaitFIFO_branchOps_branchMask),
    .branchOps_passed(requestWaitFIFO_branchOps_passed)
  );
  fifoBypassModule writeBackFIFO ( // @[replayUnit.scala 56:29]
    .clock(writeBackFIFO_clock),
    .reset(writeBackFIFO_reset),
    .write_ready(writeBackFIFO_write_ready),
    .write_data_valid(writeBackFIFO_write_data_valid),
    .write_data_address(writeBackFIFO_write_data_address),
    .write_data_data(writeBackFIFO_write_data_data),
    .read_ready(writeBackFIFO_read_ready),
    .read_data_valid(writeBackFIFO_read_data_valid),
    .read_data_address(writeBackFIFO_read_data_address),
    .read_data_data(writeBackFIFO_read_data_data)
  );
  assign requestIn_ready = requestWaitFIFO_write_ready; // @[replayUnit.scala 61:19 78:48 79:21]
  assign requestOut_request_valid = requestWaitFIFO_read_data_valid; // @[replayUnit.scala 86:22]
  assign requestOut_request_address = requestWaitFIFO_read_data_address; // @[replayUnit.scala 86:22]
  assign requestOut_request_core_instruction = requestWaitFIFO_read_data_core_instruction; // @[replayUnit.scala 86:22]
  assign requestOut_request_core_robAddr = requestWaitFIFO_read_data_core_robAddr; // @[replayUnit.scala 86:22]
  assign requestOut_request_core_prfDest = requestWaitFIFO_read_data_core_prfDest; // @[replayUnit.scala 86:22]
  assign requestOut_request_branch_valid = requestWaitFIFO_read_data_branch_valid; // @[replayUnit.scala 86:22]
  assign requestOut_request_branch_mask = requestWaitFIFO_read_data_branch_mask; // @[replayUnit.scala 86:22]
  assign requestOut_request_writeData_valid = requestWaitFIFO_read_data_writeData_valid; // @[replayUnit.scala 86:22]
  assign requestOut_request_writeData_data = requestWaitFIFO_read_data_writeData_data; // @[replayUnit.scala 86:22]
  assign requestOut_request_cacheLine_response = requestWaitFIFO_read_data_cacheLine_response; // @[replayUnit.scala 86:22]
  assign responseIn_ready = responseOut_ready; // @[replayUnit.scala 104:14]
  assign responseOut_request_valid = responseIn_request_valid; // @[replayUnit.scala 104:14]
  assign responseOut_request_address = responseIn_request_address; // @[replayUnit.scala 104:14]
  assign responseOut_request_core_instruction = responseIn_request_core_instruction; // @[replayUnit.scala 104:14]
  assign responseOut_request_core_robAddr = responseIn_request_core_robAddr; // @[replayUnit.scala 104:14]
  assign responseOut_request_core_prfDest = responseIn_request_core_prfDest; // @[replayUnit.scala 104:14]
  assign responseOut_request_branch_valid = responseIn_request_branch_valid; // @[replayUnit.scala 104:14]
  assign responseOut_request_branch_mask = responseIn_request_branch_mask; // @[replayUnit.scala 104:14]
  assign responseOut_request_writeData_valid = responseIn_request_writeData_valid; // @[replayUnit.scala 104:14]
  assign responseOut_request_writeData_data = responseIn_request_writeData_data; // @[replayUnit.scala 104:14]
  assign responseOut_request_cacheLine_cacheLine = responseIn_request_cacheLine_cacheLine; // @[replayUnit.scala 104:14]
  assign responseOut_request_cacheLine_response = responseIn_request_cacheLine_response; // @[replayUnit.scala 104:14]
  assign writeBackIn_ready = writeBackFIFO_write_ready; // @[replayUnit.scala 107:48 108:23 63:21]
  assign writeBackOut_request_valid = writeBackFIFO_read_data_valid; // @[replayUnit.scala 114:24]
  assign writeBackOut_request_address = writeBackFIFO_read_data_address; // @[replayUnit.scala 114:24]
  assign writeBackOut_request_data = writeBackFIFO_read_data_data; // @[replayUnit.scala 114:24]
  assign fenceReady = requestWaitFIFO_isEmpty; // @[replayUnit.scala 120:14]
  assign requestWaitFIFO_clock = clock;
  assign requestWaitFIFO_reset = reset;
  assign requestWaitFIFO_write_data_valid = requestIn_request_valid & requestIn_request_branch_valid &
    requestIn_request_valid; // @[replayUnit.scala 82:66 83:32 utils.scala 48:41]
  assign requestWaitFIFO_write_data_address = requestIn_request_valid & requestIn_request_branch_valid ?
    requestIn_request_address : 32'h0; // @[replayUnit.scala 82:66 83:32 utils.scala 49:41]
  assign requestWaitFIFO_write_data_core_instruction = requestIn_request_valid & requestIn_request_branch_valid ?
    requestIn_request_core_instruction : 32'h0; // @[replayUnit.scala 82:66 83:32 utils.scala 49:41]
  assign requestWaitFIFO_write_data_core_robAddr = requestIn_request_valid & requestIn_request_branch_valid ?
    requestIn_request_core_robAddr : 4'h0; // @[replayUnit.scala 82:66 83:32 utils.scala 49:41]
  assign requestWaitFIFO_write_data_core_prfDest = requestIn_request_valid & requestIn_request_branch_valid ?
    requestIn_request_core_prfDest : 6'h0; // @[replayUnit.scala 82:66 83:32 utils.scala 49:41]
  assign requestWaitFIFO_write_data_branch_valid = requestIn_request_valid & requestIn_request_branch_valid & _GEN_8; // @[replayUnit.scala 82:66 utils.scala 48:41]
  assign requestWaitFIFO_write_data_branch_mask = requestIn_request_valid & requestIn_request_branch_valid ? _GEN_7 : 5'h0
    ; // @[replayUnit.scala 82:66 utils.scala 49:41]
  assign requestWaitFIFO_write_data_writeData_valid = requestIn_request_valid & requestIn_request_branch_valid &
    requestIn_request_writeData_valid; // @[replayUnit.scala 82:66 83:32 utils.scala 48:41]
  assign requestWaitFIFO_write_data_writeData_data = requestIn_request_valid & requestIn_request_branch_valid ?
    requestIn_request_writeData_data : 64'h0; // @[replayUnit.scala 82:66 83:32 utils.scala 49:41]
  assign requestWaitFIFO_write_data_cacheLine_response = requestIn_request_valid & requestIn_request_branch_valid ?
    requestIn_request_cacheLine_response : 2'h0; // @[replayUnit.scala 82:66 83:32 utils.scala 49:41]
  assign requestWaitFIFO_read_ready = requestOut_ready; // @[replayUnit.scala 64:30 78:48 80:32]
  assign requestWaitFIFO_branchOps_valid = branchOps_valid; // @[replayUnit.scala 74:29]
  assign requestWaitFIFO_branchOps_branchMask = branchOps_branchMask; // @[replayUnit.scala 74:29]
  assign requestWaitFIFO_branchOps_passed = branchOps_passed; // @[replayUnit.scala 74:29]
  assign writeBackFIFO_clock = clock;
  assign writeBackFIFO_reset = reset;
  assign writeBackFIFO_write_data_valid = writeBackIn_request_valid; // @[replayUnit.scala 111:34 112:30 utils.scala 48:41]
  assign writeBackFIFO_write_data_address = writeBackIn_request_valid ? writeBackIn_request_address : 32'h0; // @[replayUnit.scala 111:34 112:30 utils.scala 49:41]
  assign writeBackFIFO_write_data_data = writeBackIn_request_valid ? writeBackIn_request_data : 512'h0; // @[replayUnit.scala 111:34 112:30 utils.scala 49:41]
  assign writeBackFIFO_read_ready = writeBackOut_ready; // @[replayUnit.scala 107:48 109:30 68:28]
endmodule
module fifoBaseModule(
  input         clock,
  input         reset,
  output        write_ready,
  input         write_data_valid,
  input  [31:0] write_data_address,
  input  [31:0] write_data_core_instruction,
  input  [3:0]  write_data_core_robAddr,
  input  [5:0]  write_data_core_prfDest,
  input         write_data_branch_valid,
  input  [4:0]  write_data_branch_mask,
  input  [63:0] write_data_writeData_data,
  input         read_ready,
  output        read_data_valid,
  output [31:0] read_data_address,
  output [31:0] read_data_core_instruction,
  output [3:0]  read_data_core_robAddr,
  output [5:0]  read_data_core_prfDest,
  output        read_data_branch_valid,
  output [4:0]  read_data_branch_mask,
  output [63:0] read_data_writeData_data,
  output        isEmpty
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] memReg_0_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_0_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_0_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_0_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_0_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_0_branch_mask; // @[fifo.scala 27:33]
  reg [63:0] memReg_0_writeData_data; // @[fifo.scala 27:33]
  reg [31:0] memReg_1_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_1_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_1_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_1_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_1_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_1_branch_mask; // @[fifo.scala 27:33]
  reg [63:0] memReg_1_writeData_data; // @[fifo.scala 27:33]
  reg [31:0] memReg_2_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_2_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_2_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_2_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_2_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_2_branch_mask; // @[fifo.scala 27:33]
  reg [63:0] memReg_2_writeData_data; // @[fifo.scala 27:33]
  reg [31:0] memReg_3_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_3_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_3_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_3_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_3_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_3_branch_mask; // @[fifo.scala 27:33]
  reg [63:0] memReg_3_writeData_data; // @[fifo.scala 27:33]
  reg [31:0] memReg_4_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_4_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_4_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_4_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_4_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_4_branch_mask; // @[fifo.scala 27:33]
  reg [63:0] memReg_4_writeData_data; // @[fifo.scala 27:33]
  reg [31:0] memReg_5_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_5_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_5_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_5_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_5_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_5_branch_mask; // @[fifo.scala 27:33]
  reg [63:0] memReg_5_writeData_data; // @[fifo.scala 27:33]
  reg [31:0] memReg_6_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_6_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_6_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_6_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_6_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_6_branch_mask; // @[fifo.scala 27:33]
  reg [63:0] memReg_6_writeData_data; // @[fifo.scala 27:33]
  reg [31:0] memReg_7_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_7_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_7_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_7_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_7_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_7_branch_mask; // @[fifo.scala 27:33]
  reg [63:0] memReg_7_writeData_data; // @[fifo.scala 27:33]
  reg [31:0] memReg_8_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_8_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_8_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_8_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_8_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_8_branch_mask; // @[fifo.scala 27:33]
  reg [63:0] memReg_8_writeData_data; // @[fifo.scala 27:33]
  reg [31:0] memReg_9_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_9_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_9_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_9_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_9_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_9_branch_mask; // @[fifo.scala 27:33]
  reg [63:0] memReg_9_writeData_data; // @[fifo.scala 27:33]
  reg [31:0] memReg_10_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_10_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_10_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_10_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_10_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_10_branch_mask; // @[fifo.scala 27:33]
  reg [63:0] memReg_10_writeData_data; // @[fifo.scala 27:33]
  reg [31:0] memReg_11_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_11_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_11_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_11_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_11_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_11_branch_mask; // @[fifo.scala 27:33]
  reg [63:0] memReg_11_writeData_data; // @[fifo.scala 27:33]
  reg [31:0] memReg_12_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_12_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_12_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_12_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_12_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_12_branch_mask; // @[fifo.scala 27:33]
  reg [63:0] memReg_12_writeData_data; // @[fifo.scala 27:33]
  reg [31:0] memReg_13_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_13_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_13_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_13_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_13_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_13_branch_mask; // @[fifo.scala 27:33]
  reg [63:0] memReg_13_writeData_data; // @[fifo.scala 27:33]
  reg [31:0] memReg_14_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_14_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_14_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_14_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_14_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_14_branch_mask; // @[fifo.scala 27:33]
  reg [63:0] memReg_14_writeData_data; // @[fifo.scala 27:33]
  reg [31:0] memReg_15_address; // @[fifo.scala 27:33]
  reg [31:0] memReg_15_core_instruction; // @[fifo.scala 27:33]
  reg [3:0] memReg_15_core_robAddr; // @[fifo.scala 27:33]
  reg [5:0] memReg_15_core_prfDest; // @[fifo.scala 27:33]
  reg  memReg_15_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_15_branch_mask; // @[fifo.scala 27:33]
  reg [63:0] memReg_15_writeData_data; // @[fifo.scala 27:33]
  reg [3:0] readPtr; // @[fifo.scala 33:25]
  wire [3:0] _nextVal_T_2 = readPtr + 4'h1; // @[fifo.scala 34:60]
  wire [3:0] nextRead = readPtr == 4'hf ? 4'h0 : _nextVal_T_2; // @[fifo.scala 34:22]
  wire [1:0] op = {write_data_valid,read_ready}; // @[fifo.scala 46:29]
  reg  emptyReg; // @[fifo.scala 43:25]
  wire  _T_2 = ~emptyReg; // @[fifo.scala 52:12]
  wire  _GEN_21 = 2'h2 == op ? 1'h0 : 2'h3 == op & _T_2; // @[fifo.scala 49:14]
  wire  _GEN_24 = 2'h1 == op ? _T_2 : _GEN_21; // @[fifo.scala 49:14]
  wire  incrRead = 2'h0 == op ? 1'h0 : _GEN_24; // @[fifo.scala 49:14]
  reg [3:0] writePtr; // @[fifo.scala 33:25]
  wire [3:0] _nextVal_T_5 = writePtr + 4'h1; // @[fifo.scala 34:60]
  wire [3:0] nextWrite = writePtr == 4'hf ? 4'h0 : _nextVal_T_5; // @[fifo.scala 34:22]
  reg  fullReg; // @[fifo.scala 44:34]
  wire  _T_4 = ~fullReg; // @[fifo.scala 59:12]
  wire  _GEN_18 = 2'h2 == op ? _T_4 : 2'h3 == op & _T_4; // @[fifo.scala 49:14]
  wire  _GEN_25 = 2'h1 == op ? 1'h0 : _GEN_18; // @[fifo.scala 49:14]
  wire  incrWrite = 2'h0 == op ? 1'h0 : _GEN_25; // @[fifo.scala 49:14]
  wire  _GEN_3 = ~emptyReg ? nextRead == writePtr : emptyReg; // @[fifo.scala 52:23 54:18 43:25]
  wire  _GEN_6 = ~fullReg ? 1'h0 : emptyReg; // @[fifo.scala 59:22 61:18 43:25]
  wire  _GEN_7 = ~fullReg ? nextWrite == readPtr : fullReg; // @[fifo.scala 59:22 62:17 44:34]
  wire  _fullReg_T_2 = emptyReg ? 1'h0 : nextWrite == nextRead; // @[fifo.scala 70:23]
  wire  _GEN_10 = _T_4 ? _fullReg_T_2 : fullReg; // @[fifo.scala 67:22 70:17 44:34]
  wire  _emptyReg_T_2 = fullReg ? 1'h0 : nextRead == nextWrite; // @[fifo.scala 75:24]
  wire  _GEN_11 = _T_2 ? 1'h0 : _GEN_10; // @[fifo.scala 73:23 74:17]
  wire  _GEN_12 = _T_2 ? _emptyReg_T_2 : _GEN_6; // @[fifo.scala 73:23 75:18]
  wire  _GEN_15 = 2'h3 == op ? _GEN_12 : emptyReg; // @[fifo.scala 49:14 43:25]
  wire  _GEN_16 = 2'h3 == op ? _GEN_11 : fullReg; // @[fifo.scala 49:14 44:34]
  wire  _GEN_19 = 2'h2 == op ? _GEN_6 : _GEN_15; // @[fifo.scala 49:14]
  wire  _GEN_23 = 2'h1 == op ? _GEN_3 : _GEN_19; // @[fifo.scala 49:14]
  wire  _GEN_27 = 2'h0 == op ? emptyReg : _GEN_23; // @[fifo.scala 49:14 43:25]
  wire [31:0] _GEN_431 = 4'h1 == readPtr ? memReg_1_address : memReg_0_address; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_432 = 4'h2 == readPtr ? memReg_2_address : _GEN_431; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_433 = 4'h3 == readPtr ? memReg_3_address : _GEN_432; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_434 = 4'h4 == readPtr ? memReg_4_address : _GEN_433; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_435 = 4'h5 == readPtr ? memReg_5_address : _GEN_434; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_436 = 4'h6 == readPtr ? memReg_6_address : _GEN_435; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_437 = 4'h7 == readPtr ? memReg_7_address : _GEN_436; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_438 = 4'h8 == readPtr ? memReg_8_address : _GEN_437; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_439 = 4'h9 == readPtr ? memReg_9_address : _GEN_438; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_440 = 4'ha == readPtr ? memReg_10_address : _GEN_439; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_441 = 4'hb == readPtr ? memReg_11_address : _GEN_440; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_442 = 4'hc == readPtr ? memReg_12_address : _GEN_441; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_443 = 4'hd == readPtr ? memReg_13_address : _GEN_442; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_444 = 4'he == readPtr ? memReg_14_address : _GEN_443; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_447 = 4'h1 == readPtr ? memReg_1_core_instruction : memReg_0_core_instruction; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_448 = 4'h2 == readPtr ? memReg_2_core_instruction : _GEN_447; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_449 = 4'h3 == readPtr ? memReg_3_core_instruction : _GEN_448; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_450 = 4'h4 == readPtr ? memReg_4_core_instruction : _GEN_449; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_451 = 4'h5 == readPtr ? memReg_5_core_instruction : _GEN_450; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_452 = 4'h6 == readPtr ? memReg_6_core_instruction : _GEN_451; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_453 = 4'h7 == readPtr ? memReg_7_core_instruction : _GEN_452; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_454 = 4'h8 == readPtr ? memReg_8_core_instruction : _GEN_453; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_455 = 4'h9 == readPtr ? memReg_9_core_instruction : _GEN_454; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_456 = 4'ha == readPtr ? memReg_10_core_instruction : _GEN_455; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_457 = 4'hb == readPtr ? memReg_11_core_instruction : _GEN_456; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_458 = 4'hc == readPtr ? memReg_12_core_instruction : _GEN_457; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_459 = 4'hd == readPtr ? memReg_13_core_instruction : _GEN_458; // @[fifo.scala 86:{13,13}]
  wire [31:0] _GEN_460 = 4'he == readPtr ? memReg_14_core_instruction : _GEN_459; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_463 = 4'h1 == readPtr ? memReg_1_core_robAddr : memReg_0_core_robAddr; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_464 = 4'h2 == readPtr ? memReg_2_core_robAddr : _GEN_463; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_465 = 4'h3 == readPtr ? memReg_3_core_robAddr : _GEN_464; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_466 = 4'h4 == readPtr ? memReg_4_core_robAddr : _GEN_465; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_467 = 4'h5 == readPtr ? memReg_5_core_robAddr : _GEN_466; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_468 = 4'h6 == readPtr ? memReg_6_core_robAddr : _GEN_467; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_469 = 4'h7 == readPtr ? memReg_7_core_robAddr : _GEN_468; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_470 = 4'h8 == readPtr ? memReg_8_core_robAddr : _GEN_469; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_471 = 4'h9 == readPtr ? memReg_9_core_robAddr : _GEN_470; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_472 = 4'ha == readPtr ? memReg_10_core_robAddr : _GEN_471; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_473 = 4'hb == readPtr ? memReg_11_core_robAddr : _GEN_472; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_474 = 4'hc == readPtr ? memReg_12_core_robAddr : _GEN_473; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_475 = 4'hd == readPtr ? memReg_13_core_robAddr : _GEN_474; // @[fifo.scala 86:{13,13}]
  wire [3:0] _GEN_476 = 4'he == readPtr ? memReg_14_core_robAddr : _GEN_475; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_479 = 4'h1 == readPtr ? memReg_1_core_prfDest : memReg_0_core_prfDest; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_480 = 4'h2 == readPtr ? memReg_2_core_prfDest : _GEN_479; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_481 = 4'h3 == readPtr ? memReg_3_core_prfDest : _GEN_480; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_482 = 4'h4 == readPtr ? memReg_4_core_prfDest : _GEN_481; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_483 = 4'h5 == readPtr ? memReg_5_core_prfDest : _GEN_482; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_484 = 4'h6 == readPtr ? memReg_6_core_prfDest : _GEN_483; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_485 = 4'h7 == readPtr ? memReg_7_core_prfDest : _GEN_484; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_486 = 4'h8 == readPtr ? memReg_8_core_prfDest : _GEN_485; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_487 = 4'h9 == readPtr ? memReg_9_core_prfDest : _GEN_486; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_488 = 4'ha == readPtr ? memReg_10_core_prfDest : _GEN_487; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_489 = 4'hb == readPtr ? memReg_11_core_prfDest : _GEN_488; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_490 = 4'hc == readPtr ? memReg_12_core_prfDest : _GEN_489; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_491 = 4'hd == readPtr ? memReg_13_core_prfDest : _GEN_490; // @[fifo.scala 86:{13,13}]
  wire [5:0] _GEN_492 = 4'he == readPtr ? memReg_14_core_prfDest : _GEN_491; // @[fifo.scala 86:{13,13}]
  wire  _GEN_495 = 4'h1 == readPtr ? memReg_1_branch_valid : memReg_0_branch_valid; // @[fifo.scala 86:{13,13}]
  wire  _GEN_496 = 4'h2 == readPtr ? memReg_2_branch_valid : _GEN_495; // @[fifo.scala 86:{13,13}]
  wire  _GEN_497 = 4'h3 == readPtr ? memReg_3_branch_valid : _GEN_496; // @[fifo.scala 86:{13,13}]
  wire  _GEN_498 = 4'h4 == readPtr ? memReg_4_branch_valid : _GEN_497; // @[fifo.scala 86:{13,13}]
  wire  _GEN_499 = 4'h5 == readPtr ? memReg_5_branch_valid : _GEN_498; // @[fifo.scala 86:{13,13}]
  wire  _GEN_500 = 4'h6 == readPtr ? memReg_6_branch_valid : _GEN_499; // @[fifo.scala 86:{13,13}]
  wire  _GEN_501 = 4'h7 == readPtr ? memReg_7_branch_valid : _GEN_500; // @[fifo.scala 86:{13,13}]
  wire  _GEN_502 = 4'h8 == readPtr ? memReg_8_branch_valid : _GEN_501; // @[fifo.scala 86:{13,13}]
  wire  _GEN_503 = 4'h9 == readPtr ? memReg_9_branch_valid : _GEN_502; // @[fifo.scala 86:{13,13}]
  wire  _GEN_504 = 4'ha == readPtr ? memReg_10_branch_valid : _GEN_503; // @[fifo.scala 86:{13,13}]
  wire  _GEN_505 = 4'hb == readPtr ? memReg_11_branch_valid : _GEN_504; // @[fifo.scala 86:{13,13}]
  wire  _GEN_506 = 4'hc == readPtr ? memReg_12_branch_valid : _GEN_505; // @[fifo.scala 86:{13,13}]
  wire  _GEN_507 = 4'hd == readPtr ? memReg_13_branch_valid : _GEN_506; // @[fifo.scala 86:{13,13}]
  wire  _GEN_508 = 4'he == readPtr ? memReg_14_branch_valid : _GEN_507; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_511 = 4'h1 == readPtr ? memReg_1_branch_mask : memReg_0_branch_mask; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_512 = 4'h2 == readPtr ? memReg_2_branch_mask : _GEN_511; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_513 = 4'h3 == readPtr ? memReg_3_branch_mask : _GEN_512; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_514 = 4'h4 == readPtr ? memReg_4_branch_mask : _GEN_513; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_515 = 4'h5 == readPtr ? memReg_5_branch_mask : _GEN_514; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_516 = 4'h6 == readPtr ? memReg_6_branch_mask : _GEN_515; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_517 = 4'h7 == readPtr ? memReg_7_branch_mask : _GEN_516; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_518 = 4'h8 == readPtr ? memReg_8_branch_mask : _GEN_517; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_519 = 4'h9 == readPtr ? memReg_9_branch_mask : _GEN_518; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_520 = 4'ha == readPtr ? memReg_10_branch_mask : _GEN_519; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_521 = 4'hb == readPtr ? memReg_11_branch_mask : _GEN_520; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_522 = 4'hc == readPtr ? memReg_12_branch_mask : _GEN_521; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_523 = 4'hd == readPtr ? memReg_13_branch_mask : _GEN_522; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_524 = 4'he == readPtr ? memReg_14_branch_mask : _GEN_523; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_543 = 4'h1 == readPtr ? memReg_1_writeData_data : memReg_0_writeData_data; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_544 = 4'h2 == readPtr ? memReg_2_writeData_data : _GEN_543; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_545 = 4'h3 == readPtr ? memReg_3_writeData_data : _GEN_544; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_546 = 4'h4 == readPtr ? memReg_4_writeData_data : _GEN_545; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_547 = 4'h5 == readPtr ? memReg_5_writeData_data : _GEN_546; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_548 = 4'h6 == readPtr ? memReg_6_writeData_data : _GEN_547; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_549 = 4'h7 == readPtr ? memReg_7_writeData_data : _GEN_548; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_550 = 4'h8 == readPtr ? memReg_8_writeData_data : _GEN_549; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_551 = 4'h9 == readPtr ? memReg_9_writeData_data : _GEN_550; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_552 = 4'ha == readPtr ? memReg_10_writeData_data : _GEN_551; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_553 = 4'hb == readPtr ? memReg_11_writeData_data : _GEN_552; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_554 = 4'hc == readPtr ? memReg_12_writeData_data : _GEN_553; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_555 = 4'hd == readPtr ? memReg_13_writeData_data : _GEN_554; // @[fifo.scala 86:{13,13}]
  wire [63:0] _GEN_556 = 4'he == readPtr ? memReg_14_writeData_data : _GEN_555; // @[fifo.scala 86:{13,13}]
  assign write_ready = ~fullReg; // @[fifo.scala 88:18]
  assign read_data_valid = ~emptyReg; // @[fifo.scala 87:22]
  assign read_data_address = 4'hf == readPtr ? memReg_15_address : _GEN_444; // @[fifo.scala 86:{13,13}]
  assign read_data_core_instruction = 4'hf == readPtr ? memReg_15_core_instruction : _GEN_460; // @[fifo.scala 86:{13,13}]
  assign read_data_core_robAddr = 4'hf == readPtr ? memReg_15_core_robAddr : _GEN_476; // @[fifo.scala 86:{13,13}]
  assign read_data_core_prfDest = 4'hf == readPtr ? memReg_15_core_prfDest : _GEN_492; // @[fifo.scala 86:{13,13}]
  assign read_data_branch_valid = 4'hf == readPtr ? memReg_15_branch_valid : _GEN_508; // @[fifo.scala 86:{13,13}]
  assign read_data_branch_mask = 4'hf == readPtr ? memReg_15_branch_mask : _GEN_524; // @[fifo.scala 86:{13,13}]
  assign read_data_writeData_data = 4'hf == readPtr ? memReg_15_writeData_data : _GEN_556; // @[fifo.scala 86:{13,13}]
  assign isEmpty = emptyReg; // @[fifo.scala 89:11]
  always @(posedge clock) begin
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_branch_valid <= write_data_branch_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_branch_mask <= write_data_branch_mask; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_branch_valid <= write_data_branch_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_branch_mask <= write_data_branch_mask; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_branch_valid <= write_data_branch_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_branch_mask <= write_data_branch_mask; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_branch_valid <= write_data_branch_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_branch_mask <= write_data_branch_mask; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_branch_valid <= write_data_branch_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_branch_mask <= write_data_branch_mask; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_branch_valid <= write_data_branch_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_branch_mask <= write_data_branch_mask; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_branch_valid <= write_data_branch_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_branch_mask <= write_data_branch_mask; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_branch_valid <= write_data_branch_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_branch_mask <= write_data_branch_mask; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_branch_valid <= write_data_branch_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_branch_mask <= write_data_branch_mask; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_branch_valid <= write_data_branch_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_branch_mask <= write_data_branch_mask; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_branch_valid <= write_data_branch_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_branch_mask <= write_data_branch_mask; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_branch_valid <= write_data_branch_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_branch_mask <= write_data_branch_mask; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_branch_valid <= write_data_branch_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_branch_mask <= write_data_branch_mask; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_branch_valid <= write_data_branch_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_branch_mask <= write_data_branch_mask; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_branch_valid <= write_data_branch_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_branch_mask <= write_data_branch_mask; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_core_instruction <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_core_instruction <= write_data_core_instruction; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_core_robAddr <= 4'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_core_robAddr <= write_data_core_robAddr; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_core_prfDest <= 6'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_core_prfDest <= write_data_core_prfDest; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_branch_valid <= write_data_branch_valid; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_branch_mask <= write_data_branch_mask; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_writeData_data <= 64'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (4'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_writeData_data <= write_data_writeData_data; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 33:25]
      readPtr <= 4'h0; // @[fifo.scala 33:25]
    end else if (incrRead) begin // @[fifo.scala 35:15]
      if (readPtr == 4'hf) begin // @[fifo.scala 34:22]
        readPtr <= 4'h0;
      end else begin
        readPtr <= _nextVal_T_2;
      end
    end
    emptyReg <= reset | _GEN_27; // @[fifo.scala 43:{25,25}]
    if (reset) begin // @[fifo.scala 33:25]
      writePtr <= 4'h0; // @[fifo.scala 33:25]
    end else if (incrWrite) begin // @[fifo.scala 35:15]
      if (writePtr == 4'hf) begin // @[fifo.scala 34:22]
        writePtr <= 4'h0;
      end else begin
        writePtr <= _nextVal_T_5;
      end
    end
    if (reset) begin // @[fifo.scala 44:34]
      fullReg <= 1'h0; // @[fifo.scala 44:34]
    end else if (!(2'h0 == op)) begin // @[fifo.scala 49:14]
      if (2'h1 == op) begin // @[fifo.scala 49:14]
        if (~emptyReg) begin // @[fifo.scala 52:23]
          fullReg <= 1'h0; // @[fifo.scala 53:17]
        end
      end else if (2'h2 == op) begin // @[fifo.scala 49:14]
        fullReg <= _GEN_7;
      end else begin
        fullReg <= _GEN_16;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  memReg_0_address = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  memReg_0_core_instruction = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  memReg_0_core_robAddr = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  memReg_0_core_prfDest = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  memReg_0_branch_valid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  memReg_0_branch_mask = _RAND_5[4:0];
  _RAND_6 = {2{`RANDOM}};
  memReg_0_writeData_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  memReg_1_address = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  memReg_1_core_instruction = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  memReg_1_core_robAddr = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  memReg_1_core_prfDest = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  memReg_1_branch_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  memReg_1_branch_mask = _RAND_12[4:0];
  _RAND_13 = {2{`RANDOM}};
  memReg_1_writeData_data = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  memReg_2_address = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  memReg_2_core_instruction = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  memReg_2_core_robAddr = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  memReg_2_core_prfDest = _RAND_17[5:0];
  _RAND_18 = {1{`RANDOM}};
  memReg_2_branch_valid = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  memReg_2_branch_mask = _RAND_19[4:0];
  _RAND_20 = {2{`RANDOM}};
  memReg_2_writeData_data = _RAND_20[63:0];
  _RAND_21 = {1{`RANDOM}};
  memReg_3_address = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  memReg_3_core_instruction = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  memReg_3_core_robAddr = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  memReg_3_core_prfDest = _RAND_24[5:0];
  _RAND_25 = {1{`RANDOM}};
  memReg_3_branch_valid = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  memReg_3_branch_mask = _RAND_26[4:0];
  _RAND_27 = {2{`RANDOM}};
  memReg_3_writeData_data = _RAND_27[63:0];
  _RAND_28 = {1{`RANDOM}};
  memReg_4_address = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  memReg_4_core_instruction = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  memReg_4_core_robAddr = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  memReg_4_core_prfDest = _RAND_31[5:0];
  _RAND_32 = {1{`RANDOM}};
  memReg_4_branch_valid = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  memReg_4_branch_mask = _RAND_33[4:0];
  _RAND_34 = {2{`RANDOM}};
  memReg_4_writeData_data = _RAND_34[63:0];
  _RAND_35 = {1{`RANDOM}};
  memReg_5_address = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  memReg_5_core_instruction = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  memReg_5_core_robAddr = _RAND_37[3:0];
  _RAND_38 = {1{`RANDOM}};
  memReg_5_core_prfDest = _RAND_38[5:0];
  _RAND_39 = {1{`RANDOM}};
  memReg_5_branch_valid = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  memReg_5_branch_mask = _RAND_40[4:0];
  _RAND_41 = {2{`RANDOM}};
  memReg_5_writeData_data = _RAND_41[63:0];
  _RAND_42 = {1{`RANDOM}};
  memReg_6_address = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  memReg_6_core_instruction = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  memReg_6_core_robAddr = _RAND_44[3:0];
  _RAND_45 = {1{`RANDOM}};
  memReg_6_core_prfDest = _RAND_45[5:0];
  _RAND_46 = {1{`RANDOM}};
  memReg_6_branch_valid = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  memReg_6_branch_mask = _RAND_47[4:0];
  _RAND_48 = {2{`RANDOM}};
  memReg_6_writeData_data = _RAND_48[63:0];
  _RAND_49 = {1{`RANDOM}};
  memReg_7_address = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  memReg_7_core_instruction = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  memReg_7_core_robAddr = _RAND_51[3:0];
  _RAND_52 = {1{`RANDOM}};
  memReg_7_core_prfDest = _RAND_52[5:0];
  _RAND_53 = {1{`RANDOM}};
  memReg_7_branch_valid = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  memReg_7_branch_mask = _RAND_54[4:0];
  _RAND_55 = {2{`RANDOM}};
  memReg_7_writeData_data = _RAND_55[63:0];
  _RAND_56 = {1{`RANDOM}};
  memReg_8_address = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  memReg_8_core_instruction = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  memReg_8_core_robAddr = _RAND_58[3:0];
  _RAND_59 = {1{`RANDOM}};
  memReg_8_core_prfDest = _RAND_59[5:0];
  _RAND_60 = {1{`RANDOM}};
  memReg_8_branch_valid = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  memReg_8_branch_mask = _RAND_61[4:0];
  _RAND_62 = {2{`RANDOM}};
  memReg_8_writeData_data = _RAND_62[63:0];
  _RAND_63 = {1{`RANDOM}};
  memReg_9_address = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  memReg_9_core_instruction = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  memReg_9_core_robAddr = _RAND_65[3:0];
  _RAND_66 = {1{`RANDOM}};
  memReg_9_core_prfDest = _RAND_66[5:0];
  _RAND_67 = {1{`RANDOM}};
  memReg_9_branch_valid = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  memReg_9_branch_mask = _RAND_68[4:0];
  _RAND_69 = {2{`RANDOM}};
  memReg_9_writeData_data = _RAND_69[63:0];
  _RAND_70 = {1{`RANDOM}};
  memReg_10_address = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  memReg_10_core_instruction = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  memReg_10_core_robAddr = _RAND_72[3:0];
  _RAND_73 = {1{`RANDOM}};
  memReg_10_core_prfDest = _RAND_73[5:0];
  _RAND_74 = {1{`RANDOM}};
  memReg_10_branch_valid = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  memReg_10_branch_mask = _RAND_75[4:0];
  _RAND_76 = {2{`RANDOM}};
  memReg_10_writeData_data = _RAND_76[63:0];
  _RAND_77 = {1{`RANDOM}};
  memReg_11_address = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  memReg_11_core_instruction = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  memReg_11_core_robAddr = _RAND_79[3:0];
  _RAND_80 = {1{`RANDOM}};
  memReg_11_core_prfDest = _RAND_80[5:0];
  _RAND_81 = {1{`RANDOM}};
  memReg_11_branch_valid = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  memReg_11_branch_mask = _RAND_82[4:0];
  _RAND_83 = {2{`RANDOM}};
  memReg_11_writeData_data = _RAND_83[63:0];
  _RAND_84 = {1{`RANDOM}};
  memReg_12_address = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  memReg_12_core_instruction = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  memReg_12_core_robAddr = _RAND_86[3:0];
  _RAND_87 = {1{`RANDOM}};
  memReg_12_core_prfDest = _RAND_87[5:0];
  _RAND_88 = {1{`RANDOM}};
  memReg_12_branch_valid = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  memReg_12_branch_mask = _RAND_89[4:0];
  _RAND_90 = {2{`RANDOM}};
  memReg_12_writeData_data = _RAND_90[63:0];
  _RAND_91 = {1{`RANDOM}};
  memReg_13_address = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  memReg_13_core_instruction = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  memReg_13_core_robAddr = _RAND_93[3:0];
  _RAND_94 = {1{`RANDOM}};
  memReg_13_core_prfDest = _RAND_94[5:0];
  _RAND_95 = {1{`RANDOM}};
  memReg_13_branch_valid = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  memReg_13_branch_mask = _RAND_96[4:0];
  _RAND_97 = {2{`RANDOM}};
  memReg_13_writeData_data = _RAND_97[63:0];
  _RAND_98 = {1{`RANDOM}};
  memReg_14_address = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  memReg_14_core_instruction = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  memReg_14_core_robAddr = _RAND_100[3:0];
  _RAND_101 = {1{`RANDOM}};
  memReg_14_core_prfDest = _RAND_101[5:0];
  _RAND_102 = {1{`RANDOM}};
  memReg_14_branch_valid = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  memReg_14_branch_mask = _RAND_103[4:0];
  _RAND_104 = {2{`RANDOM}};
  memReg_14_writeData_data = _RAND_104[63:0];
  _RAND_105 = {1{`RANDOM}};
  memReg_15_address = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  memReg_15_core_instruction = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  memReg_15_core_robAddr = _RAND_107[3:0];
  _RAND_108 = {1{`RANDOM}};
  memReg_15_core_prfDest = _RAND_108[5:0];
  _RAND_109 = {1{`RANDOM}};
  memReg_15_branch_valid = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  memReg_15_branch_mask = _RAND_110[4:0];
  _RAND_111 = {2{`RANDOM}};
  memReg_15_writeData_data = _RAND_111[63:0];
  _RAND_112 = {1{`RANDOM}};
  readPtr = _RAND_112[3:0];
  _RAND_113 = {1{`RANDOM}};
  emptyReg = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  writePtr = _RAND_114[3:0];
  _RAND_115 = {1{`RANDOM}};
  fullReg = _RAND_115[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module moduleCounter(
  input   clock,
  input   reset,
  output  count,
  input   incrm
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  cntReg; // @[utils.scala 17:23]
  assign count = cntReg; // @[utils.scala 20:9]
  always @(posedge clock) begin
    if (reset) begin // @[utils.scala 17:23]
      cntReg <= 1'h0; // @[utils.scala 17:23]
    end else if (incrm & cntReg) begin // @[utils.scala 18:16]
      cntReg <= 1'h0;
    end else if (incrm) begin // @[utils.scala 19:20]
      cntReg <= cntReg + 1'h1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cntReg = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module peripheralUnit(
  input         clock,
  input         reset,
  output        request_ready,
  input         request_request_valid,
  input  [31:0] request_request_address,
  input  [31:0] request_request_core_instruction,
  input  [3:0]  request_request_core_robAddr,
  input  [5:0]  request_request_core_prfDest,
  input         request_request_branch_valid,
  input  [4:0]  request_request_branch_mask,
  input         request_request_writeData_valid,
  input  [63:0] request_request_writeData_data,
  input         responseOut_ready,
  output        responseOut_request_valid,
  output [31:0] responseOut_request_address,
  output [31:0] responseOut_request_core_instruction,
  output [3:0]  responseOut_request_core_robAddr,
  output [5:0]  responseOut_request_core_prfDest,
  output        responseOut_request_branch_valid,
  output [4:0]  responseOut_request_branch_mask,
  output [63:0] responseOut_request_writeData_data,
  output [31:0] bus_AWADDR,
  output [7:0]  bus_AWLEN,
  output [2:0]  bus_AWSIZE,
  output [1:0]  bus_AWBURST,
  output [2:0]  bus_AWPROT,
  output        bus_AWVALID,
  input         bus_AWREADY,
  output [31:0] bus_WDATA,
  output [3:0]  bus_WSTRB,
  output        bus_WLAST,
  output        bus_WVALID,
  input         bus_WREADY,
  input  [1:0]  bus_BID,
  input  [1:0]  bus_BRESP,
  input         bus_BVALID,
  output        bus_BREADY,
  output [31:0] bus_ARADDR,
  output [7:0]  bus_ARLEN,
  output [2:0]  bus_ARSIZE,
  output [1:0]  bus_ARBURST,
  output [2:0]  bus_ARPROT,
  output        bus_ARVALID,
  input         bus_ARREADY,
  input  [1:0]  bus_RID,
  input  [31:0] bus_RDATA,
  input  [1:0]  bus_RRESP,
  input         bus_RLAST,
  input         bus_RVALID,
  output        bus_RREADY,
  output        writeInstructionCommit_ready,
  input         writeInstructionCommit_fired,
  input         branchOps_valid,
  input  [4:0]  branchOps_branchMask,
  input         branchOps_passed
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
`endif // RANDOMIZE_REG_INIT
  wire  peripheralMSHR_clock; // @[peripheralUnit.scala 82:30]
  wire  peripheralMSHR_reset; // @[peripheralUnit.scala 82:30]
  wire  peripheralMSHR_write_ready; // @[peripheralUnit.scala 82:30]
  wire  peripheralMSHR_write_data_valid; // @[peripheralUnit.scala 82:30]
  wire [31:0] peripheralMSHR_write_data_address; // @[peripheralUnit.scala 82:30]
  wire [31:0] peripheralMSHR_write_data_core_instruction; // @[peripheralUnit.scala 82:30]
  wire [3:0] peripheralMSHR_write_data_core_robAddr; // @[peripheralUnit.scala 82:30]
  wire [5:0] peripheralMSHR_write_data_core_prfDest; // @[peripheralUnit.scala 82:30]
  wire  peripheralMSHR_write_data_branch_valid; // @[peripheralUnit.scala 82:30]
  wire [4:0] peripheralMSHR_write_data_branch_mask; // @[peripheralUnit.scala 82:30]
  wire [63:0] peripheralMSHR_write_data_writeData_data; // @[peripheralUnit.scala 82:30]
  wire  peripheralMSHR_read_ready; // @[peripheralUnit.scala 82:30]
  wire  peripheralMSHR_read_data_valid; // @[peripheralUnit.scala 82:30]
  wire [31:0] peripheralMSHR_read_data_address; // @[peripheralUnit.scala 82:30]
  wire [31:0] peripheralMSHR_read_data_core_instruction; // @[peripheralUnit.scala 82:30]
  wire [3:0] peripheralMSHR_read_data_core_robAddr; // @[peripheralUnit.scala 82:30]
  wire [5:0] peripheralMSHR_read_data_core_prfDest; // @[peripheralUnit.scala 82:30]
  wire  peripheralMSHR_read_data_branch_valid; // @[peripheralUnit.scala 82:30]
  wire [4:0] peripheralMSHR_read_data_branch_mask; // @[peripheralUnit.scala 82:30]
  wire [63:0] peripheralMSHR_read_data_writeData_data; // @[peripheralUnit.scala 82:30]
  wire  peripheralMSHR_isEmpty; // @[peripheralUnit.scala 82:30]
  wire  writeCounter_clock; // @[peripheralUnit.scala 114:28]
  wire  writeCounter_reset; // @[peripheralUnit.scala 114:28]
  wire  writeCounter_count; // @[peripheralUnit.scala 114:28]
  wire  writeCounter_incrm; // @[peripheralUnit.scala 114:28]
  wire  readCounter_clock; // @[peripheralUnit.scala 197:27]
  wire  readCounter_reset; // @[peripheralUnit.scala 197:27]
  wire  readCounter_count; // @[peripheralUnit.scala 197:27]
  wire  readCounter_incrm; // @[peripheralUnit.scala 197:27]
  reg  requestBuffer_valid; // @[peripheralUnit.scala 69:30]
  reg [31:0] requestBuffer_address; // @[peripheralUnit.scala 69:30]
  reg [31:0] requestBuffer_core_instruction; // @[peripheralUnit.scala 69:30]
  reg [3:0] requestBuffer_core_robAddr; // @[peripheralUnit.scala 69:30]
  reg [5:0] requestBuffer_core_prfDest; // @[peripheralUnit.scala 69:30]
  reg  requestBuffer_branch_valid; // @[peripheralUnit.scala 69:30]
  reg [4:0] requestBuffer_branch_mask; // @[peripheralUnit.scala 69:30]
  reg  requestBuffer_writeData_valid; // @[peripheralUnit.scala 69:30]
  reg [63:0] requestBuffer_writeData_data; // @[peripheralUnit.scala 69:30]
  reg  readRequestBuffer_valid; // @[peripheralUnit.scala 70:34]
  reg [31:0] readRequestBuffer_address; // @[peripheralUnit.scala 70:34]
  reg [31:0] readRequestBuffer_core_instruction; // @[peripheralUnit.scala 70:34]
  reg [3:0] readRequestBuffer_core_robAddr; // @[peripheralUnit.scala 70:34]
  reg [5:0] readRequestBuffer_core_prfDest; // @[peripheralUnit.scala 70:34]
  reg  readRequestBuffer_branch_valid; // @[peripheralUnit.scala 70:34]
  reg [4:0] readRequestBuffer_branch_mask; // @[peripheralUnit.scala 70:34]
  reg [63:0] readRequestBuffer_writeData_data; // @[peripheralUnit.scala 70:34]
  reg  writeRequestBuffer_valid; // @[peripheralUnit.scala 71:35]
  reg [31:0] writeRequestBuffer_address; // @[peripheralUnit.scala 71:35]
  reg [31:0] writeRequestBuffer_core_instruction; // @[peripheralUnit.scala 71:35]
  reg  writeRequestBuffer_branch_valid; // @[peripheralUnit.scala 71:35]
  reg [63:0] writeRequestBuffer_writeData_data; // @[peripheralUnit.scala 71:35]
  reg  responseOutBuffer_valid; // @[peripheralUnit.scala 73:34]
  reg [31:0] responseOutBuffer_address; // @[peripheralUnit.scala 73:34]
  reg [31:0] responseOutBuffer_core_instruction; // @[peripheralUnit.scala 73:34]
  reg [3:0] responseOutBuffer_core_robAddr; // @[peripheralUnit.scala 73:34]
  reg [5:0] responseOutBuffer_core_prfDest; // @[peripheralUnit.scala 73:34]
  reg  responseOutBuffer_branch_valid; // @[peripheralUnit.scala 73:34]
  reg [4:0] responseOutBuffer_branch_mask; // @[peripheralUnit.scala 73:34]
  reg [63:0] responseOutBuffer_writeData_data; // @[peripheralUnit.scala 73:34]
  reg  writeCommitInstructionBuffer; // @[peripheralUnit.scala 76:45]
  wire  _GEN_0 = writeInstructionCommit_fired ? 1'h0 : writeCommitInstructionBuffer; // @[peripheralUnit.scala 78:37 79:34 76:45]
  wire [4:0] _T_4 = requestBuffer_branch_mask & branchOps_branchMask; // @[utils.scala 62:31]
  wire  _T_5 = |_T_4; // @[utils.scala 62:55]
  wire [4:0] _readRequestBuffer_branch_mask_T = requestBuffer_branch_mask ^ branchOps_branchMask; // @[utils.scala 63:42]
  wire [4:0] _GEN_1 = |_T_4 ? _readRequestBuffer_branch_mask_T : requestBuffer_branch_mask; // @[utils.scala 62:60 63:23 65:23]
  wire  _GEN_2 = _T_5 ? 1'h0 : requestBuffer_branch_valid; // @[utils.scala 70:60 71:24 74:24]
  wire [4:0] _GEN_3 = _T_5 ? 5'h0 : requestBuffer_branch_mask; // @[utils.scala 70:60 72:23 75:23]
  wire [4:0] _GEN_4 = branchOps_passed ? _GEN_1 : _GEN_3; // @[utils.scala 60:30]
  wire  _GEN_5 = branchOps_passed ? requestBuffer_branch_valid : _GEN_2; // @[utils.scala 60:30 67:22]
  wire  _GEN_7 = branchOps_valid ? _GEN_5 : requestBuffer_branch_valid; // @[utils.scala 59:26 79:22]
  wire  _GEN_15 = ~writeRequestBuffer_valid & requestBuffer_writeData_valid & requestBuffer_branch_valid ?
    requestBuffer_valid : writeRequestBuffer_valid; // @[peripheralUnit.scala 97:105 99:26 71:35]
  wire  _GEN_28 = ~readRequestBuffer_valid & ~requestBuffer_writeData_valid ? requestBuffer_valid :
    readRequestBuffer_valid; // @[peripheralUnit.scala 92:69 94:25 70:34]
  wire  _GEN_41 = ~readRequestBuffer_valid & ~requestBuffer_writeData_valid ? writeRequestBuffer_valid : _GEN_15; // @[peripheralUnit.scala 71:35 92:69]
  wire  _GEN_66 = requestBuffer_valid & requestBuffer_branch_valid ? _GEN_28 : readRequestBuffer_valid; // @[peripheralUnit.scala 70:34 90:58]
  wire  _GEN_79 = requestBuffer_valid & requestBuffer_branch_valid ? _GEN_41 : writeRequestBuffer_valid; // @[peripheralUnit.scala 71:35 90:58]
  reg [1:0] writeAXIState; // @[peripheralUnit.scala 113:30]
  wire [1:0] sizeByIns = writeRequestBuffer_core_instruction[13:12]; // @[peripheralUnit.scala 123:58]
  wire [3:0] _sizePerBeat_T = 4'h1 << sizeByIns; // @[peripheralUnit.scala 124:30]
  wire [7:0] sizePerBeat = _sizePerBeat_T * 4'h8; // @[peripheralUnit.scala 124:44]
  wire [7:0] _bus_AWLEN_T_1 = sizePerBeat + 8'h20; // @[peripheralUnit.scala 129:34]
  wire [7:0] _bus_AWLEN_T_3 = _bus_AWLEN_T_1 - 8'h1; // @[peripheralUnit.scala 129:47]
  wire [7:0] _bus_AWLEN_T_4 = _bus_AWLEN_T_3 / 6'h20; // @[peripheralUnit.scala 129:54]
  wire [7:0] _bus_AWLEN_T_6 = _bus_AWLEN_T_4 - 8'h1; // @[peripheralUnit.scala 129:68]
  wire [5:0] _bus_AWSIZE_T_1 = 6'h20 / 4'h8; // @[peripheralUnit.scala 130:79]
  wire [1:0] bus_AWSIZE_hi = _bus_AWSIZE_T_1[5:4]; // @[CircuitMath.scala 33:17]
  wire [3:0] bus_AWSIZE_lo = _bus_AWSIZE_T_1[3:0]; // @[CircuitMath.scala 34:17]
  wire  bus_AWSIZE_useHi = |bus_AWSIZE_hi; // @[CircuitMath.scala 35:22]
  wire [1:0] _bus_AWSIZE_T_6 = bus_AWSIZE_lo[2] ? 2'h2 : {{1'd0}, bus_AWSIZE_lo[1]}; // @[CircuitMath.scala 30:10]
  wire [1:0] _bus_AWSIZE_T_7 = bus_AWSIZE_lo[3] ? 2'h3 : _bus_AWSIZE_T_6; // @[CircuitMath.scala 30:10]
  wire [1:0] _bus_AWSIZE_T_8 = bus_AWSIZE_useHi ? {{1'd0}, bus_AWSIZE_hi[1]} : _bus_AWSIZE_T_7; // @[CircuitMath.scala 36:21]
  wire [2:0] _bus_AWSIZE_T_9 = {bus_AWSIZE_useHi,_bus_AWSIZE_T_8}; // @[Cat.scala 33:92]
  wire [2:0] _bus_AWSIZE_T_10 = sizePerBeat <= 8'h20 ? {{1'd0}, sizeByIns} : _bus_AWSIZE_T_9; // @[peripheralUnit.scala 130:24]
  wire [7:0] _GEN_8 = {{7'd0}, writeCounter_count}; // @[peripheralUnit.scala 139:39]
  wire [31:0] writeChunks_0 = writeRequestBuffer_writeData_data[31:0]; // @[peripheralUnit.scala 143:42]
  wire [31:0] writeChunks_1 = writeRequestBuffer_writeData_data[63:32]; // @[peripheralUnit.scala 143:42]
  wire  _T_18 = bus_WREADY & bus_AWREADY; // @[peripheralUnit.scala 145:23]
  wire [31:0] _GEN_104 = writeCounter_count ? writeChunks_1 : writeChunks_0; // @[peripheralUnit.scala 148:{17,17}]
  wire  _writeRequestBuffer_valid_T_1 = bus_BVALID & bus_BID == 2'h0; // @[peripheralUnit.scala 153:48]
  wire  _writeRequestBuffer_valid_T_2 = bus_BRESP == 2'h0; // @[peripheralUnit.scala 153:81]
  wire [1:0] _writeAXIState_T_8 = _writeRequestBuffer_valid_T_2 ? 2'h0 : 2'h1; // @[peripheralUnit.scala 156:28]
  wire [1:0] _writeAXIState_T_9 = _writeRequestBuffer_valid_T_1 ? _writeAXIState_T_8 : 2'h2; // @[peripheralUnit.scala 155:27]
  wire  _GEN_107 = 2'h2 == writeAXIState | _GEN_0; // @[peripheralUnit.scala 117:25 154:36]
  wire [31:0] _GEN_111 = 2'h1 == writeAXIState ? writeRequestBuffer_address : 32'h0; // @[peripheralUnit.scala 117:25 128:18 38:14]
  wire [7:0] _GEN_112 = 2'h1 == writeAXIState ? _bus_AWLEN_T_6 : 8'h0; // @[peripheralUnit.scala 117:25 129:17 39:13]
  wire [2:0] _GEN_113 = 2'h1 == writeAXIState ? _bus_AWSIZE_T_10 : 3'h0; // @[peripheralUnit.scala 117:25 130:18 40:14]
  wire [1:0] _GEN_114 = 2'h1 == writeAXIState ? 2'h2 : 2'h0; // @[peripheralUnit.scala 117:25 134:18 44:14]
  wire [3:0] _GEN_115 = 2'h1 == writeAXIState ? 4'hf : 4'h0; // @[peripheralUnit.scala 117:25 138:17 49:13]
  wire  _GEN_116 = 2'h1 == writeAXIState & _GEN_8 == bus_ARLEN; // @[peripheralUnit.scala 117:25 139:17 50:13]
  wire [31:0] _GEN_118 = 2'h1 == writeAXIState ? _GEN_104 : 32'h0; // @[peripheralUnit.scala 117:25 148:17 48:13]
  wire  _GEN_120 = 2'h1 == writeAXIState ? 1'h0 : 2'h2 == writeAXIState; // @[peripheralUnit.scala 117:25 53:14]
  wire  _GEN_125 = 2'h0 == writeAXIState ? 1'h0 : 2'h1 == writeAXIState; // @[peripheralUnit.scala 117:25 46:15]
  wire [1:0] _GEN_130 = 2'h0 == writeAXIState ? 2'h0 : _GEN_114; // @[peripheralUnit.scala 117:25 44:14]
  reg  readAXIRequestState; // @[peripheralUnit.scala 163:36]
  wire [1:0] sizeByIns_1 = readRequestBuffer_core_instruction[13:12]; // @[peripheralUnit.scala 169:57]
  wire [3:0] _sizePerBeat_T_1 = 4'h1 << sizeByIns_1; // @[peripheralUnit.scala 170:30]
  wire [7:0] sizePerBeat_1 = _sizePerBeat_T_1 * 4'h8; // @[peripheralUnit.scala 170:44]
  wire [7:0] _bus_ARLEN_T_1 = sizePerBeat_1 + 8'h20; // @[peripheralUnit.scala 175:34]
  wire [7:0] _bus_ARLEN_T_3 = _bus_ARLEN_T_1 - 8'h1; // @[peripheralUnit.scala 175:47]
  wire [7:0] _bus_ARLEN_T_4 = _bus_ARLEN_T_3 / 6'h20; // @[peripheralUnit.scala 175:54]
  wire [7:0] _bus_ARLEN_T_6 = _bus_ARLEN_T_4 - 8'h1; // @[peripheralUnit.scala 175:68]
  wire [2:0] _bus_ARSIZE_T_10 = sizePerBeat_1 <= 8'h20 ? {{1'd0}, sizeByIns_1} : _bus_AWSIZE_T_9; // @[peripheralUnit.scala 176:24]
  wire [63:0] _GEN_141 = bus_ARREADY ? readRequestBuffer_writeData_data : 64'h0; // @[peripheralUnit.scala 185:24 186:35 utils.scala 49:41]
  wire [4:0] _GEN_143 = bus_ARREADY ? readRequestBuffer_branch_mask : 5'h0; // @[peripheralUnit.scala 185:24 186:35 utils.scala 49:41]
  wire  _GEN_144 = bus_ARREADY & readRequestBuffer_branch_valid; // @[peripheralUnit.scala 185:24 186:35 utils.scala 48:41]
  wire [5:0] _GEN_145 = bus_ARREADY ? readRequestBuffer_core_prfDest : 6'h0; // @[peripheralUnit.scala 185:24 186:35 utils.scala 49:41]
  wire [3:0] _GEN_146 = bus_ARREADY ? readRequestBuffer_core_robAddr : 4'h0; // @[peripheralUnit.scala 185:24 186:35 utils.scala 49:41]
  wire [31:0] _GEN_147 = bus_ARREADY ? readRequestBuffer_core_instruction : 32'h0; // @[peripheralUnit.scala 185:24 186:35 utils.scala 49:41]
  wire [31:0] _GEN_148 = bus_ARREADY ? readRequestBuffer_address : 32'h0; // @[peripheralUnit.scala 185:24 186:35 utils.scala 49:41]
  wire  _GEN_149 = bus_ARREADY & readRequestBuffer_valid; // @[peripheralUnit.scala 185:24 186:35 utils.scala 48:41]
  wire [31:0] _GEN_152 = readAXIRequestState ? readRequestBuffer_address : 32'h0; // @[peripheralUnit.scala 164:31 174:18 56:14]
  wire [7:0] _GEN_153 = readAXIRequestState ? _bus_ARLEN_T_6 : 8'h0; // @[peripheralUnit.scala 164:31 175:17 57:13]
  wire [2:0] _GEN_154 = readAXIRequestState ? _bus_ARSIZE_T_10 : 3'h0; // @[peripheralUnit.scala 164:31 176:18 58:14]
  wire [1:0] _GEN_155 = readAXIRequestState ? 2'h2 : 2'h0; // @[peripheralUnit.scala 164:31 180:18 62:14]
  wire [63:0] _GEN_160 = readAXIRequestState ? _GEN_141 : 64'h0; // @[peripheralUnit.scala 164:31 utils.scala 49:41]
  wire [4:0] _GEN_162 = readAXIRequestState ? _GEN_143 : 5'h0; // @[peripheralUnit.scala 164:31 utils.scala 49:41]
  wire [5:0] _GEN_164 = readAXIRequestState ? _GEN_145 : 6'h0; // @[peripheralUnit.scala 164:31 utils.scala 49:41]
  wire [3:0] _GEN_165 = readAXIRequestState ? _GEN_146 : 4'h0; // @[peripheralUnit.scala 164:31 utils.scala 49:41]
  wire [31:0] _GEN_166 = readAXIRequestState ? _GEN_147 : 32'h0; // @[peripheralUnit.scala 164:31 utils.scala 49:41]
  wire [31:0] _GEN_167 = readAXIRequestState ? _GEN_148 : 32'h0; // @[peripheralUnit.scala 164:31 utils.scala 49:41]
  wire  _GEN_171 = ~readAXIRequestState ? 1'h0 : readAXIRequestState; // @[peripheralUnit.scala 164:31 64:15]
  wire [1:0] _GEN_176 = ~readAXIRequestState ? 2'h0 : _GEN_155; // @[peripheralUnit.scala 164:31 62:14]
  reg [1:0] readAXIResponseState; // @[peripheralUnit.scala 194:37]
  reg [31:0] readDataVec_0; // @[peripheralUnit.scala 195:28]
  reg [31:0] readDataVec_1; // @[peripheralUnit.scala 195:28]
  reg  responseValid; // @[peripheralUnit.scala 196:30]
  wire  _T_23 = ~peripheralMSHR_isEmpty; // @[peripheralUnit.scala 204:12]
  wire  _T_26 = bus_RVALID & bus_RID == 2'h0; // @[peripheralUnit.scala 213:23]
  wire [31:0] _GEN_203 = ~readCounter_count ? bus_RDATA : readDataVec_0; // @[peripheralUnit.scala 195:28 215:{40,40}]
  wire [31:0] _GEN_204 = readCounter_count ? bus_RDATA : readDataVec_1; // @[peripheralUnit.scala 195:28 215:{40,40}]
  wire  _GEN_208 = bus_RVALID & bus_RID == 2'h0 ? bus_RRESP == 2'h0 & responseValid : responseValid; // @[peripheralUnit.scala 213:42 216:23 196:30]
  wire [63:0] doubleWordChoosen = {readDataVec_1,readDataVec_0}; // @[Cat.scala 33:92]
  wire [7:0] byteChunks_0 = doubleWordChoosen[7:0]; // @[peripheralUnit.scala 226:26]
  wire [7:0] byteChunks_1 = doubleWordChoosen[15:8]; // @[peripheralUnit.scala 226:26]
  wire [7:0] byteChunks_2 = doubleWordChoosen[23:16]; // @[peripheralUnit.scala 226:26]
  wire [7:0] byteChunks_3 = doubleWordChoosen[31:24]; // @[peripheralUnit.scala 226:26]
  wire [15:0] halfwordChoosed = {byteChunks_1,byteChunks_0}; // @[Cat.scala 33:92]
  wire [31:0] wordChoosed = {byteChunks_3,byteChunks_2,byteChunks_1,byteChunks_0}; // @[Cat.scala 33:92]
  wire [55:0] _responseOutBuffer_writeData_data_T_3 = byteChunks_0[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _responseOutBuffer_writeData_data_T_4 = {_responseOutBuffer_writeData_data_T_3,byteChunks_0}; // @[Cat.scala 33:92]
  wire [63:0] _responseOutBuffer_writeData_data_T_5 = responseOutBuffer_core_instruction[14] ? {{56'd0}, byteChunks_0}
     : _responseOutBuffer_writeData_data_T_4; // @[peripheralUnit.scala 232:60]
  wire [47:0] _responseOutBuffer_writeData_data_T_9 = halfwordChoosed[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _responseOutBuffer_writeData_data_T_10 = {_responseOutBuffer_writeData_data_T_9,byteChunks_1,byteChunks_0}
    ; // @[Cat.scala 33:92]
  wire [63:0] _responseOutBuffer_writeData_data_T_11 = responseOutBuffer_core_instruction[14] ? {{48'd0},
    halfwordChoosed} : _responseOutBuffer_writeData_data_T_10; // @[peripheralUnit.scala 234:60]
  wire [31:0] _responseOutBuffer_writeData_data_T_15 = wordChoosed[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _responseOutBuffer_writeData_data_T_16 = {_responseOutBuffer_writeData_data_T_15,byteChunks_3,byteChunks_2
    ,byteChunks_1,byteChunks_0}; // @[Cat.scala 33:92]
  wire [63:0] _responseOutBuffer_writeData_data_T_17 = responseOutBuffer_core_instruction[14] ? {{32'd0}, wordChoosed}
     : _responseOutBuffer_writeData_data_T_16; // @[peripheralUnit.scala 236:60]
  wire [63:0] _responseOutBuffer_writeData_data_T_19 = responseOutBuffer_core_instruction[14] ? 64'h0 :
    doubleWordChoosen; // @[peripheralUnit.scala 238:60]
  wire [63:0] _GEN_209 = 2'h3 == responseOutBuffer_core_instruction[13:12] ? _responseOutBuffer_writeData_data_T_19 :
    responseOutBuffer_writeData_data; // @[peripheralUnit.scala 231:57 238:54 73:34]
  wire [63:0] _GEN_210 = 2'h2 == responseOutBuffer_core_instruction[13:12] ? _responseOutBuffer_writeData_data_T_17 :
    _GEN_209; // @[peripheralUnit.scala 231:57 236:54]
  wire [63:0] _GEN_211 = 2'h1 == responseOutBuffer_core_instruction[13:12] ? _responseOutBuffer_writeData_data_T_11 :
    _GEN_210; // @[peripheralUnit.scala 231:57 234:54]
  wire [63:0] _GEN_212 = 2'h0 == responseOutBuffer_core_instruction[13:12] ? _responseOutBuffer_writeData_data_T_5 :
    _GEN_211; // @[peripheralUnit.scala 231:57 232:54]
  wire  _GEN_213 = responseOutBuffer_valid & responseOut_ready ? 1'h0 : 1'h1; // @[peripheralUnit.scala 241:31 242:57 243:33]
  wire [1:0] _readAXIResponseState_T_8 = responseOut_ready & responseOutBuffer_valid ? 2'h0 : 2'h2; // @[peripheralUnit.scala 245:34]
  wire  _GEN_221 = 2'h1 == readAXIResponseState ? _GEN_208 : responseValid; // @[peripheralUnit.scala 196:30 200:31]
  wire  _GEN_244 = 2'h0 == readAXIResponseState ? responseValid : _GEN_221; // @[peripheralUnit.scala 196:30 200:31]
  fifoBaseModule peripheralMSHR ( // @[peripheralUnit.scala 82:30]
    .clock(peripheralMSHR_clock),
    .reset(peripheralMSHR_reset),
    .write_ready(peripheralMSHR_write_ready),
    .write_data_valid(peripheralMSHR_write_data_valid),
    .write_data_address(peripheralMSHR_write_data_address),
    .write_data_core_instruction(peripheralMSHR_write_data_core_instruction),
    .write_data_core_robAddr(peripheralMSHR_write_data_core_robAddr),
    .write_data_core_prfDest(peripheralMSHR_write_data_core_prfDest),
    .write_data_branch_valid(peripheralMSHR_write_data_branch_valid),
    .write_data_branch_mask(peripheralMSHR_write_data_branch_mask),
    .write_data_writeData_data(peripheralMSHR_write_data_writeData_data),
    .read_ready(peripheralMSHR_read_ready),
    .read_data_valid(peripheralMSHR_read_data_valid),
    .read_data_address(peripheralMSHR_read_data_address),
    .read_data_core_instruction(peripheralMSHR_read_data_core_instruction),
    .read_data_core_robAddr(peripheralMSHR_read_data_core_robAddr),
    .read_data_core_prfDest(peripheralMSHR_read_data_core_prfDest),
    .read_data_branch_valid(peripheralMSHR_read_data_branch_valid),
    .read_data_branch_mask(peripheralMSHR_read_data_branch_mask),
    .read_data_writeData_data(peripheralMSHR_read_data_writeData_data),
    .isEmpty(peripheralMSHR_isEmpty)
  );
  moduleCounter writeCounter ( // @[peripheralUnit.scala 114:28]
    .clock(writeCounter_clock),
    .reset(writeCounter_reset),
    .count(writeCounter_count),
    .incrm(writeCounter_incrm)
  );
  moduleCounter readCounter ( // @[peripheralUnit.scala 197:27]
    .clock(readCounter_clock),
    .reset(readCounter_reset),
    .count(readCounter_count),
    .incrm(readCounter_incrm)
  );
  assign request_ready = requestBuffer_valid & requestBuffer_branch_valid ? 1'h0 : ~writeCommitInstructionBuffer; // @[peripheralUnit.scala 104:19 90:58 91:19]
  assign responseOut_request_valid = responseOutBuffer_valid; // @[peripheralUnit.scala 74:23]
  assign responseOut_request_address = responseOutBuffer_address; // @[peripheralUnit.scala 74:23]
  assign responseOut_request_core_instruction = responseOutBuffer_core_instruction; // @[peripheralUnit.scala 74:23]
  assign responseOut_request_core_robAddr = responseOutBuffer_core_robAddr; // @[peripheralUnit.scala 74:23]
  assign responseOut_request_core_prfDest = responseOutBuffer_core_prfDest; // @[peripheralUnit.scala 74:23]
  assign responseOut_request_branch_valid = responseOutBuffer_branch_valid; // @[peripheralUnit.scala 74:23]
  assign responseOut_request_branch_mask = responseOutBuffer_branch_mask; // @[peripheralUnit.scala 74:23]
  assign responseOut_request_writeData_data = responseOutBuffer_writeData_data; // @[peripheralUnit.scala 74:23]
  assign bus_AWADDR = 2'h0 == writeAXIState ? 32'h0 : _GEN_111; // @[peripheralUnit.scala 117:25 38:14]
  assign bus_AWLEN = 2'h0 == writeAXIState ? 8'h0 : _GEN_112; // @[peripheralUnit.scala 117:25 39:13]
  assign bus_AWSIZE = 2'h0 == writeAXIState ? 3'h0 : _GEN_113; // @[peripheralUnit.scala 117:25 40:14]
  assign bus_AWBURST = {{1'd0}, _GEN_125};
  assign bus_AWPROT = {{1'd0}, _GEN_130};
  assign bus_AWVALID = 2'h0 == writeAXIState ? 1'h0 : 2'h1 == writeAXIState; // @[peripheralUnit.scala 117:25 46:15]
  assign bus_WDATA = 2'h0 == writeAXIState ? 32'h0 : _GEN_118; // @[peripheralUnit.scala 117:25 48:13]
  assign bus_WSTRB = 2'h0 == writeAXIState ? 4'h0 : _GEN_115; // @[peripheralUnit.scala 117:25 49:13]
  assign bus_WLAST = 2'h0 == writeAXIState ? 1'h0 : _GEN_116; // @[peripheralUnit.scala 117:25 50:13]
  assign bus_WVALID = 2'h0 == writeAXIState ? 1'h0 : 2'h1 == writeAXIState; // @[peripheralUnit.scala 117:25 46:15]
  assign bus_BREADY = 2'h0 == writeAXIState ? 1'h0 : _GEN_120; // @[peripheralUnit.scala 117:25 53:14]
  assign bus_ARADDR = ~readAXIRequestState ? 32'h0 : _GEN_152; // @[peripheralUnit.scala 164:31 56:14]
  assign bus_ARLEN = ~readAXIRequestState ? 8'h0 : _GEN_153; // @[peripheralUnit.scala 164:31 57:13]
  assign bus_ARSIZE = ~readAXIRequestState ? 3'h0 : _GEN_154; // @[peripheralUnit.scala 164:31 58:14]
  assign bus_ARBURST = {{1'd0}, _GEN_171};
  assign bus_ARPROT = {{1'd0}, _GEN_176};
  assign bus_ARVALID = ~readAXIRequestState ? 1'h0 : readAXIRequestState; // @[peripheralUnit.scala 164:31 64:15]
  assign bus_RREADY = 2'h0 == readAXIResponseState ? 1'h0 : 2'h1 == readAXIResponseState; // @[peripheralUnit.scala 200:31 66:14]
  assign writeInstructionCommit_ready = writeCommitInstructionBuffer; // @[peripheralUnit.scala 77:32]
  assign peripheralMSHR_clock = clock;
  assign peripheralMSHR_reset = reset;
  assign peripheralMSHR_write_data_valid = ~readAXIRequestState ? 1'h0 : readAXIRequestState & _GEN_149; // @[peripheralUnit.scala 164:31 utils.scala 48:41]
  assign peripheralMSHR_write_data_address = ~readAXIRequestState ? 32'h0 : _GEN_167; // @[peripheralUnit.scala 164:31 utils.scala 49:41]
  assign peripheralMSHR_write_data_core_instruction = ~readAXIRequestState ? 32'h0 : _GEN_166; // @[peripheralUnit.scala 164:31 utils.scala 49:41]
  assign peripheralMSHR_write_data_core_robAddr = ~readAXIRequestState ? 4'h0 : _GEN_165; // @[peripheralUnit.scala 164:31 utils.scala 49:41]
  assign peripheralMSHR_write_data_core_prfDest = ~readAXIRequestState ? 6'h0 : _GEN_164; // @[peripheralUnit.scala 164:31 utils.scala 49:41]
  assign peripheralMSHR_write_data_branch_valid = ~readAXIRequestState ? 1'h0 : readAXIRequestState & _GEN_144; // @[peripheralUnit.scala 164:31 utils.scala 48:41]
  assign peripheralMSHR_write_data_branch_mask = ~readAXIRequestState ? 5'h0 : _GEN_162; // @[peripheralUnit.scala 164:31 utils.scala 49:41]
  assign peripheralMSHR_write_data_writeData_data = ~readAXIRequestState ? 64'h0 : _GEN_160; // @[peripheralUnit.scala 164:31 utils.scala 49:41]
  assign peripheralMSHR_read_ready = 2'h0 == readAXIResponseState & _T_23; // @[peripheralUnit.scala 200:31 87:29]
  assign writeCounter_clock = clock;
  assign writeCounter_reset = 2'h0 == writeAXIState; // @[peripheralUnit.scala 117:25]
  assign writeCounter_incrm = 2'h0 == writeAXIState ? 1'h0 : 2'h1 == writeAXIState & _T_18; // @[peripheralUnit.scala 115:22 117:25]
  assign readCounter_clock = clock;
  assign readCounter_reset = 2'h0 == readAXIResponseState; // @[peripheralUnit.scala 200:31]
  assign readCounter_incrm = 2'h0 == readAXIResponseState ? 1'h0 : 2'h1 == readAXIResponseState & _T_26; // @[peripheralUnit.scala 198:21 200:31]
  always @(posedge clock) begin
    if (reset) begin // @[peripheralUnit.scala 69:30]
      requestBuffer_valid <= 1'h0; // @[peripheralUnit.scala 69:30]
    end else if (requestBuffer_valid & requestBuffer_branch_valid) begin // @[peripheralUnit.scala 90:58]
      if (~readRequestBuffer_valid & ~requestBuffer_writeData_valid) begin // @[peripheralUnit.scala 92:69]
        requestBuffer_valid <= 1'h0; // @[peripheralUnit.scala 96:27]
      end else if (~writeRequestBuffer_valid & requestBuffer_writeData_valid & requestBuffer_branch_valid) begin // @[peripheralUnit.scala 97:105]
        requestBuffer_valid <= 1'h0; // @[peripheralUnit.scala 101:27]
      end
    end else if (request_request_valid & request_request_branch_valid) begin // @[peripheralUnit.scala 105:64]
      requestBuffer_valid <= request_request_valid; // @[peripheralUnit.scala 106:21]
    end
    if (reset) begin // @[peripheralUnit.scala 69:30]
      requestBuffer_address <= 32'h0; // @[peripheralUnit.scala 69:30]
    end else if (!(requestBuffer_valid & requestBuffer_branch_valid)) begin // @[peripheralUnit.scala 90:58]
      if (request_request_valid & request_request_branch_valid) begin // @[peripheralUnit.scala 105:64]
        requestBuffer_address <= request_request_address; // @[peripheralUnit.scala 106:21]
      end
    end
    if (reset) begin // @[peripheralUnit.scala 69:30]
      requestBuffer_core_instruction <= 32'h0; // @[peripheralUnit.scala 69:30]
    end else if (!(requestBuffer_valid & requestBuffer_branch_valid)) begin // @[peripheralUnit.scala 90:58]
      if (request_request_valid & request_request_branch_valid) begin // @[peripheralUnit.scala 105:64]
        requestBuffer_core_instruction <= request_request_core_instruction; // @[peripheralUnit.scala 106:21]
      end
    end
    if (reset) begin // @[peripheralUnit.scala 69:30]
      requestBuffer_core_robAddr <= 4'h0; // @[peripheralUnit.scala 69:30]
    end else if (!(requestBuffer_valid & requestBuffer_branch_valid)) begin // @[peripheralUnit.scala 90:58]
      if (request_request_valid & request_request_branch_valid) begin // @[peripheralUnit.scala 105:64]
        requestBuffer_core_robAddr <= request_request_core_robAddr; // @[peripheralUnit.scala 106:21]
      end
    end
    if (reset) begin // @[peripheralUnit.scala 69:30]
      requestBuffer_core_prfDest <= 6'h0; // @[peripheralUnit.scala 69:30]
    end else if (!(requestBuffer_valid & requestBuffer_branch_valid)) begin // @[peripheralUnit.scala 90:58]
      if (request_request_valid & request_request_branch_valid) begin // @[peripheralUnit.scala 105:64]
        requestBuffer_core_prfDest <= request_request_core_prfDest; // @[peripheralUnit.scala 106:21]
      end
    end
    if (reset) begin // @[peripheralUnit.scala 69:30]
      requestBuffer_branch_valid <= 1'h0; // @[peripheralUnit.scala 69:30]
    end else if (!(requestBuffer_valid & requestBuffer_branch_valid)) begin // @[peripheralUnit.scala 90:58]
      if (request_request_valid & request_request_branch_valid) begin // @[peripheralUnit.scala 105:64]
        requestBuffer_branch_valid <= request_request_branch_valid; // @[peripheralUnit.scala 106:21]
      end
    end
    if (reset) begin // @[peripheralUnit.scala 69:30]
      requestBuffer_branch_mask <= 5'h0; // @[peripheralUnit.scala 69:30]
    end else if (!(requestBuffer_valid & requestBuffer_branch_valid)) begin // @[peripheralUnit.scala 90:58]
      if (request_request_valid & request_request_branch_valid) begin // @[peripheralUnit.scala 105:64]
        requestBuffer_branch_mask <= request_request_branch_mask; // @[peripheralUnit.scala 106:21]
      end
    end
    if (reset) begin // @[peripheralUnit.scala 69:30]
      requestBuffer_writeData_valid <= 1'h0; // @[peripheralUnit.scala 69:30]
    end else if (!(requestBuffer_valid & requestBuffer_branch_valid)) begin // @[peripheralUnit.scala 90:58]
      if (request_request_valid & request_request_branch_valid) begin // @[peripheralUnit.scala 105:64]
        requestBuffer_writeData_valid <= request_request_writeData_valid; // @[peripheralUnit.scala 106:21]
      end
    end
    if (reset) begin // @[peripheralUnit.scala 69:30]
      requestBuffer_writeData_data <= 64'h0; // @[peripheralUnit.scala 69:30]
    end else if (!(requestBuffer_valid & requestBuffer_branch_valid)) begin // @[peripheralUnit.scala 90:58]
      if (request_request_valid & request_request_branch_valid) begin // @[peripheralUnit.scala 105:64]
        requestBuffer_writeData_data <= request_request_writeData_data; // @[peripheralUnit.scala 106:21]
      end
    end
    if (reset) begin // @[peripheralUnit.scala 70:34]
      readRequestBuffer_valid <= 1'h0; // @[peripheralUnit.scala 70:34]
    end else if (~readAXIRequestState) begin // @[peripheralUnit.scala 164:31]
      readRequestBuffer_valid <= _GEN_66;
    end else if (readAXIRequestState) begin // @[peripheralUnit.scala 164:31]
      readRequestBuffer_valid <= ~bus_ARREADY; // @[peripheralUnit.scala 183:31]
    end else begin
      readRequestBuffer_valid <= _GEN_66;
    end
    if (reset) begin // @[peripheralUnit.scala 70:34]
      readRequestBuffer_address <= 32'h0; // @[peripheralUnit.scala 70:34]
    end else if (requestBuffer_valid & requestBuffer_branch_valid) begin // @[peripheralUnit.scala 90:58]
      if (~readRequestBuffer_valid & ~requestBuffer_writeData_valid) begin // @[peripheralUnit.scala 92:69]
        readRequestBuffer_address <= requestBuffer_address; // @[peripheralUnit.scala 94:25]
      end
    end
    if (reset) begin // @[peripheralUnit.scala 70:34]
      readRequestBuffer_core_instruction <= 32'h0; // @[peripheralUnit.scala 70:34]
    end else if (requestBuffer_valid & requestBuffer_branch_valid) begin // @[peripheralUnit.scala 90:58]
      if (~readRequestBuffer_valid & ~requestBuffer_writeData_valid) begin // @[peripheralUnit.scala 92:69]
        readRequestBuffer_core_instruction <= requestBuffer_core_instruction; // @[peripheralUnit.scala 94:25]
      end
    end
    if (reset) begin // @[peripheralUnit.scala 70:34]
      readRequestBuffer_core_robAddr <= 4'h0; // @[peripheralUnit.scala 70:34]
    end else if (requestBuffer_valid & requestBuffer_branch_valid) begin // @[peripheralUnit.scala 90:58]
      if (~readRequestBuffer_valid & ~requestBuffer_writeData_valid) begin // @[peripheralUnit.scala 92:69]
        readRequestBuffer_core_robAddr <= requestBuffer_core_robAddr; // @[peripheralUnit.scala 94:25]
      end
    end
    if (reset) begin // @[peripheralUnit.scala 70:34]
      readRequestBuffer_core_prfDest <= 6'h0; // @[peripheralUnit.scala 70:34]
    end else if (requestBuffer_valid & requestBuffer_branch_valid) begin // @[peripheralUnit.scala 90:58]
      if (~readRequestBuffer_valid & ~requestBuffer_writeData_valid) begin // @[peripheralUnit.scala 92:69]
        readRequestBuffer_core_prfDest <= requestBuffer_core_prfDest; // @[peripheralUnit.scala 94:25]
      end
    end
    if (reset) begin // @[peripheralUnit.scala 70:34]
      readRequestBuffer_branch_valid <= 1'h0; // @[peripheralUnit.scala 70:34]
    end else if (requestBuffer_valid & requestBuffer_branch_valid) begin // @[peripheralUnit.scala 90:58]
      if (~readRequestBuffer_valid & ~requestBuffer_writeData_valid) begin // @[peripheralUnit.scala 92:69]
        if (branchOps_valid) begin // @[utils.scala 59:26]
          readRequestBuffer_branch_valid <= _GEN_5;
        end else begin
          readRequestBuffer_branch_valid <= requestBuffer_branch_valid; // @[utils.scala 79:22]
        end
      end
    end
    if (reset) begin // @[peripheralUnit.scala 70:34]
      readRequestBuffer_branch_mask <= 5'h0; // @[peripheralUnit.scala 70:34]
    end else if (requestBuffer_valid & requestBuffer_branch_valid) begin // @[peripheralUnit.scala 90:58]
      if (~readRequestBuffer_valid & ~requestBuffer_writeData_valid) begin // @[peripheralUnit.scala 92:69]
        if (branchOps_valid) begin // @[utils.scala 59:26]
          readRequestBuffer_branch_mask <= _GEN_4;
        end else begin
          readRequestBuffer_branch_mask <= requestBuffer_branch_mask; // @[utils.scala 80:21]
        end
      end
    end
    if (reset) begin // @[peripheralUnit.scala 70:34]
      readRequestBuffer_writeData_data <= 64'h0; // @[peripheralUnit.scala 70:34]
    end else if (requestBuffer_valid & requestBuffer_branch_valid) begin // @[peripheralUnit.scala 90:58]
      if (~readRequestBuffer_valid & ~requestBuffer_writeData_valid) begin // @[peripheralUnit.scala 92:69]
        readRequestBuffer_writeData_data <= requestBuffer_writeData_data; // @[peripheralUnit.scala 94:25]
      end
    end
    if (reset) begin // @[peripheralUnit.scala 71:35]
      writeRequestBuffer_valid <= 1'h0; // @[peripheralUnit.scala 71:35]
    end else if (2'h0 == writeAXIState) begin // @[peripheralUnit.scala 117:25]
      writeRequestBuffer_valid <= _GEN_79;
    end else if (2'h1 == writeAXIState) begin // @[peripheralUnit.scala 117:25]
      writeRequestBuffer_valid <= _GEN_79;
    end else if (2'h2 == writeAXIState) begin // @[peripheralUnit.scala 117:25]
      writeRequestBuffer_valid <= ~(bus_BVALID & bus_BID == 2'h0 & bus_BRESP == 2'h0); // @[peripheralUnit.scala 153:32]
    end else begin
      writeRequestBuffer_valid <= _GEN_79;
    end
    if (reset) begin // @[peripheralUnit.scala 71:35]
      writeRequestBuffer_address <= 32'h0; // @[peripheralUnit.scala 71:35]
    end else if (requestBuffer_valid & requestBuffer_branch_valid) begin // @[peripheralUnit.scala 90:58]
      if (!(~readRequestBuffer_valid & ~requestBuffer_writeData_valid)) begin // @[peripheralUnit.scala 92:69]
        if (~writeRequestBuffer_valid & requestBuffer_writeData_valid & requestBuffer_branch_valid) begin // @[peripheralUnit.scala 97:105]
          writeRequestBuffer_address <= requestBuffer_address; // @[peripheralUnit.scala 99:26]
        end
      end
    end
    if (reset) begin // @[peripheralUnit.scala 71:35]
      writeRequestBuffer_core_instruction <= 32'h0; // @[peripheralUnit.scala 71:35]
    end else if (requestBuffer_valid & requestBuffer_branch_valid) begin // @[peripheralUnit.scala 90:58]
      if (!(~readRequestBuffer_valid & ~requestBuffer_writeData_valid)) begin // @[peripheralUnit.scala 92:69]
        if (~writeRequestBuffer_valid & requestBuffer_writeData_valid & requestBuffer_branch_valid) begin // @[peripheralUnit.scala 97:105]
          writeRequestBuffer_core_instruction <= requestBuffer_core_instruction; // @[peripheralUnit.scala 99:26]
        end
      end
    end
    if (reset) begin // @[peripheralUnit.scala 71:35]
      writeRequestBuffer_branch_valid <= 1'h0; // @[peripheralUnit.scala 71:35]
    end else if (requestBuffer_valid & requestBuffer_branch_valid) begin // @[peripheralUnit.scala 90:58]
      if (!(~readRequestBuffer_valid & ~requestBuffer_writeData_valid)) begin // @[peripheralUnit.scala 92:69]
        if (~writeRequestBuffer_valid & requestBuffer_writeData_valid & requestBuffer_branch_valid) begin // @[peripheralUnit.scala 97:105]
          writeRequestBuffer_branch_valid <= _GEN_7;
        end
      end
    end
    if (reset) begin // @[peripheralUnit.scala 71:35]
      writeRequestBuffer_writeData_data <= 64'h0; // @[peripheralUnit.scala 71:35]
    end else if (requestBuffer_valid & requestBuffer_branch_valid) begin // @[peripheralUnit.scala 90:58]
      if (!(~readRequestBuffer_valid & ~requestBuffer_writeData_valid)) begin // @[peripheralUnit.scala 92:69]
        if (~writeRequestBuffer_valid & requestBuffer_writeData_valid & requestBuffer_branch_valid) begin // @[peripheralUnit.scala 97:105]
          writeRequestBuffer_writeData_data <= requestBuffer_writeData_data; // @[peripheralUnit.scala 99:26]
        end
      end
    end
    if (reset) begin // @[peripheralUnit.scala 73:34]
      responseOutBuffer_valid <= 1'h0; // @[peripheralUnit.scala 73:34]
    end else if (2'h0 == readAXIResponseState) begin // @[peripheralUnit.scala 200:31]
      responseOutBuffer_valid <= 1'h0; // @[peripheralUnit.scala 208:31]
    end else if (!(2'h1 == readAXIResponseState)) begin // @[peripheralUnit.scala 200:31]
      if (2'h2 == readAXIResponseState) begin // @[peripheralUnit.scala 200:31]
        responseOutBuffer_valid <= _GEN_213;
      end
    end
    if (reset) begin // @[peripheralUnit.scala 73:34]
      responseOutBuffer_address <= 32'h0; // @[peripheralUnit.scala 73:34]
    end else if (2'h0 == readAXIResponseState) begin // @[peripheralUnit.scala 200:31]
      if (~peripheralMSHR_isEmpty) begin // @[peripheralUnit.scala 204:36]
        responseOutBuffer_address <= peripheralMSHR_read_data_address; // @[peripheralUnit.scala 206:27]
      end
    end
    if (reset) begin // @[peripheralUnit.scala 73:34]
      responseOutBuffer_core_instruction <= 32'h0; // @[peripheralUnit.scala 73:34]
    end else if (2'h0 == readAXIResponseState) begin // @[peripheralUnit.scala 200:31]
      if (~peripheralMSHR_isEmpty) begin // @[peripheralUnit.scala 204:36]
        responseOutBuffer_core_instruction <= peripheralMSHR_read_data_core_instruction; // @[peripheralUnit.scala 206:27]
      end
    end
    if (reset) begin // @[peripheralUnit.scala 73:34]
      responseOutBuffer_core_robAddr <= 4'h0; // @[peripheralUnit.scala 73:34]
    end else if (2'h0 == readAXIResponseState) begin // @[peripheralUnit.scala 200:31]
      if (~peripheralMSHR_isEmpty) begin // @[peripheralUnit.scala 204:36]
        responseOutBuffer_core_robAddr <= peripheralMSHR_read_data_core_robAddr; // @[peripheralUnit.scala 206:27]
      end
    end
    if (reset) begin // @[peripheralUnit.scala 73:34]
      responseOutBuffer_core_prfDest <= 6'h0; // @[peripheralUnit.scala 73:34]
    end else if (2'h0 == readAXIResponseState) begin // @[peripheralUnit.scala 200:31]
      if (~peripheralMSHR_isEmpty) begin // @[peripheralUnit.scala 204:36]
        responseOutBuffer_core_prfDest <= peripheralMSHR_read_data_core_prfDest; // @[peripheralUnit.scala 206:27]
      end
    end
    if (reset) begin // @[peripheralUnit.scala 73:34]
      responseOutBuffer_branch_valid <= 1'h0; // @[peripheralUnit.scala 73:34]
    end else if (2'h0 == readAXIResponseState) begin // @[peripheralUnit.scala 200:31]
      if (~peripheralMSHR_isEmpty) begin // @[peripheralUnit.scala 204:36]
        responseOutBuffer_branch_valid <= peripheralMSHR_read_data_branch_valid; // @[peripheralUnit.scala 206:27]
      end
    end
    if (reset) begin // @[peripheralUnit.scala 73:34]
      responseOutBuffer_branch_mask <= 5'h0; // @[peripheralUnit.scala 73:34]
    end else if (2'h0 == readAXIResponseState) begin // @[peripheralUnit.scala 200:31]
      if (~peripheralMSHR_isEmpty) begin // @[peripheralUnit.scala 204:36]
        responseOutBuffer_branch_mask <= peripheralMSHR_read_data_branch_mask; // @[peripheralUnit.scala 206:27]
      end
    end
    if (reset) begin // @[peripheralUnit.scala 73:34]
      responseOutBuffer_writeData_data <= 64'h0; // @[peripheralUnit.scala 73:34]
    end else if (2'h0 == readAXIResponseState) begin // @[peripheralUnit.scala 200:31]
      if (~peripheralMSHR_isEmpty) begin // @[peripheralUnit.scala 204:36]
        responseOutBuffer_writeData_data <= peripheralMSHR_read_data_writeData_data; // @[peripheralUnit.scala 206:27]
      end
    end else if (!(2'h1 == readAXIResponseState)) begin // @[peripheralUnit.scala 200:31]
      if (2'h2 == readAXIResponseState) begin // @[peripheralUnit.scala 200:31]
        responseOutBuffer_writeData_data <= _GEN_212;
      end
    end
    if (reset) begin // @[peripheralUnit.scala 76:45]
      writeCommitInstructionBuffer <= 1'h0; // @[peripheralUnit.scala 76:45]
    end else if (2'h0 == writeAXIState) begin // @[peripheralUnit.scala 117:25]
      writeCommitInstructionBuffer <= _GEN_0;
    end else if (2'h1 == writeAXIState) begin // @[peripheralUnit.scala 117:25]
      writeCommitInstructionBuffer <= _GEN_0;
    end else begin
      writeCommitInstructionBuffer <= _GEN_107;
    end
    if (reset) begin // @[peripheralUnit.scala 113:30]
      writeAXIState <= 2'h0; // @[peripheralUnit.scala 113:30]
    end else if (2'h0 == writeAXIState) begin // @[peripheralUnit.scala 117:25]
      if (writeRequestBuffer_valid & writeRequestBuffer_branch_valid) begin // @[peripheralUnit.scala 120:29]
        writeAXIState <= 2'h1;
      end else begin
        writeAXIState <= 2'h0;
      end
    end else if (2'h1 == writeAXIState) begin // @[peripheralUnit.scala 117:25]
      if (bus_WLAST & bus_WREADY & bus_AWREADY) begin // @[peripheralUnit.scala 149:27]
        writeAXIState <= 2'h2;
      end else begin
        writeAXIState <= 2'h1;
      end
    end else if (2'h2 == writeAXIState) begin // @[peripheralUnit.scala 117:25]
      writeAXIState <= _writeAXIState_T_9; // @[peripheralUnit.scala 155:21]
    end
    if (reset) begin // @[peripheralUnit.scala 163:36]
      readAXIRequestState <= 1'h0; // @[peripheralUnit.scala 163:36]
    end else if (~readAXIRequestState) begin // @[peripheralUnit.scala 164:31]
      readAXIRequestState <= readRequestBuffer_valid & readRequestBuffer_branch_valid & peripheralMSHR_write_ready; // @[peripheralUnit.scala 166:27]
    end else if (readAXIRequestState) begin // @[peripheralUnit.scala 164:31]
      if (bus_ARREADY) begin // @[peripheralUnit.scala 188:33]
        readAXIRequestState <= 1'h0;
      end else begin
        readAXIRequestState <= 1'h1;
      end
    end
    if (reset) begin // @[peripheralUnit.scala 194:37]
      readAXIResponseState <= 2'h0; // @[peripheralUnit.scala 194:37]
    end else if (2'h0 == readAXIResponseState) begin // @[peripheralUnit.scala 200:31]
      if (peripheralMSHR_read_data_valid & peripheralMSHR_read_data_branch_valid & _T_23) begin // @[peripheralUnit.scala 209:34]
        readAXIResponseState <= 2'h1;
      end else begin
        readAXIResponseState <= 2'h0;
      end
    end else if (2'h1 == readAXIResponseState) begin // @[peripheralUnit.scala 200:31]
      if (bus_RLAST & bus_RVALID & responseValid) begin // @[peripheralUnit.scala 219:34]
        readAXIResponseState <= 2'h2;
      end else begin
        readAXIResponseState <= 2'h1;
      end
    end else if (2'h2 == readAXIResponseState) begin // @[peripheralUnit.scala 200:31]
      readAXIResponseState <= _readAXIResponseState_T_8; // @[peripheralUnit.scala 245:28]
    end
    if (reset) begin // @[peripheralUnit.scala 195:28]
      readDataVec_0 <= 32'h0; // @[peripheralUnit.scala 195:28]
    end else if (!(2'h0 == readAXIResponseState)) begin // @[peripheralUnit.scala 200:31]
      if (2'h1 == readAXIResponseState) begin // @[peripheralUnit.scala 200:31]
        if (bus_RVALID & bus_RID == 2'h0) begin // @[peripheralUnit.scala 213:42]
          readDataVec_0 <= _GEN_203;
        end
      end
    end
    if (reset) begin // @[peripheralUnit.scala 195:28]
      readDataVec_1 <= 32'h0; // @[peripheralUnit.scala 195:28]
    end else if (!(2'h0 == readAXIResponseState)) begin // @[peripheralUnit.scala 200:31]
      if (2'h1 == readAXIResponseState) begin // @[peripheralUnit.scala 200:31]
        if (bus_RVALID & bus_RID == 2'h0) begin // @[peripheralUnit.scala 213:42]
          readDataVec_1 <= _GEN_204;
        end
      end
    end
    responseValid <= reset | _GEN_244; // @[peripheralUnit.scala 196:{30,30}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  requestBuffer_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  requestBuffer_address = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  requestBuffer_core_instruction = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  requestBuffer_core_robAddr = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  requestBuffer_core_prfDest = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  requestBuffer_branch_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  requestBuffer_branch_mask = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  requestBuffer_writeData_valid = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  requestBuffer_writeData_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  readRequestBuffer_valid = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  readRequestBuffer_address = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  readRequestBuffer_core_instruction = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  readRequestBuffer_core_robAddr = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  readRequestBuffer_core_prfDest = _RAND_13[5:0];
  _RAND_14 = {1{`RANDOM}};
  readRequestBuffer_branch_valid = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  readRequestBuffer_branch_mask = _RAND_15[4:0];
  _RAND_16 = {2{`RANDOM}};
  readRequestBuffer_writeData_data = _RAND_16[63:0];
  _RAND_17 = {1{`RANDOM}};
  writeRequestBuffer_valid = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  writeRequestBuffer_address = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  writeRequestBuffer_core_instruction = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  writeRequestBuffer_branch_valid = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  writeRequestBuffer_writeData_data = _RAND_21[63:0];
  _RAND_22 = {1{`RANDOM}};
  responseOutBuffer_valid = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  responseOutBuffer_address = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  responseOutBuffer_core_instruction = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  responseOutBuffer_core_robAddr = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  responseOutBuffer_core_prfDest = _RAND_26[5:0];
  _RAND_27 = {1{`RANDOM}};
  responseOutBuffer_branch_valid = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  responseOutBuffer_branch_mask = _RAND_28[4:0];
  _RAND_29 = {2{`RANDOM}};
  responseOutBuffer_writeData_data = _RAND_29[63:0];
  _RAND_30 = {1{`RANDOM}};
  writeCommitInstructionBuffer = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  writeAXIState = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  readAXIRequestState = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  readAXIResponseState = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  readDataVec_0 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  readDataVec_1 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  responseValid = _RAND_36[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module moduleCounter_2(
  input        clock,
  input        reset,
  output [2:0] count,
  input        incrm
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] cntReg; // @[utils.scala 17:23]
  wire [2:0] _cntReg_T_3 = cntReg + 3'h1; // @[utils.scala 19:35]
  assign count = cntReg; // @[utils.scala 20:9]
  always @(posedge clock) begin
    if (reset) begin // @[utils.scala 17:23]
      cntReg <= 3'h0; // @[utils.scala 17:23]
    end else if (incrm & cntReg == 3'h7) begin // @[utils.scala 18:16]
      cntReg <= 3'h0;
    end else if (incrm) begin // @[utils.scala 19:20]
      cntReg <= _cntReg_T_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cntReg = _RAND_0[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ACEUnit(
  input          clock,
  input          reset,
  output         readRequest_ready,
  input          readRequest_request_valid,
  input  [31:0]  readRequest_request_address,
  input  [31:0]  readRequest_request_core_instruction,
  input  [3:0]   readRequest_request_core_robAddr,
  input  [5:0]   readRequest_request_core_prfDest,
  input          readRequest_request_branch_valid,
  input  [4:0]   readRequest_request_branch_mask,
  input          readRequest_request_writeData_valid,
  input  [63:0]  readRequest_request_writeData_data,
  input  [1:0]   readRequest_request_cacheLine_response,
  input          readResponse_ready,
  output         readResponse_request_valid,
  output [31:0]  readResponse_request_address,
  output [31:0]  readResponse_request_core_instruction,
  output [3:0]   readResponse_request_core_robAddr,
  output [5:0]   readResponse_request_core_prfDest,
  output         readResponse_request_branch_valid,
  output [4:0]   readResponse_request_branch_mask,
  output         readResponse_request_writeData_valid,
  output [63:0]  readResponse_request_writeData_data,
  output [511:0] readResponse_request_cacheLine_cacheLine,
  output [1:0]   readResponse_request_cacheLine_response,
  output         writeRequest_ready,
  input          writeRequest_request_valid,
  input  [31:0]  writeRequest_request_address,
  input  [511:0] writeRequest_request_data,
  input          coherencyRequest_ready,
  output         coherencyRequest_request_valid,
  output [31:0]  coherencyRequest_request_address,
  output [1:0]   coherencyRequest_request_response,
  output         coherencyResponse_ready,
  input          coherencyResponse_request_valid,
  input  [1:0]   coherencyResponse_request_response,
  input  [511:0] coherencyResponse_request_cacheLine,
  input          coherencyResponse_request_dataValid,
  output         fenceReady,
  input          branchOps_valid,
  input  [4:0]   branchOps_branchMask,
  input          branchOps_passed,
  output [31:0]  bus_AWADDR,
  output         bus_AWVALID,
  input          bus_AWREADY,
  output [63:0]  bus_WDATA,
  output         bus_WLAST,
  output         bus_WVALID,
  input          bus_WREADY,
  input  [1:0]   bus_BRESP,
  input          bus_BVALID,
  output         bus_BREADY,
  output [31:0]  bus_ARADDR,
  output         bus_ARVALID,
  input          bus_ARREADY,
  input  [63:0]  bus_RDATA,
  input          bus_RLAST,
  input          bus_RVALID,
  output         bus_RREADY,
  output [2:0]   bus_AWSNOOP,
  output [3:0]   bus_ARSNOOP,
  input  [3:0]   bus_RRESP,
  input          bus_ACVALID,
  output         bus_ACREADY,
  input  [31:0]  bus_ACADDR,
  input  [3:0]   bus_ACSNOOP,
  output         bus_CRVALID,
  input          bus_CRREADY,
  output [4:0]   bus_CRRESP,
  output         bus_CDVALID,
  input          bus_CDREADY,
  output [63:0]  bus_CDDATA,
  output         bus_CDLAST
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [511:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [511:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [511:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
`endif // RANDOMIZE_REG_INIT
  wire  ACEMSHR_clock; // @[ACEUnit.scala 106:25]
  wire  ACEMSHR_reset; // @[ACEUnit.scala 106:25]
  wire  ACEMSHR_write_ready; // @[ACEUnit.scala 106:25]
  wire  ACEMSHR_write_data_valid; // @[ACEUnit.scala 106:25]
  wire [31:0] ACEMSHR_write_data_address; // @[ACEUnit.scala 106:25]
  wire [31:0] ACEMSHR_write_data_core_instruction; // @[ACEUnit.scala 106:25]
  wire [3:0] ACEMSHR_write_data_core_robAddr; // @[ACEUnit.scala 106:25]
  wire [5:0] ACEMSHR_write_data_core_prfDest; // @[ACEUnit.scala 106:25]
  wire  ACEMSHR_write_data_branch_valid; // @[ACEUnit.scala 106:25]
  wire [4:0] ACEMSHR_write_data_branch_mask; // @[ACEUnit.scala 106:25]
  wire  ACEMSHR_write_data_writeData_valid; // @[ACEUnit.scala 106:25]
  wire [63:0] ACEMSHR_write_data_writeData_data; // @[ACEUnit.scala 106:25]
  wire [1:0] ACEMSHR_write_data_cacheLine_response; // @[ACEUnit.scala 106:25]
  wire  ACEMSHR_read_ready; // @[ACEUnit.scala 106:25]
  wire  ACEMSHR_read_data_valid; // @[ACEUnit.scala 106:25]
  wire [31:0] ACEMSHR_read_data_address; // @[ACEUnit.scala 106:25]
  wire [31:0] ACEMSHR_read_data_core_instruction; // @[ACEUnit.scala 106:25]
  wire [3:0] ACEMSHR_read_data_core_robAddr; // @[ACEUnit.scala 106:25]
  wire [5:0] ACEMSHR_read_data_core_prfDest; // @[ACEUnit.scala 106:25]
  wire  ACEMSHR_read_data_branch_valid; // @[ACEUnit.scala 106:25]
  wire [4:0] ACEMSHR_read_data_branch_mask; // @[ACEUnit.scala 106:25]
  wire  ACEMSHR_read_data_writeData_valid; // @[ACEUnit.scala 106:25]
  wire [63:0] ACEMSHR_read_data_writeData_data; // @[ACEUnit.scala 106:25]
  wire [1:0] ACEMSHR_read_data_cacheLine_response; // @[ACEUnit.scala 106:25]
  wire  ACEMSHR_isEmpty; // @[ACEUnit.scala 106:25]
  wire  ACEMSHR_branchOps_valid; // @[ACEUnit.scala 106:25]
  wire [4:0] ACEMSHR_branchOps_branchMask; // @[ACEUnit.scala 106:25]
  wire  ACEMSHR_branchOps_passed; // @[ACEUnit.scala 106:25]
  wire  writeCounter_clock; // @[ACEUnit.scala 170:28]
  wire  writeCounter_reset; // @[ACEUnit.scala 170:28]
  wire [2:0] writeCounter_count; // @[ACEUnit.scala 170:28]
  wire  writeCounter_incrm; // @[ACEUnit.scala 170:28]
  wire  readCounter_clock; // @[ACEUnit.scala 265:27]
  wire  readCounter_reset; // @[ACEUnit.scala 265:27]
  wire [2:0] readCounter_count; // @[ACEUnit.scala 265:27]
  wire  readCounter_incrm; // @[ACEUnit.scala 265:27]
  wire  coherentCounter_clock; // @[ACEUnit.scala 327:31]
  wire  coherentCounter_reset; // @[ACEUnit.scala 327:31]
  wire [2:0] coherentCounter_count; // @[ACEUnit.scala 327:31]
  wire  coherentCounter_incrm; // @[ACEUnit.scala 327:31]
  reg  readBuffer_valid; // @[ACEUnit.scala 104:28]
  reg [31:0] readBuffer_address; // @[ACEUnit.scala 104:28]
  reg [31:0] readBuffer_core_instruction; // @[ACEUnit.scala 104:28]
  reg [3:0] readBuffer_core_robAddr; // @[ACEUnit.scala 104:28]
  reg [5:0] readBuffer_core_prfDest; // @[ACEUnit.scala 104:28]
  reg  readBuffer_branch_valid; // @[ACEUnit.scala 104:28]
  reg [4:0] readBuffer_branch_mask; // @[ACEUnit.scala 104:28]
  reg  readBuffer_writeData_valid; // @[ACEUnit.scala 104:28]
  reg [63:0] readBuffer_writeData_data; // @[ACEUnit.scala 104:28]
  reg [1:0] readBuffer_cacheLine_response; // @[ACEUnit.scala 104:28]
  reg  responseBuffer_valid; // @[ACEUnit.scala 105:31]
  reg [31:0] responseBuffer_address; // @[ACEUnit.scala 105:31]
  reg [31:0] responseBuffer_core_instruction; // @[ACEUnit.scala 105:31]
  reg [3:0] responseBuffer_core_robAddr; // @[ACEUnit.scala 105:31]
  reg [5:0] responseBuffer_core_prfDest; // @[ACEUnit.scala 105:31]
  reg  responseBuffer_branch_valid; // @[ACEUnit.scala 105:31]
  reg [4:0] responseBuffer_branch_mask; // @[ACEUnit.scala 105:31]
  reg  responseBuffer_writeData_valid; // @[ACEUnit.scala 105:31]
  reg [63:0] responseBuffer_writeData_data; // @[ACEUnit.scala 105:31]
  reg [511:0] responseBuffer_cacheLine_cacheLine; // @[ACEUnit.scala 105:31]
  reg [1:0] responseBuffer_cacheLine_response; // @[ACEUnit.scala 105:31]
  reg  writeBuffer_valid; // @[ACEUnit.scala 111:28]
  reg [31:0] writeBuffer_address; // @[ACEUnit.scala 111:28]
  reg [511:0] writeBuffer_data; // @[ACEUnit.scala 111:28]
  reg  coherencyRequestBuffer_valid; // @[ACEUnit.scala 112:39]
  reg [31:0] coherencyRequestBuffer_address; // @[ACEUnit.scala 112:39]
  reg [1:0] coherencyRequestBuffer_response; // @[ACEUnit.scala 112:39]
  reg  coherencyResponseBuffer_valid; // @[ACEUnit.scala 113:40]
  reg [1:0] coherencyResponseBuffer_response; // @[ACEUnit.scala 113:40]
  reg [511:0] coherencyResponseBuffer_cacheLine; // @[ACEUnit.scala 113:40]
  reg  coherencyResponseBuffer_dataValid; // @[ACEUnit.scala 113:40]
  wire  isCoherencyAddressMatchWire = responseBuffer_address[31:6] == coherencyRequestBuffer_address[31:6]; // @[ACEUnit.scala 119:107]
  wire  _T = ~writeBuffer_valid; // @[ACEUnit.scala 121:38]
  wire  _T_1 = writeRequest_request_valid & ~writeBuffer_valid; // @[ACEUnit.scala 121:35]
  wire  _GEN_0 = writeBuffer_valid & writeBuffer_address[31:6] == coherencyRequestBuffer_address[31:6]; // @[ACEUnit.scala 123:33 124:30]
  wire  isWriteAddressMatchWire = writeRequest_request_valid & ~writeBuffer_valid ? writeRequest_request_address[31:6]
     == coherencyRequestBuffer_address[31:6] : _GEN_0; // @[ACEUnit.scala 121:57 122:29]
  wire  _readRequest_ready_T = ~readBuffer_valid; // @[ACEUnit.scala 128:24]
  wire [4:0] _T_4 = readRequest_request_branch_mask & branchOps_branchMask; // @[utils.scala 62:31]
  wire  _T_5 = |_T_4; // @[utils.scala 62:55]
  wire [4:0] _readBuffer_branch_mask_T = readRequest_request_branch_mask ^ branchOps_branchMask; // @[utils.scala 63:42]
  wire [4:0] _GEN_2 = |_T_4 ? _readBuffer_branch_mask_T : readRequest_request_branch_mask; // @[utils.scala 62:60 63:23 65:23]
  wire  _GEN_3 = _T_5 ? 1'h0 : readRequest_request_branch_valid; // @[utils.scala 70:60 71:24 74:24]
  wire [4:0] _GEN_4 = _T_5 ? 5'h0 : readRequest_request_branch_mask; // @[utils.scala 70:60 72:23 75:23]
  wire [4:0] _GEN_5 = branchOps_passed ? _GEN_2 : _GEN_4; // @[utils.scala 60:30]
  wire  _GEN_6 = branchOps_passed ? readRequest_request_branch_valid : _GEN_3; // @[utils.scala 60:30 67:22]
  wire [4:0] _GEN_7 = branchOps_valid ? _GEN_5 : readRequest_request_branch_mask; // @[utils.scala 59:26 80:21]
  wire  _GEN_8 = branchOps_valid ? _GEN_6 : readRequest_request_branch_valid; // @[utils.scala 59:26 79:22]
  wire  _GEN_9 = readRequest_request_valid & readRequest_request_branch_valid & readRequest_ready ?
    readRequest_request_valid : readBuffer_valid; // @[ACEUnit.scala 129:91 130:16 104:28]
  wire  _GEN_14 = readRequest_request_valid & readRequest_request_branch_valid & readRequest_ready ? _GEN_8 :
    readBuffer_branch_valid; // @[ACEUnit.scala 104:28 129:91]
  wire [4:0] _GEN_15 = readRequest_request_valid & readRequest_request_branch_valid & readRequest_ready ? _GEN_7 :
    readBuffer_branch_mask; // @[ACEUnit.scala 104:28 129:91]
  wire [4:0] _T_8 = readBuffer_branch_mask & branchOps_branchMask; // @[utils.scala 122:29]
  wire  _T_9 = |_T_8; // @[utils.scala 122:53]
  wire [4:0] _readBuffer_branch_mask_T_1 = readBuffer_branch_mask ^ branchOps_branchMask; // @[utils.scala 123:40]
  wire [4:0] _GEN_21 = |_T_8 ? _readBuffer_branch_mask_T_1 : _GEN_15; // @[utils.scala 122:58 123:25]
  wire  _GEN_22 = _T_9 ? 1'h0 : _GEN_14; // @[utils.scala 127:58 128:26]
  wire [4:0] _GEN_23 = _T_9 ? 5'h0 : _GEN_15; // @[utils.scala 127:58 129:25]
  wire [4:0] _GEN_24 = branchOps_passed ? _GEN_21 : _GEN_23; // @[utils.scala 121:32]
  wire  _GEN_25 = branchOps_passed ? readBuffer_branch_valid : _GEN_22; // @[utils.scala 121:32 125:24]
  wire [4:0] _T_12 = responseBuffer_branch_mask & branchOps_branchMask; // @[utils.scala 92:27]
  wire  _T_13 = |_T_12; // @[utils.scala 92:51]
  wire [4:0] _readResponse_request_branch_mask_T = responseBuffer_branch_mask ^ branchOps_branchMask; // @[utils.scala 93:42]
  wire [4:0] _GEN_32 = |_T_12 ? _readResponse_request_branch_mask_T : responseBuffer_branch_mask; // @[utils.scala 92:56 93:27 96:27]
  wire [4:0] _GEN_33 = _T_13 ? 5'h0 : responseBuffer_branch_mask; // @[utils.scala 101:56 102:27 106:27]
  wire  _GEN_34 = _T_13 ? 1'h0 : responseBuffer_branch_valid; // @[utils.scala 101:56 103:28 107:28]
  wire [4:0] _GEN_35 = branchOps_passed ? _GEN_32 : _GEN_33; // @[utils.scala 90:30]
  wire  _GEN_36 = branchOps_passed ? responseBuffer_branch_valid : _GEN_34; // @[utils.scala 90:30 98:26]
  wire  _GEN_39 = _T & writeRequest_request_valid ? writeRequest_request_valid : writeBuffer_valid; // @[ACEUnit.scala 147:57 148:17 111:28]
  wire  _coherencyResponse_ready_T = ~coherencyResponseBuffer_valid; // @[ACEUnit.scala 155:30]
  wire  isWireACEBusy = _T_1 | writeBuffer_valid; // @[ACEUnit.scala 173:69]
  reg [1:0] writeACEState; // @[ACEUnit.scala 169:30]
  wire [31:0] _bus_AWADDR_T_1 = {writeBuffer_address[31:6],6'h0}; // @[Cat.scala 33:92]
  wire [63:0] writeChunks__0 = writeBuffer_data[63:0]; // @[ACEUnit.scala 205:25]
  wire [63:0] writeChunks__1 = writeBuffer_data[127:64]; // @[ACEUnit.scala 205:25]
  wire [63:0] writeChunks__2 = writeBuffer_data[191:128]; // @[ACEUnit.scala 205:25]
  wire [63:0] writeChunks__3 = writeBuffer_data[255:192]; // @[ACEUnit.scala 205:25]
  wire [63:0] writeChunks__4 = writeBuffer_data[319:256]; // @[ACEUnit.scala 205:25]
  wire [63:0] writeChunks__5 = writeBuffer_data[383:320]; // @[ACEUnit.scala 205:25]
  wire [63:0] writeChunks__6 = writeBuffer_data[447:384]; // @[ACEUnit.scala 205:25]
  wire [63:0] writeChunks__7 = writeBuffer_data[511:448]; // @[ACEUnit.scala 205:25]
  wire [63:0] _GEN_53 = 3'h1 == writeCounter_count ? writeChunks__1 : writeChunks__0; // @[ACEUnit.scala 210:{17,17}]
  wire [63:0] _GEN_54 = 3'h2 == writeCounter_count ? writeChunks__2 : _GEN_53; // @[ACEUnit.scala 210:{17,17}]
  wire [63:0] _GEN_55 = 3'h3 == writeCounter_count ? writeChunks__3 : _GEN_54; // @[ACEUnit.scala 210:{17,17}]
  wire [63:0] _GEN_56 = 3'h4 == writeCounter_count ? writeChunks__4 : _GEN_55; // @[ACEUnit.scala 210:{17,17}]
  wire [63:0] _GEN_57 = 3'h5 == writeCounter_count ? writeChunks__5 : _GEN_56; // @[ACEUnit.scala 210:{17,17}]
  wire [63:0] _GEN_58 = 3'h6 == writeCounter_count ? writeChunks__6 : _GEN_57; // @[ACEUnit.scala 210:{17,17}]
  wire [63:0] _GEN_59 = 3'h7 == writeCounter_count ? writeChunks__7 : _GEN_58; // @[ACEUnit.scala 210:{17,17}]
  wire [1:0] _writeACEState_T_3 = bus_WLAST & bus_WREADY ? 2'h3 : 2'h2; // @[ACEUnit.scala 211:27]
  wire  _writeBuffer_valid_T_2 = bus_BRESP == 2'h0; // @[ACEUnit.scala 215:74]
  wire [1:0] _writeACEState_T_7 = _writeBuffer_valid_T_2 ? 2'h0 : 2'h1; // @[ACEUnit.scala 218:28]
  wire [1:0] _writeACEState_T_8 = bus_BVALID ? _writeACEState_T_7 : 2'h3; // @[ACEUnit.scala 217:27]
  wire  _GEN_61 = 2'h3 == writeACEState ? ~(bus_BVALID & bus_BRESP == 2'h0) : _GEN_39; // @[ACEUnit.scala 174:25 215:25]
  wire [1:0] _GEN_62 = 2'h3 == writeACEState ? _writeACEState_T_8 : writeACEState; // @[ACEUnit.scala 174:25 217:21 169:30]
  wire  _GEN_65 = 2'h2 == writeACEState & writeCounter_count == 3'h7; // @[ACEUnit.scala 174:25 201:17 68:13]
  wire [63:0] _GEN_67 = 2'h2 == writeACEState ? _GEN_59 : 64'h0; // @[ACEUnit.scala 174:25 210:17 66:13]
  wire  _GEN_69 = 2'h2 == writeACEState ? 1'h0 : 2'h3 == writeACEState; // @[ACEUnit.scala 174:25 71:14]
  wire [31:0] _GEN_73 = 2'h1 == writeACEState ? _bus_AWADDR_T_1 : 32'h0; // @[ACEUnit.scala 174:25 183:18 56:14]
  wire [1:0] _GEN_75 = 2'h1 == writeACEState ? 2'h3 : 2'h0; // @[ACEUnit.scala 174:25 185:18 58:14]
  wire  _GEN_79 = 2'h1 == writeACEState ? 1'h0 : 2'h2 == writeACEState; // @[ACEUnit.scala 174:25 69:14]
  wire  _GEN_81 = 2'h1 == writeACEState ? 1'h0 : _GEN_65; // @[ACEUnit.scala 174:25 68:13]
  wire  _GEN_82 = 2'h1 == writeACEState ? 1'h0 : 2'h2 == writeACEState & bus_WREADY; // @[ACEUnit.scala 171:22 174:25]
  wire [63:0] _GEN_83 = 2'h1 == writeACEState ? 64'h0 : _GEN_67; // @[ACEUnit.scala 174:25 66:13]
  wire  _GEN_84 = 2'h1 == writeACEState ? 1'h0 : _GEN_69; // @[ACEUnit.scala 174:25 71:14]
  wire [1:0] _GEN_92 = 2'h0 == writeACEState ? 2'h0 : _GEN_75; // @[ACEUnit.scala 174:25 58:14]
  reg  readACERequestState; // @[ACEUnit.scala 224:36]
  reg [1:0] coherentAXIState; // @[ACEUnit.scala 326:33]
  wire  isCoherencyIdle = coherentAXIState == 2'h0; // @[ACEUnit.scala 329:40]
  wire [31:0] _bus_ARADDR_T_1 = {readBuffer_address[31:6],6'h0}; // @[Cat.scala 33:92]
  wire [3:0] _GEN_102 = 2'h3 == readBuffer_cacheLine_response ? 4'hb : 4'h1; // @[ACEUnit.scala 242:19 243:49 246:34]
  wire [3:0] _GEN_103 = 2'h1 == readBuffer_cacheLine_response ? 4'h7 : _GEN_102; // @[ACEUnit.scala 243:49 245:34]
  wire [3:0] _GEN_104 = 2'h0 == readBuffer_cacheLine_response ? 4'h1 : _GEN_103; // @[ACEUnit.scala 243:49 244:34]
  wire [4:0] _GEN_105 = _T_9 ? _readBuffer_branch_mask_T_1 : readBuffer_branch_mask; // @[utils.scala 92:56 93:27 96:27]
  wire [4:0] _GEN_106 = _T_9 ? 5'h0 : readBuffer_branch_mask; // @[utils.scala 101:56 102:27 106:27]
  wire  _GEN_107 = _T_9 ? 1'h0 : readBuffer_branch_valid; // @[utils.scala 101:56 103:28 107:28]
  wire [4:0] _GEN_108 = branchOps_passed ? _GEN_105 : _GEN_106; // @[utils.scala 90:30]
  wire  _GEN_109 = branchOps_passed ? readBuffer_branch_valid : _GEN_107; // @[utils.scala 90:30 98:26]
  wire [4:0] _GEN_110 = branchOps_valid ? _GEN_108 : readBuffer_branch_mask; // @[utils.scala 111:23 89:27]
  wire  _GEN_111 = branchOps_valid ? _GEN_109 : readBuffer_branch_valid; // @[utils.scala 112:24 89:27]
  wire [1:0] _GEN_113 = bus_ARREADY ? readBuffer_cacheLine_response : 2'h0; // @[ACEUnit.scala 251:24 252:28 utils.scala 49:41]
  wire [63:0] _GEN_115 = bus_ARREADY ? readBuffer_writeData_data : 64'h0; // @[ACEUnit.scala 251:24 252:28 utils.scala 49:41]
  wire  _GEN_116 = bus_ARREADY & readBuffer_writeData_valid; // @[ACEUnit.scala 251:24 252:28 utils.scala 48:41]
  wire [4:0] _GEN_117 = bus_ARREADY ? _GEN_110 : 5'h0; // @[ACEUnit.scala 251:24 utils.scala 49:41]
  wire  _GEN_118 = bus_ARREADY & _GEN_111; // @[ACEUnit.scala 251:24 utils.scala 48:41]
  wire [5:0] _GEN_119 = bus_ARREADY ? readBuffer_core_prfDest : 6'h0; // @[ACEUnit.scala 251:24 252:28 utils.scala 49:41]
  wire [3:0] _GEN_120 = bus_ARREADY ? readBuffer_core_robAddr : 4'h0; // @[ACEUnit.scala 251:24 252:28 utils.scala 49:41]
  wire [31:0] _GEN_121 = bus_ARREADY ? readBuffer_core_instruction : 32'h0; // @[ACEUnit.scala 251:24 252:28 utils.scala 49:41]
  wire [31:0] _GEN_122 = bus_ARREADY ? readBuffer_address : 32'h0; // @[ACEUnit.scala 251:24 252:28 utils.scala 49:41]
  wire  _GEN_123 = bus_ARREADY & readBuffer_valid; // @[ACEUnit.scala 251:24 252:28 utils.scala 48:41]
  wire [31:0] _GEN_127 = readACERequestState ? _bus_ARADDR_T_1 : 32'h0; // @[ACEUnit.scala 225:31 232:18 74:14]
  wire [3:0] _GEN_132 = readACERequestState ? _GEN_104 : 4'h0; // @[ACEUnit.scala 225:31 92:15]
  wire [1:0] _GEN_134 = readACERequestState ? _GEN_113 : 2'h0; // @[ACEUnit.scala 225:31 utils.scala 49:41]
  wire [63:0] _GEN_136 = readACERequestState ? _GEN_115 : 64'h0; // @[ACEUnit.scala 225:31 utils.scala 49:41]
  wire [4:0] _GEN_138 = readACERequestState ? _GEN_117 : 5'h0; // @[ACEUnit.scala 225:31 utils.scala 49:41]
  wire [5:0] _GEN_140 = readACERequestState ? _GEN_119 : 6'h0; // @[ACEUnit.scala 225:31 utils.scala 49:41]
  wire [3:0] _GEN_141 = readACERequestState ? _GEN_120 : 4'h0; // @[ACEUnit.scala 225:31 utils.scala 49:41]
  wire [31:0] _GEN_142 = readACERequestState ? _GEN_121 : 32'h0; // @[ACEUnit.scala 225:31 utils.scala 49:41]
  wire [31:0] _GEN_143 = readACERequestState ? _GEN_122 : 32'h0; // @[ACEUnit.scala 225:31 utils.scala 49:41]
  reg [1:0] readACEResponseState; // @[ACEUnit.scala 261:37]
  reg [63:0] readDataVec_0; // @[ACEUnit.scala 262:28]
  reg [63:0] readDataVec_1; // @[ACEUnit.scala 262:28]
  reg [63:0] readDataVec_2; // @[ACEUnit.scala 262:28]
  reg [63:0] readDataVec_3; // @[ACEUnit.scala 262:28]
  reg [63:0] readDataVec_4; // @[ACEUnit.scala 262:28]
  reg [63:0] readDataVec_5; // @[ACEUnit.scala 262:28]
  reg [63:0] readDataVec_6; // @[ACEUnit.scala 262:28]
  reg [63:0] readDataVec_7; // @[ACEUnit.scala 262:28]
  reg  readResponseValid; // @[ACEUnit.scala 263:34]
  reg [1:0] readResponseReg; // @[ACEUnit.scala 264:32]
  wire  _T_34 = ~ACEMSHR_isEmpty; // @[ACEUnit.scala 272:12]
  wire  _GEN_175 = ~ACEMSHR_isEmpty ? ACEMSHR_read_data_branch_valid : responseBuffer_branch_valid; // @[ACEUnit.scala 272:29 274:24 105:31]
  wire [4:0] _GEN_176 = ~ACEMSHR_isEmpty ? ACEMSHR_read_data_branch_mask : responseBuffer_branch_mask; // @[ACEUnit.scala 272:29 274:24 105:31]
  wire  isCleanUniqueWire = responseBuffer_cacheLine_response == 2'h3; // @[ACEUnit.scala 281:65]
  wire  _readResponseValid_T_2 = bus_RRESP[1:0] == 2'h0 & readResponseValid; // @[ACEUnit.scala 286:33]
  wire [63:0] _GEN_182 = 3'h0 == readCounter_count ? bus_RDATA : readDataVec_0; // @[ACEUnit.scala 262:28 291:{42,42}]
  wire [63:0] _GEN_183 = 3'h1 == readCounter_count ? bus_RDATA : readDataVec_1; // @[ACEUnit.scala 262:28 291:{42,42}]
  wire [63:0] _GEN_184 = 3'h2 == readCounter_count ? bus_RDATA : readDataVec_2; // @[ACEUnit.scala 262:28 291:{42,42}]
  wire [63:0] _GEN_185 = 3'h3 == readCounter_count ? bus_RDATA : readDataVec_3; // @[ACEUnit.scala 262:28 291:{42,42}]
  wire [63:0] _GEN_186 = 3'h4 == readCounter_count ? bus_RDATA : readDataVec_4; // @[ACEUnit.scala 262:28 291:{42,42}]
  wire [63:0] _GEN_187 = 3'h5 == readCounter_count ? bus_RDATA : readDataVec_5; // @[ACEUnit.scala 262:28 291:{42,42}]
  wire [63:0] _GEN_188 = 3'h6 == readCounter_count ? bus_RDATA : readDataVec_6; // @[ACEUnit.scala 262:28 291:{42,42}]
  wire [63:0] _GEN_189 = 3'h7 == readCounter_count ? bus_RDATA : readDataVec_7; // @[ACEUnit.scala 262:28 291:{42,42}]
  wire [63:0] _GEN_191 = bus_RVALID ? _GEN_182 : readDataVec_0; // @[ACEUnit.scala 262:28 289:45]
  wire [63:0] _GEN_192 = bus_RVALID ? _GEN_183 : readDataVec_1; // @[ACEUnit.scala 262:28 289:45]
  wire [63:0] _GEN_193 = bus_RVALID ? _GEN_184 : readDataVec_2; // @[ACEUnit.scala 262:28 289:45]
  wire [63:0] _GEN_194 = bus_RVALID ? _GEN_185 : readDataVec_3; // @[ACEUnit.scala 262:28 289:45]
  wire [63:0] _GEN_195 = bus_RVALID ? _GEN_186 : readDataVec_4; // @[ACEUnit.scala 262:28 289:45]
  wire [63:0] _GEN_196 = bus_RVALID ? _GEN_187 : readDataVec_5; // @[ACEUnit.scala 262:28 289:45]
  wire [63:0] _GEN_197 = bus_RVALID ? _GEN_188 : readDataVec_6; // @[ACEUnit.scala 262:28 289:45]
  wire [63:0] _GEN_198 = bus_RVALID ? _GEN_189 : readDataVec_7; // @[ACEUnit.scala 262:28 289:45]
  wire  _GEN_199 = bus_RVALID ? _readResponseValid_T_2 : readResponseValid; // @[ACEUnit.scala 289:45 292:29 263:34]
  wire [1:0] _GEN_200 = bus_RVALID ? bus_RRESP[3:2] : readResponseReg; // @[ACEUnit.scala 289:45 293:27 264:32]
  wire  _GEN_202 = isCleanUniqueWire ? bus_RRESP[1:0] == 2'h0 & readResponseValid : _GEN_199; // @[ACEUnit.scala 284:30 286:27]
  wire  _GEN_203 = isCleanUniqueWire | (readCounter_count != 3'h0 | bus_RVALID & readCounter_count == 3'h0); // @[ACEUnit.scala 284:30 287:24 295:24]
  wire  _GEN_204 = isCleanUniqueWire ? 1'h0 : bus_RVALID; // @[ACEUnit.scala 266:21 284:30]
  wire [1:0] _readACEResponseState_T_5 = bus_RVALID ? 2'h2 : 2'h1; // @[ACEUnit.scala 300:36]
  wire [1:0] _readACEResponseState_T_8 = bus_RLAST & bus_RVALID & readResponseValid ? 2'h2 : 2'h1; // @[ACEUnit.scala 302:36]
  wire [511:0] _responseBuffer_cacheLine_cacheLine_T = {readDataVec_7,readDataVec_6,readDataVec_5,readDataVec_4,
    readDataVec_3,readDataVec_2,readDataVec_1,readDataVec_0}; // @[Cat.scala 33:92]
  wire  _GEN_214 = responseBuffer_valid & readResponse_ready ? 1'h0 : 1'h1; // @[ACEUnit.scala 306:28 310:55 311:30]
  wire [1:0] _readACEResponseState_T_9 = readResponse_ready ? 2'h0 : 2'h2; // @[ACEUnit.scala 316:34]
  wire  _GEN_222 = 2'h1 == readACEResponseState ? _GEN_202 : readResponseValid; // @[ACEUnit.scala 268:32 263:34]
  wire  _GEN_223 = 2'h1 == readACEResponseState ? _GEN_203 : 2'h2 == readACEResponseState; // @[ACEUnit.scala 268:32]
  wire  _GEN_244 = 2'h0 == readACEResponseState ? _GEN_175 : responseBuffer_branch_valid; // @[ACEUnit.scala 105:31 268:32]
  wire [4:0] _GEN_245 = 2'h0 == readACEResponseState ? _GEN_176 : responseBuffer_branch_mask; // @[ACEUnit.scala 105:31 268:32]
  wire  _GEN_254 = 2'h0 == readACEResponseState ? readResponseValid : _GEN_222; // @[ACEUnit.scala 268:32 263:34]
  wire  isReadRespBusy = 2'h0 == readACEResponseState ? 1'h0 : _GEN_223; // @[ACEUnit.scala 268:32]
  wire [4:0] _GEN_265 = _T_13 ? _readResponse_request_branch_mask_T : _GEN_245; // @[utils.scala 122:58 123:25]
  wire  _GEN_266 = _T_13 ? 1'h0 : _GEN_244; // @[utils.scala 127:58 128:26]
  wire [4:0] _GEN_267 = _T_13 ? 5'h0 : _GEN_245; // @[utils.scala 127:58 129:25]
  reg  coherentRequestSend; // @[ACEUnit.scala 328:36]
  wire  _coherencyRequestBuffer_response_T_1 = bus_ACSNOOP == 4'h7; // @[ACEUnit.scala 341:91]
  wire  _coherencyRequestBuffer_response_T_2 = bus_ACSNOOP == 4'h9 | bus_ACSNOOP == 4'h7; // @[ACEUnit.scala 341:75]
  wire  _coherencyRequestBuffer_response_T_5 = bus_ACSNOOP == 4'h1 | _coherencyRequestBuffer_response_T_1; // @[ACEUnit.scala 342:76]
  wire [1:0] _coherencyRequestBuffer_response_T_6 = {_coherencyRequestBuffer_response_T_2,
    _coherencyRequestBuffer_response_T_5}; // @[Cat.scala 33:92]
  wire  _coherencyRequestBuffer_valid_T = coherencyRequest_ready ? 1'h0 : 1'h1; // @[ACEUnit.scala 348:43]
  wire  _coherencyRequestBuffer_valid_T_2 = isReadRespBusy & isCoherencyAddressMatchWire ? 1'h0 : 1'h1; // @[ACEUnit.scala 351:46]
  wire  _GEN_274 = ~coherentRequestSend ? _coherencyRequestBuffer_valid_T_2 : coherencyRequestBuffer_valid; // @[ACEUnit.scala 350:35 112:39 351:40]
  wire  _GEN_275 = ~coherentRequestSend ? _coherencyRequestBuffer_valid_T_2 : coherentRequestSend; // @[ACEUnit.scala 350:35 352:31 328:36]
  wire [1:0] _coherentAXIState_T_1 = writeBuffer_valid ? 2'h2 : 2'h1; // @[ACEUnit.scala 357:32]
  wire [1:0] _coherentAXIState_T_2 = coherencyResponse_request_valid ? 2'h2 : 2'h1; // @[ACEUnit.scala 359:32]
  wire [4:0] _bus_CRRESP_T_2 = {1'h0,coherencyResponseBuffer_response[1],coherencyResponseBuffer_response[0],1'h0,
    coherencyResponseBuffer_dataValid}; // @[Cat.scala 33:92]
  wire [4:0] _bus_CRRESP_T_3 = coherencyResponseBuffer_valid ? _bus_CRRESP_T_2 : 5'h0; // @[ACEUnit.scala 368:24]
  wire [1:0] _coherentAXIState_T_3 = coherencyResponseBuffer_dataValid ? 2'h3 : 2'h0; // @[ACEUnit.scala 371:32]
  wire [1:0] _GEN_279 = bus_CRREADY ? _coherentAXIState_T_3 : 2'h2; // @[ACEUnit.scala 370:24 371:26 373:26]
  wire [63:0] writeChunks_1_0 = coherencyResponseBuffer_cacheLine[63:0]; // @[ACEUnit.scala 381:42]
  wire [63:0] writeChunks_1_1 = coherencyResponseBuffer_cacheLine[127:64]; // @[ACEUnit.scala 381:42]
  wire [63:0] writeChunks_1_2 = coherencyResponseBuffer_cacheLine[191:128]; // @[ACEUnit.scala 381:42]
  wire [63:0] writeChunks_1_3 = coherencyResponseBuffer_cacheLine[255:192]; // @[ACEUnit.scala 381:42]
  wire [63:0] writeChunks_1_4 = coherencyResponseBuffer_cacheLine[319:256]; // @[ACEUnit.scala 381:42]
  wire [63:0] writeChunks_1_5 = coherencyResponseBuffer_cacheLine[383:320]; // @[ACEUnit.scala 381:42]
  wire [63:0] writeChunks_1_6 = coherencyResponseBuffer_cacheLine[447:384]; // @[ACEUnit.scala 381:42]
  wire [63:0] writeChunks_1_7 = coherencyResponseBuffer_cacheLine[511:448]; // @[ACEUnit.scala 381:42]
  wire [63:0] _GEN_282 = 3'h1 == coherentCounter_count ? writeChunks_1_1 : writeChunks_1_0; // @[ACEUnit.scala 386:{18,18}]
  wire [63:0] _GEN_283 = 3'h2 == coherentCounter_count ? writeChunks_1_2 : _GEN_282; // @[ACEUnit.scala 386:{18,18}]
  wire [63:0] _GEN_284 = 3'h3 == coherentCounter_count ? writeChunks_1_3 : _GEN_283; // @[ACEUnit.scala 386:{18,18}]
  wire [63:0] _GEN_285 = 3'h4 == coherentCounter_count ? writeChunks_1_4 : _GEN_284; // @[ACEUnit.scala 386:{18,18}]
  wire [63:0] _GEN_286 = 3'h5 == coherentCounter_count ? writeChunks_1_5 : _GEN_285; // @[ACEUnit.scala 386:{18,18}]
  wire [63:0] _GEN_287 = 3'h6 == coherentCounter_count ? writeChunks_1_6 : _GEN_286; // @[ACEUnit.scala 386:{18,18}]
  wire [63:0] _GEN_288 = 3'h7 == coherentCounter_count ? writeChunks_1_7 : _GEN_287; // @[ACEUnit.scala 386:{18,18}]
  wire [1:0] _coherentAXIState_T_5 = bus_CDLAST & bus_CDREADY ? 2'h0 : 2'h3; // @[ACEUnit.scala 389:30]
  wire [63:0] _GEN_291 = 2'h3 == coherentAXIState ? _GEN_288 : 64'h0; // @[ACEUnit.scala 101:14 332:27 386:18]
  wire  _GEN_292 = 2'h3 == coherentAXIState & coherentCounter_count == 3'h7; // @[ACEUnit.scala 102:14 332:27 387:18]
  wire [1:0] _GEN_293 = 2'h3 == coherentAXIState ? _coherentAXIState_T_5 : coherentAXIState; // @[ACEUnit.scala 332:27 389:24 326:33]
  wire [4:0] _GEN_296 = 2'h2 == coherentAXIState ? _bus_CRRESP_T_3 : 5'h0; // @[ACEUnit.scala 332:27 368:18 98:14]
  wire  _GEN_298 = 2'h2 == coherentAXIState ? 1'h0 : 2'h3 == coherentAXIState; // @[ACEUnit.scala 100:15 332:27]
  wire  _GEN_299 = 2'h2 == coherentAXIState ? 1'h0 : 2'h3 == coherentAXIState & bus_CDREADY; // @[ACEUnit.scala 330:25 332:27]
  wire [63:0] _GEN_300 = 2'h2 == coherentAXIState ? 64'h0 : _GEN_291; // @[ACEUnit.scala 101:14 332:27]
  wire  _GEN_301 = 2'h2 == coherentAXIState ? 1'h0 : _GEN_292; // @[ACEUnit.scala 102:14 332:27]
  wire  _GEN_305 = 2'h1 == coherentAXIState ? 1'h0 : 2'h2 == coherentAXIState; // @[ACEUnit.scala 332:27 97:15]
  wire [4:0] _GEN_306 = 2'h1 == coherentAXIState ? 5'h0 : _GEN_296; // @[ACEUnit.scala 332:27 98:14]
  wire  _GEN_307 = 2'h1 == coherentAXIState ? 1'h0 : _GEN_298; // @[ACEUnit.scala 100:15 332:27]
  wire  _GEN_308 = 2'h1 == coherentAXIState ? 1'h0 : _GEN_299; // @[ACEUnit.scala 330:25 332:27]
  wire [63:0] _GEN_309 = 2'h1 == coherentAXIState ? 64'h0 : _GEN_300; // @[ACEUnit.scala 101:14 332:27]
  wire  _GEN_310 = 2'h1 == coherentAXIState ? 1'h0 : _GEN_301; // @[ACEUnit.scala 102:14 332:27]
  fifoWithBranchOps ACEMSHR ( // @[ACEUnit.scala 106:25]
    .clock(ACEMSHR_clock),
    .reset(ACEMSHR_reset),
    .write_ready(ACEMSHR_write_ready),
    .write_data_valid(ACEMSHR_write_data_valid),
    .write_data_address(ACEMSHR_write_data_address),
    .write_data_core_instruction(ACEMSHR_write_data_core_instruction),
    .write_data_core_robAddr(ACEMSHR_write_data_core_robAddr),
    .write_data_core_prfDest(ACEMSHR_write_data_core_prfDest),
    .write_data_branch_valid(ACEMSHR_write_data_branch_valid),
    .write_data_branch_mask(ACEMSHR_write_data_branch_mask),
    .write_data_writeData_valid(ACEMSHR_write_data_writeData_valid),
    .write_data_writeData_data(ACEMSHR_write_data_writeData_data),
    .write_data_cacheLine_response(ACEMSHR_write_data_cacheLine_response),
    .read_ready(ACEMSHR_read_ready),
    .read_data_valid(ACEMSHR_read_data_valid),
    .read_data_address(ACEMSHR_read_data_address),
    .read_data_core_instruction(ACEMSHR_read_data_core_instruction),
    .read_data_core_robAddr(ACEMSHR_read_data_core_robAddr),
    .read_data_core_prfDest(ACEMSHR_read_data_core_prfDest),
    .read_data_branch_valid(ACEMSHR_read_data_branch_valid),
    .read_data_branch_mask(ACEMSHR_read_data_branch_mask),
    .read_data_writeData_valid(ACEMSHR_read_data_writeData_valid),
    .read_data_writeData_data(ACEMSHR_read_data_writeData_data),
    .read_data_cacheLine_response(ACEMSHR_read_data_cacheLine_response),
    .isEmpty(ACEMSHR_isEmpty),
    .branchOps_valid(ACEMSHR_branchOps_valid),
    .branchOps_branchMask(ACEMSHR_branchOps_branchMask),
    .branchOps_passed(ACEMSHR_branchOps_passed)
  );
  moduleCounter_2 writeCounter ( // @[ACEUnit.scala 170:28]
    .clock(writeCounter_clock),
    .reset(writeCounter_reset),
    .count(writeCounter_count),
    .incrm(writeCounter_incrm)
  );
  moduleCounter_2 readCounter ( // @[ACEUnit.scala 265:27]
    .clock(readCounter_clock),
    .reset(readCounter_reset),
    .count(readCounter_count),
    .incrm(readCounter_incrm)
  );
  moduleCounter_2 coherentCounter ( // @[ACEUnit.scala 327:31]
    .clock(coherentCounter_clock),
    .reset(coherentCounter_reset),
    .count(coherentCounter_count),
    .incrm(coherentCounter_incrm)
  );
  assign readRequest_ready = ~readBuffer_valid; // @[ACEUnit.scala 128:24]
  assign readResponse_request_valid = responseBuffer_valid; // @[ACEUnit.scala 138:24]
  assign readResponse_request_address = responseBuffer_address; // @[ACEUnit.scala 138:24]
  assign readResponse_request_core_instruction = responseBuffer_core_instruction; // @[ACEUnit.scala 138:24]
  assign readResponse_request_core_robAddr = responseBuffer_core_robAddr; // @[ACEUnit.scala 138:24]
  assign readResponse_request_core_prfDest = responseBuffer_core_prfDest; // @[ACEUnit.scala 138:24]
  assign readResponse_request_branch_valid = branchOps_valid ? _GEN_36 : responseBuffer_branch_valid; // @[utils.scala 112:24 89:27]
  assign readResponse_request_branch_mask = branchOps_valid ? _GEN_35 : responseBuffer_branch_mask; // @[utils.scala 111:23 89:27]
  assign readResponse_request_writeData_valid = responseBuffer_writeData_valid; // @[ACEUnit.scala 138:24]
  assign readResponse_request_writeData_data = responseBuffer_writeData_data; // @[ACEUnit.scala 138:24]
  assign readResponse_request_cacheLine_cacheLine = responseBuffer_cacheLine_cacheLine; // @[ACEUnit.scala 138:24]
  assign readResponse_request_cacheLine_response = responseBuffer_cacheLine_response; // @[ACEUnit.scala 138:24]
  assign writeRequest_ready = ~writeBuffer_valid; // @[ACEUnit.scala 146:25]
  assign coherencyRequest_request_valid = coherencyRequestBuffer_valid; // @[ACEUnit.scala 152:28]
  assign coherencyRequest_request_address = coherencyRequestBuffer_address; // @[ACEUnit.scala 152:28]
  assign coherencyRequest_request_response = coherencyRequestBuffer_response; // @[ACEUnit.scala 152:28]
  assign coherencyResponse_ready = ~coherencyResponseBuffer_valid; // @[ACEUnit.scala 155:30]
  assign fenceReady = _readRequest_ready_T & ~responseBuffer_valid & ACEMSHR_isEmpty; // @[ACEUnit.scala 392:60]
  assign bus_AWADDR = 2'h0 == writeACEState ? 32'h0 : _GEN_73; // @[ACEUnit.scala 174:25 56:14]
  assign bus_AWVALID = 2'h0 == writeACEState ? 1'h0 : 2'h1 == writeACEState; // @[ACEUnit.scala 174:25 64:15]
  assign bus_WDATA = 2'h0 == writeACEState ? 64'h0 : _GEN_83; // @[ACEUnit.scala 174:25 66:13]
  assign bus_WLAST = 2'h0 == writeACEState ? 1'h0 : _GEN_81; // @[ACEUnit.scala 174:25 68:13]
  assign bus_WVALID = 2'h0 == writeACEState ? 1'h0 : _GEN_79; // @[ACEUnit.scala 174:25 69:14]
  assign bus_BREADY = 2'h0 == writeACEState ? 1'h0 : _GEN_84; // @[ACEUnit.scala 174:25 71:14]
  assign bus_ARADDR = ~readACERequestState ? 32'h0 : _GEN_127; // @[ACEUnit.scala 225:31 74:14]
  assign bus_ARVALID = ~readACERequestState ? 1'h0 : readACERequestState; // @[ACEUnit.scala 225:31 82:15]
  assign bus_RREADY = 2'h0 == readACEResponseState ? 1'h0 : 2'h1 == readACEResponseState; // @[ACEUnit.scala 268:32 84:14]
  assign bus_AWSNOOP = {{1'd0}, _GEN_92};
  assign bus_ARSNOOP = ~readACERequestState ? 4'h0 : _GEN_132; // @[ACEUnit.scala 225:31 92:15]
  assign bus_ACREADY = 2'h0 == coherentAXIState; // @[ACEUnit.scala 332:27]
  assign bus_CRVALID = 2'h0 == coherentAXIState ? 1'h0 : _GEN_305; // @[ACEUnit.scala 332:27 97:15]
  assign bus_CRRESP = 2'h0 == coherentAXIState ? 5'h0 : _GEN_306; // @[ACEUnit.scala 332:27 98:14]
  assign bus_CDVALID = 2'h0 == coherentAXIState ? 1'h0 : _GEN_307; // @[ACEUnit.scala 100:15 332:27]
  assign bus_CDDATA = 2'h0 == coherentAXIState ? 64'h0 : _GEN_309; // @[ACEUnit.scala 101:14 332:27]
  assign bus_CDLAST = 2'h0 == coherentAXIState ? 1'h0 : _GEN_310; // @[ACEUnit.scala 102:14 332:27]
  assign ACEMSHR_clock = clock;
  assign ACEMSHR_reset = reset;
  assign ACEMSHR_write_data_valid = ~readACERequestState ? 1'h0 : readACERequestState & _GEN_123; // @[ACEUnit.scala 225:31 utils.scala 48:41]
  assign ACEMSHR_write_data_address = ~readACERequestState ? 32'h0 : _GEN_143; // @[ACEUnit.scala 225:31 utils.scala 49:41]
  assign ACEMSHR_write_data_core_instruction = ~readACERequestState ? 32'h0 : _GEN_142; // @[ACEUnit.scala 225:31 utils.scala 49:41]
  assign ACEMSHR_write_data_core_robAddr = ~readACERequestState ? 4'h0 : _GEN_141; // @[ACEUnit.scala 225:31 utils.scala 49:41]
  assign ACEMSHR_write_data_core_prfDest = ~readACERequestState ? 6'h0 : _GEN_140; // @[ACEUnit.scala 225:31 utils.scala 49:41]
  assign ACEMSHR_write_data_branch_valid = ~readACERequestState ? 1'h0 : readACERequestState & _GEN_118; // @[ACEUnit.scala 225:31 utils.scala 48:41]
  assign ACEMSHR_write_data_branch_mask = ~readACERequestState ? 5'h0 : _GEN_138; // @[ACEUnit.scala 225:31 utils.scala 49:41]
  assign ACEMSHR_write_data_writeData_valid = ~readACERequestState ? 1'h0 : readACERequestState & _GEN_116; // @[ACEUnit.scala 225:31 utils.scala 48:41]
  assign ACEMSHR_write_data_writeData_data = ~readACERequestState ? 64'h0 : _GEN_136; // @[ACEUnit.scala 225:31 utils.scala 49:41]
  assign ACEMSHR_write_data_cacheLine_response = ~readACERequestState ? 2'h0 : _GEN_134; // @[ACEUnit.scala 225:31 utils.scala 49:41]
  assign ACEMSHR_read_ready = 2'h0 == readACEResponseState & _T_34; // @[ACEUnit.scala 142:22 268:32]
  assign ACEMSHR_branchOps_valid = branchOps_valid; // @[ACEUnit.scala 143:21]
  assign ACEMSHR_branchOps_branchMask = branchOps_branchMask; // @[ACEUnit.scala 143:21]
  assign ACEMSHR_branchOps_passed = branchOps_passed; // @[ACEUnit.scala 143:21]
  assign writeCounter_clock = clock;
  assign writeCounter_reset = 2'h0 == writeACEState; // @[ACEUnit.scala 174:25]
  assign writeCounter_incrm = 2'h0 == writeACEState ? 1'h0 : _GEN_82; // @[ACEUnit.scala 171:22 174:25]
  assign readCounter_clock = clock;
  assign readCounter_reset = 2'h0 == readACEResponseState; // @[ACEUnit.scala 268:32]
  assign readCounter_incrm = 2'h0 == readACEResponseState ? 1'h0 : 2'h1 == readACEResponseState & _GEN_204; // @[ACEUnit.scala 266:21 268:32]
  assign coherentCounter_clock = clock;
  assign coherentCounter_reset = 2'h0 == coherentAXIState ? 1'h0 : _GEN_305; // @[ACEUnit.scala 332:27 97:15]
  assign coherentCounter_incrm = 2'h0 == coherentAXIState ? 1'h0 : _GEN_308; // @[ACEUnit.scala 330:25 332:27]
  always @(posedge clock) begin
    if (reset) begin // @[ACEUnit.scala 104:28]
      readBuffer_valid <= 1'h0; // @[ACEUnit.scala 104:28]
    end else if (~readACERequestState) begin // @[ACEUnit.scala 225:31]
      readBuffer_valid <= _GEN_9;
    end else if (readACERequestState) begin // @[ACEUnit.scala 225:31]
      if (bus_ARREADY) begin // @[ACEUnit.scala 251:24]
        readBuffer_valid <= 1'h0; // @[ACEUnit.scala 254:26]
      end else begin
        readBuffer_valid <= _GEN_9;
      end
    end else begin
      readBuffer_valid <= _GEN_9;
    end
    if (reset) begin // @[ACEUnit.scala 104:28]
      readBuffer_address <= 32'h0; // @[ACEUnit.scala 104:28]
    end else if (readRequest_request_valid & readRequest_request_branch_valid & readRequest_ready) begin // @[ACEUnit.scala 129:91]
      readBuffer_address <= readRequest_request_address; // @[ACEUnit.scala 130:16]
    end
    if (reset) begin // @[ACEUnit.scala 104:28]
      readBuffer_core_instruction <= 32'h0; // @[ACEUnit.scala 104:28]
    end else if (readRequest_request_valid & readRequest_request_branch_valid & readRequest_ready) begin // @[ACEUnit.scala 129:91]
      readBuffer_core_instruction <= readRequest_request_core_instruction; // @[ACEUnit.scala 130:16]
    end
    if (reset) begin // @[ACEUnit.scala 104:28]
      readBuffer_core_robAddr <= 4'h0; // @[ACEUnit.scala 104:28]
    end else if (readRequest_request_valid & readRequest_request_branch_valid & readRequest_ready) begin // @[ACEUnit.scala 129:91]
      readBuffer_core_robAddr <= readRequest_request_core_robAddr; // @[ACEUnit.scala 130:16]
    end
    if (reset) begin // @[ACEUnit.scala 104:28]
      readBuffer_core_prfDest <= 6'h0; // @[ACEUnit.scala 104:28]
    end else if (readRequest_request_valid & readRequest_request_branch_valid & readRequest_ready) begin // @[ACEUnit.scala 129:91]
      readBuffer_core_prfDest <= readRequest_request_core_prfDest; // @[ACEUnit.scala 130:16]
    end
    if (reset) begin // @[ACEUnit.scala 104:28]
      readBuffer_branch_valid <= 1'h0; // @[ACEUnit.scala 104:28]
    end else if (readBuffer_valid) begin // @[ACEUnit.scala 133:25]
      if (readBuffer_branch_valid) begin // @[utils.scala 119:24]
        if (branchOps_valid) begin // @[utils.scala 120:29]
          readBuffer_branch_valid <= _GEN_25;
        end else begin
          readBuffer_branch_valid <= _GEN_14;
        end
      end else begin
        readBuffer_branch_valid <= _GEN_14;
      end
    end else begin
      readBuffer_branch_valid <= _GEN_14;
    end
    if (reset) begin // @[ACEUnit.scala 104:28]
      readBuffer_branch_mask <= 5'h0; // @[ACEUnit.scala 104:28]
    end else if (readBuffer_valid) begin // @[ACEUnit.scala 133:25]
      if (readBuffer_branch_valid) begin // @[utils.scala 119:24]
        if (branchOps_valid) begin // @[utils.scala 120:29]
          readBuffer_branch_mask <= _GEN_24;
        end else begin
          readBuffer_branch_mask <= _GEN_15;
        end
      end else begin
        readBuffer_branch_mask <= _GEN_15;
      end
    end else begin
      readBuffer_branch_mask <= _GEN_15;
    end
    if (reset) begin // @[ACEUnit.scala 104:28]
      readBuffer_writeData_valid <= 1'h0; // @[ACEUnit.scala 104:28]
    end else if (readRequest_request_valid & readRequest_request_branch_valid & readRequest_ready) begin // @[ACEUnit.scala 129:91]
      readBuffer_writeData_valid <= readRequest_request_writeData_valid; // @[ACEUnit.scala 130:16]
    end
    if (reset) begin // @[ACEUnit.scala 104:28]
      readBuffer_writeData_data <= 64'h0; // @[ACEUnit.scala 104:28]
    end else if (readRequest_request_valid & readRequest_request_branch_valid & readRequest_ready) begin // @[ACEUnit.scala 129:91]
      readBuffer_writeData_data <= readRequest_request_writeData_data; // @[ACEUnit.scala 130:16]
    end
    if (reset) begin // @[ACEUnit.scala 104:28]
      readBuffer_cacheLine_response <= 2'h0; // @[ACEUnit.scala 104:28]
    end else if (readRequest_request_valid & readRequest_request_branch_valid & readRequest_ready) begin // @[ACEUnit.scala 129:91]
      readBuffer_cacheLine_response <= readRequest_request_cacheLine_response; // @[ACEUnit.scala 130:16]
    end
    if (reset) begin // @[ACEUnit.scala 105:31]
      responseBuffer_valid <= 1'h0; // @[ACEUnit.scala 105:31]
    end else if (2'h0 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
      responseBuffer_valid <= 1'h0; // @[ACEUnit.scala 276:28]
    end else if (!(2'h1 == readACEResponseState)) begin // @[ACEUnit.scala 268:32]
      if (2'h2 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
        responseBuffer_valid <= _GEN_214;
      end
    end
    if (reset) begin // @[ACEUnit.scala 105:31]
      responseBuffer_address <= 32'h0; // @[ACEUnit.scala 105:31]
    end else if (2'h0 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
      if (~ACEMSHR_isEmpty) begin // @[ACEUnit.scala 272:29]
        responseBuffer_address <= ACEMSHR_read_data_address; // @[ACEUnit.scala 274:24]
      end
    end
    if (reset) begin // @[ACEUnit.scala 105:31]
      responseBuffer_core_instruction <= 32'h0; // @[ACEUnit.scala 105:31]
    end else if (2'h0 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
      if (~ACEMSHR_isEmpty) begin // @[ACEUnit.scala 272:29]
        responseBuffer_core_instruction <= ACEMSHR_read_data_core_instruction; // @[ACEUnit.scala 274:24]
      end
    end
    if (reset) begin // @[ACEUnit.scala 105:31]
      responseBuffer_core_robAddr <= 4'h0; // @[ACEUnit.scala 105:31]
    end else if (2'h0 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
      if (~ACEMSHR_isEmpty) begin // @[ACEUnit.scala 272:29]
        responseBuffer_core_robAddr <= ACEMSHR_read_data_core_robAddr; // @[ACEUnit.scala 274:24]
      end
    end
    if (reset) begin // @[ACEUnit.scala 105:31]
      responseBuffer_core_prfDest <= 6'h0; // @[ACEUnit.scala 105:31]
    end else if (2'h0 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
      if (~ACEMSHR_isEmpty) begin // @[ACEUnit.scala 272:29]
        responseBuffer_core_prfDest <= ACEMSHR_read_data_core_prfDest; // @[ACEUnit.scala 274:24]
      end
    end
    if (reset) begin // @[ACEUnit.scala 105:31]
      responseBuffer_branch_valid <= 1'h0; // @[ACEUnit.scala 105:31]
    end else if (responseBuffer_branch_valid) begin // @[utils.scala 119:24]
      if (branchOps_valid) begin // @[utils.scala 120:29]
        if (!(branchOps_passed)) begin // @[utils.scala 121:32]
          responseBuffer_branch_valid <= _GEN_266;
        end
      end else begin
        responseBuffer_branch_valid <= _GEN_244;
      end
    end else begin
      responseBuffer_branch_valid <= _GEN_244;
    end
    if (reset) begin // @[ACEUnit.scala 105:31]
      responseBuffer_branch_mask <= 5'h0; // @[ACEUnit.scala 105:31]
    end else if (responseBuffer_branch_valid) begin // @[utils.scala 119:24]
      if (branchOps_valid) begin // @[utils.scala 120:29]
        if (branchOps_passed) begin // @[utils.scala 121:32]
          responseBuffer_branch_mask <= _GEN_265;
        end else begin
          responseBuffer_branch_mask <= _GEN_267;
        end
      end else begin
        responseBuffer_branch_mask <= _GEN_245;
      end
    end else begin
      responseBuffer_branch_mask <= _GEN_245;
    end
    if (reset) begin // @[ACEUnit.scala 105:31]
      responseBuffer_writeData_valid <= 1'h0; // @[ACEUnit.scala 105:31]
    end else if (2'h0 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
      if (~ACEMSHR_isEmpty) begin // @[ACEUnit.scala 272:29]
        responseBuffer_writeData_valid <= ACEMSHR_read_data_writeData_valid; // @[ACEUnit.scala 274:24]
      end
    end
    if (reset) begin // @[ACEUnit.scala 105:31]
      responseBuffer_writeData_data <= 64'h0; // @[ACEUnit.scala 105:31]
    end else if (2'h0 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
      if (~ACEMSHR_isEmpty) begin // @[ACEUnit.scala 272:29]
        responseBuffer_writeData_data <= ACEMSHR_read_data_writeData_data; // @[ACEUnit.scala 274:24]
      end
    end
    if (reset) begin // @[ACEUnit.scala 105:31]
      responseBuffer_cacheLine_cacheLine <= 512'h0; // @[ACEUnit.scala 105:31]
    end else if (2'h0 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
      if (~ACEMSHR_isEmpty) begin // @[ACEUnit.scala 272:29]
        responseBuffer_cacheLine_cacheLine <= 512'h0; // @[ACEUnit.scala 274:24]
      end
    end else if (!(2'h1 == readACEResponseState)) begin // @[ACEUnit.scala 268:32]
      if (2'h2 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
        responseBuffer_cacheLine_cacheLine <= _responseBuffer_cacheLine_cacheLine_T; // @[ACEUnit.scala 307:42]
      end
    end
    if (reset) begin // @[ACEUnit.scala 105:31]
      responseBuffer_cacheLine_response <= 2'h0; // @[ACEUnit.scala 105:31]
    end else if (2'h0 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
      if (~ACEMSHR_isEmpty) begin // @[ACEUnit.scala 272:29]
        responseBuffer_cacheLine_response <= ACEMSHR_read_data_cacheLine_response; // @[ACEUnit.scala 274:24]
      end
    end else if (!(2'h1 == readACEResponseState)) begin // @[ACEUnit.scala 268:32]
      if (2'h2 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
        responseBuffer_cacheLine_response <= readResponseReg; // @[ACEUnit.scala 308:41]
      end
    end
    if (reset) begin // @[ACEUnit.scala 111:28]
      writeBuffer_valid <= 1'h0; // @[ACEUnit.scala 111:28]
    end else if (2'h0 == writeACEState) begin // @[ACEUnit.scala 174:25]
      writeBuffer_valid <= _GEN_39;
    end else if (2'h1 == writeACEState) begin // @[ACEUnit.scala 174:25]
      writeBuffer_valid <= _GEN_39;
    end else if (2'h2 == writeACEState) begin // @[ACEUnit.scala 174:25]
      writeBuffer_valid <= _GEN_39;
    end else begin
      writeBuffer_valid <= _GEN_61;
    end
    if (reset) begin // @[ACEUnit.scala 111:28]
      writeBuffer_address <= 32'h0; // @[ACEUnit.scala 111:28]
    end else if (_T & writeRequest_request_valid) begin // @[ACEUnit.scala 147:57]
      writeBuffer_address <= writeRequest_request_address; // @[ACEUnit.scala 148:17]
    end
    if (reset) begin // @[ACEUnit.scala 111:28]
      writeBuffer_data <= 512'h0; // @[ACEUnit.scala 111:28]
    end else if (_T & writeRequest_request_valid) begin // @[ACEUnit.scala 147:57]
      writeBuffer_data <= writeRequest_request_data; // @[ACEUnit.scala 148:17]
    end
    if (reset) begin // @[ACEUnit.scala 112:39]
      coherencyRequestBuffer_valid <= 1'h0; // @[ACEUnit.scala 112:39]
    end else if (2'h0 == coherentAXIState) begin // @[ACEUnit.scala 332:27]
      coherencyRequestBuffer_valid <= 1'h0; // @[ACEUnit.scala 339:36]
    end else if (2'h1 == coherentAXIState) begin // @[ACEUnit.scala 332:27]
      if (coherencyRequestBuffer_valid) begin // @[ACEUnit.scala 347:41]
        coherencyRequestBuffer_valid <= _coherencyRequestBuffer_valid_T; // @[ACEUnit.scala 348:37]
      end else begin
        coherencyRequestBuffer_valid <= _GEN_274;
      end
    end
    if (reset) begin // @[ACEUnit.scala 112:39]
      coherencyRequestBuffer_address <= 32'h0; // @[ACEUnit.scala 112:39]
    end else if (2'h0 == coherentAXIState) begin // @[ACEUnit.scala 332:27]
      coherencyRequestBuffer_address <= bus_ACADDR; // @[ACEUnit.scala 340:38]
    end
    if (reset) begin // @[ACEUnit.scala 112:39]
      coherencyRequestBuffer_response <= 2'h0; // @[ACEUnit.scala 112:39]
    end else if (2'h0 == coherentAXIState) begin // @[ACEUnit.scala 332:27]
      coherencyRequestBuffer_response <= _coherencyRequestBuffer_response_T_6; // @[ACEUnit.scala 341:39]
    end
    if (reset) begin // @[ACEUnit.scala 113:40]
      coherencyResponseBuffer_valid <= 1'h0; // @[ACEUnit.scala 113:40]
    end else if (2'h0 == coherentAXIState) begin // @[ACEUnit.scala 332:27]
      coherencyResponseBuffer_valid <= 1'h0; // @[ACEUnit.scala 337:37]
    end else if (_coherencyResponse_ready_T) begin // @[ACEUnit.scala 156:39]
      coherencyResponseBuffer_valid <= coherencyResponse_request_valid; // @[ACEUnit.scala 163:29]
    end
    if (reset) begin // @[ACEUnit.scala 113:40]
      coherencyResponseBuffer_response <= 2'h0; // @[ACEUnit.scala 113:40]
    end else if (_coherencyResponse_ready_T) begin // @[ACEUnit.scala 156:39]
      coherencyResponseBuffer_response <= coherencyResponse_request_response; // @[ACEUnit.scala 163:29]
    end
    if (reset) begin // @[ACEUnit.scala 113:40]
      coherencyResponseBuffer_cacheLine <= 512'h0; // @[ACEUnit.scala 113:40]
    end else if (_coherencyResponse_ready_T) begin // @[ACEUnit.scala 156:39]
      coherencyResponseBuffer_cacheLine <= coherencyResponse_request_cacheLine; // @[ACEUnit.scala 163:29]
    end
    if (reset) begin // @[ACEUnit.scala 113:40]
      coherencyResponseBuffer_dataValid <= 1'h0; // @[ACEUnit.scala 113:40]
    end else if (_coherencyResponse_ready_T) begin // @[ACEUnit.scala 156:39]
      coherencyResponseBuffer_dataValid <= coherencyResponse_request_dataValid; // @[ACEUnit.scala 163:29]
    end
    if (reset) begin // @[ACEUnit.scala 169:30]
      writeACEState <= 2'h0; // @[ACEUnit.scala 169:30]
    end else if (2'h0 == writeACEState) begin // @[ACEUnit.scala 174:25]
      if (writeBuffer_valid) begin // @[ACEUnit.scala 178:29]
        writeACEState <= 2'h1;
      end else begin
        writeACEState <= 2'h0;
      end
    end else if (2'h1 == writeACEState) begin // @[ACEUnit.scala 174:25]
      if (bus_AWREADY) begin // @[ACEUnit.scala 195:27]
        writeACEState <= 2'h2;
      end else begin
        writeACEState <= 2'h1;
      end
    end else if (2'h2 == writeACEState) begin // @[ACEUnit.scala 174:25]
      writeACEState <= _writeACEState_T_3; // @[ACEUnit.scala 211:21]
    end else begin
      writeACEState <= _GEN_62;
    end
    if (reset) begin // @[ACEUnit.scala 224:36]
      readACERequestState <= 1'h0; // @[ACEUnit.scala 224:36]
    end else if (~readACERequestState) begin // @[ACEUnit.scala 225:31]
      readACERequestState <= readBuffer_valid & isCoherencyIdle; // @[ACEUnit.scala 227:27]
    end else if (readACERequestState) begin // @[ACEUnit.scala 225:31]
      if (bus_ARREADY) begin // @[ACEUnit.scala 256:33]
        readACERequestState <= 1'h0;
      end else begin
        readACERequestState <= 1'h1;
      end
    end
    if (reset) begin // @[ACEUnit.scala 326:33]
      coherentAXIState <= 2'h0; // @[ACEUnit.scala 326:33]
    end else if (2'h0 == coherentAXIState) begin // @[ACEUnit.scala 332:27]
      if (bus_ACVALID) begin // @[ACEUnit.scala 343:30]
        coherentAXIState <= 2'h1;
      end else begin
        coherentAXIState <= 2'h0;
      end
    end else if (2'h1 == coherentAXIState) begin // @[ACEUnit.scala 332:27]
      if (isWriteAddressMatchWire & isWireACEBusy) begin // @[ACEUnit.scala 356:53]
        coherentAXIState <= _coherentAXIState_T_1; // @[ACEUnit.scala 357:26]
      end else begin
        coherentAXIState <= _coherentAXIState_T_2; // @[ACEUnit.scala 359:26]
      end
    end else if (2'h2 == coherentAXIState) begin // @[ACEUnit.scala 332:27]
      coherentAXIState <= _GEN_279;
    end else begin
      coherentAXIState <= _GEN_293;
    end
    if (reset) begin // @[ACEUnit.scala 261:37]
      readACEResponseState <= 2'h0; // @[ACEUnit.scala 261:37]
    end else if (2'h0 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
      if (ACEMSHR_read_data_valid & _T_34) begin // @[ACEUnit.scala 278:34]
        readACEResponseState <= 2'h1;
      end else begin
        readACEResponseState <= 2'h0;
      end
    end else if (2'h1 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
      if (isCleanUniqueWire) begin // @[ACEUnit.scala 299:30]
        readACEResponseState <= _readACEResponseState_T_5; // @[ACEUnit.scala 300:30]
      end else begin
        readACEResponseState <= _readACEResponseState_T_8; // @[ACEUnit.scala 302:30]
      end
    end else if (2'h2 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
      readACEResponseState <= _readACEResponseState_T_9; // @[ACEUnit.scala 316:28]
    end
    if (reset) begin // @[ACEUnit.scala 262:28]
      readDataVec_0 <= 64'h0; // @[ACEUnit.scala 262:28]
    end else if (!(2'h0 == readACEResponseState)) begin // @[ACEUnit.scala 268:32]
      if (2'h1 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
        if (!(isCleanUniqueWire)) begin // @[ACEUnit.scala 284:30]
          readDataVec_0 <= _GEN_191;
        end
      end
    end
    if (reset) begin // @[ACEUnit.scala 262:28]
      readDataVec_1 <= 64'h0; // @[ACEUnit.scala 262:28]
    end else if (!(2'h0 == readACEResponseState)) begin // @[ACEUnit.scala 268:32]
      if (2'h1 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
        if (!(isCleanUniqueWire)) begin // @[ACEUnit.scala 284:30]
          readDataVec_1 <= _GEN_192;
        end
      end
    end
    if (reset) begin // @[ACEUnit.scala 262:28]
      readDataVec_2 <= 64'h0; // @[ACEUnit.scala 262:28]
    end else if (!(2'h0 == readACEResponseState)) begin // @[ACEUnit.scala 268:32]
      if (2'h1 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
        if (!(isCleanUniqueWire)) begin // @[ACEUnit.scala 284:30]
          readDataVec_2 <= _GEN_193;
        end
      end
    end
    if (reset) begin // @[ACEUnit.scala 262:28]
      readDataVec_3 <= 64'h0; // @[ACEUnit.scala 262:28]
    end else if (!(2'h0 == readACEResponseState)) begin // @[ACEUnit.scala 268:32]
      if (2'h1 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
        if (!(isCleanUniqueWire)) begin // @[ACEUnit.scala 284:30]
          readDataVec_3 <= _GEN_194;
        end
      end
    end
    if (reset) begin // @[ACEUnit.scala 262:28]
      readDataVec_4 <= 64'h0; // @[ACEUnit.scala 262:28]
    end else if (!(2'h0 == readACEResponseState)) begin // @[ACEUnit.scala 268:32]
      if (2'h1 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
        if (!(isCleanUniqueWire)) begin // @[ACEUnit.scala 284:30]
          readDataVec_4 <= _GEN_195;
        end
      end
    end
    if (reset) begin // @[ACEUnit.scala 262:28]
      readDataVec_5 <= 64'h0; // @[ACEUnit.scala 262:28]
    end else if (!(2'h0 == readACEResponseState)) begin // @[ACEUnit.scala 268:32]
      if (2'h1 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
        if (!(isCleanUniqueWire)) begin // @[ACEUnit.scala 284:30]
          readDataVec_5 <= _GEN_196;
        end
      end
    end
    if (reset) begin // @[ACEUnit.scala 262:28]
      readDataVec_6 <= 64'h0; // @[ACEUnit.scala 262:28]
    end else if (!(2'h0 == readACEResponseState)) begin // @[ACEUnit.scala 268:32]
      if (2'h1 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
        if (!(isCleanUniqueWire)) begin // @[ACEUnit.scala 284:30]
          readDataVec_6 <= _GEN_197;
        end
      end
    end
    if (reset) begin // @[ACEUnit.scala 262:28]
      readDataVec_7 <= 64'h0; // @[ACEUnit.scala 262:28]
    end else if (!(2'h0 == readACEResponseState)) begin // @[ACEUnit.scala 268:32]
      if (2'h1 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
        if (!(isCleanUniqueWire)) begin // @[ACEUnit.scala 284:30]
          readDataVec_7 <= _GEN_198;
        end
      end
    end
    readResponseValid <= reset | _GEN_254; // @[ACEUnit.scala 263:{34,34}]
    if (reset) begin // @[ACEUnit.scala 264:32]
      readResponseReg <= 2'h0; // @[ACEUnit.scala 264:32]
    end else if (!(2'h0 == readACEResponseState)) begin // @[ACEUnit.scala 268:32]
      if (2'h1 == readACEResponseState) begin // @[ACEUnit.scala 268:32]
        if (isCleanUniqueWire) begin // @[ACEUnit.scala 284:30]
          readResponseReg <= bus_RRESP[3:2]; // @[ACEUnit.scala 285:25]
        end else begin
          readResponseReg <= _GEN_200;
        end
      end
    end
    if (reset) begin // @[ACEUnit.scala 328:36]
      coherentRequestSend <= 1'h0; // @[ACEUnit.scala 328:36]
    end else if (2'h0 == coherentAXIState) begin // @[ACEUnit.scala 332:27]
      coherentRequestSend <= 1'h0; // @[ACEUnit.scala 334:27]
    end else if (2'h1 == coherentAXIState) begin // @[ACEUnit.scala 332:27]
      if (!(coherencyRequestBuffer_valid)) begin // @[ACEUnit.scala 347:41]
        coherentRequestSend <= _GEN_275;
      end
    end else if (2'h2 == coherentAXIState) begin // @[ACEUnit.scala 332:27]
      coherentRequestSend <= 1'h0; // @[ACEUnit.scala 363:27]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  readBuffer_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  readBuffer_address = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  readBuffer_core_instruction = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  readBuffer_core_robAddr = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  readBuffer_core_prfDest = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  readBuffer_branch_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  readBuffer_branch_mask = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  readBuffer_writeData_valid = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  readBuffer_writeData_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  readBuffer_cacheLine_response = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  responseBuffer_valid = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  responseBuffer_address = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  responseBuffer_core_instruction = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  responseBuffer_core_robAddr = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  responseBuffer_core_prfDest = _RAND_14[5:0];
  _RAND_15 = {1{`RANDOM}};
  responseBuffer_branch_valid = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  responseBuffer_branch_mask = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  responseBuffer_writeData_valid = _RAND_17[0:0];
  _RAND_18 = {2{`RANDOM}};
  responseBuffer_writeData_data = _RAND_18[63:0];
  _RAND_19 = {16{`RANDOM}};
  responseBuffer_cacheLine_cacheLine = _RAND_19[511:0];
  _RAND_20 = {1{`RANDOM}};
  responseBuffer_cacheLine_response = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  writeBuffer_valid = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  writeBuffer_address = _RAND_22[31:0];
  _RAND_23 = {16{`RANDOM}};
  writeBuffer_data = _RAND_23[511:0];
  _RAND_24 = {1{`RANDOM}};
  coherencyRequestBuffer_valid = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  coherencyRequestBuffer_address = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  coherencyRequestBuffer_response = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  coherencyResponseBuffer_valid = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  coherencyResponseBuffer_response = _RAND_28[1:0];
  _RAND_29 = {16{`RANDOM}};
  coherencyResponseBuffer_cacheLine = _RAND_29[511:0];
  _RAND_30 = {1{`RANDOM}};
  coherencyResponseBuffer_dataValid = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  writeACEState = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  readACERequestState = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  coherentAXIState = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  readACEResponseState = _RAND_34[1:0];
  _RAND_35 = {2{`RANDOM}};
  readDataVec_0 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  readDataVec_1 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  readDataVec_2 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  readDataVec_3 = _RAND_38[63:0];
  _RAND_39 = {2{`RANDOM}};
  readDataVec_4 = _RAND_39[63:0];
  _RAND_40 = {2{`RANDOM}};
  readDataVec_5 = _RAND_40[63:0];
  _RAND_41 = {2{`RANDOM}};
  readDataVec_6 = _RAND_41[63:0];
  _RAND_42 = {2{`RANDOM}};
  readDataVec_7 = _RAND_42[63:0];
  _RAND_43 = {1{`RANDOM}};
  readResponseValid = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  readResponseReg = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  coherentRequestSend = _RAND_45[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module fifoRecordInvalidateI(
  input         clock,
  input         reset,
  input         write_data_valid,
  input  [31:0] write_data_address,
  input         write_data_branch_valid,
  input  [4:0]  write_data_branch_mask,
  input         read_ready,
  output        read_data_valid,
  output        read_data_branch_valid,
  output        isEmpty,
  input         branchOps_valid,
  input  [4:0]  branchOps_branchMask,
  input         branchOps_passed,
  output        isFull,
  input  [31:0] invalidateAddr,
  input         invalidateEnable
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
`endif // RANDOMIZE_REG_INIT
  reg  memReg_0_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_0_address; // @[fifo.scala 27:33]
  reg  memReg_0_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_0_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_1_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_1_address; // @[fifo.scala 27:33]
  reg  memReg_1_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_1_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_2_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_2_address; // @[fifo.scala 27:33]
  reg  memReg_2_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_2_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_3_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_3_address; // @[fifo.scala 27:33]
  reg  memReg_3_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_3_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_4_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_4_address; // @[fifo.scala 27:33]
  reg  memReg_4_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_4_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_5_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_5_address; // @[fifo.scala 27:33]
  reg  memReg_5_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_5_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_6_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_6_address; // @[fifo.scala 27:33]
  reg  memReg_6_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_6_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_7_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_7_address; // @[fifo.scala 27:33]
  reg  memReg_7_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_7_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_8_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_8_address; // @[fifo.scala 27:33]
  reg  memReg_8_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_8_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_9_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_9_address; // @[fifo.scala 27:33]
  reg  memReg_9_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_9_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_10_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_10_address; // @[fifo.scala 27:33]
  reg  memReg_10_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_10_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_11_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_11_address; // @[fifo.scala 27:33]
  reg  memReg_11_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_11_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_12_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_12_address; // @[fifo.scala 27:33]
  reg  memReg_12_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_12_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_13_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_13_address; // @[fifo.scala 27:33]
  reg  memReg_13_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_13_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_14_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_14_address; // @[fifo.scala 27:33]
  reg  memReg_14_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_14_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_15_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_15_address; // @[fifo.scala 27:33]
  reg  memReg_15_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_15_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_16_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_16_address; // @[fifo.scala 27:33]
  reg  memReg_16_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_16_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_17_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_17_address; // @[fifo.scala 27:33]
  reg  memReg_17_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_17_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_18_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_18_address; // @[fifo.scala 27:33]
  reg  memReg_18_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_18_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_19_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_19_address; // @[fifo.scala 27:33]
  reg  memReg_19_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_19_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_20_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_20_address; // @[fifo.scala 27:33]
  reg  memReg_20_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_20_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_21_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_21_address; // @[fifo.scala 27:33]
  reg  memReg_21_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_21_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_22_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_22_address; // @[fifo.scala 27:33]
  reg  memReg_22_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_22_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_23_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_23_address; // @[fifo.scala 27:33]
  reg  memReg_23_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_23_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_24_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_24_address; // @[fifo.scala 27:33]
  reg  memReg_24_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_24_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_25_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_25_address; // @[fifo.scala 27:33]
  reg  memReg_25_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_25_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_26_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_26_address; // @[fifo.scala 27:33]
  reg  memReg_26_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_26_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_27_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_27_address; // @[fifo.scala 27:33]
  reg  memReg_27_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_27_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_28_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_28_address; // @[fifo.scala 27:33]
  reg  memReg_28_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_28_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_29_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_29_address; // @[fifo.scala 27:33]
  reg  memReg_29_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_29_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_30_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_30_address; // @[fifo.scala 27:33]
  reg  memReg_30_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_30_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_31_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_31_address; // @[fifo.scala 27:33]
  reg  memReg_31_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_31_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_32_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_32_address; // @[fifo.scala 27:33]
  reg  memReg_32_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_32_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_33_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_33_address; // @[fifo.scala 27:33]
  reg  memReg_33_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_33_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_34_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_34_address; // @[fifo.scala 27:33]
  reg  memReg_34_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_34_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_35_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_35_address; // @[fifo.scala 27:33]
  reg  memReg_35_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_35_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_36_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_36_address; // @[fifo.scala 27:33]
  reg  memReg_36_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_36_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_37_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_37_address; // @[fifo.scala 27:33]
  reg  memReg_37_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_37_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_38_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_38_address; // @[fifo.scala 27:33]
  reg  memReg_38_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_38_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_39_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_39_address; // @[fifo.scala 27:33]
  reg  memReg_39_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_39_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_40_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_40_address; // @[fifo.scala 27:33]
  reg  memReg_40_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_40_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_41_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_41_address; // @[fifo.scala 27:33]
  reg  memReg_41_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_41_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_42_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_42_address; // @[fifo.scala 27:33]
  reg  memReg_42_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_42_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_43_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_43_address; // @[fifo.scala 27:33]
  reg  memReg_43_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_43_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_44_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_44_address; // @[fifo.scala 27:33]
  reg  memReg_44_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_44_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_45_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_45_address; // @[fifo.scala 27:33]
  reg  memReg_45_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_45_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_46_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_46_address; // @[fifo.scala 27:33]
  reg  memReg_46_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_46_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_47_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_47_address; // @[fifo.scala 27:33]
  reg  memReg_47_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_47_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_48_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_48_address; // @[fifo.scala 27:33]
  reg  memReg_48_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_48_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_49_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_49_address; // @[fifo.scala 27:33]
  reg  memReg_49_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_49_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_50_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_50_address; // @[fifo.scala 27:33]
  reg  memReg_50_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_50_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_51_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_51_address; // @[fifo.scala 27:33]
  reg  memReg_51_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_51_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_52_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_52_address; // @[fifo.scala 27:33]
  reg  memReg_52_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_52_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_53_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_53_address; // @[fifo.scala 27:33]
  reg  memReg_53_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_53_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_54_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_54_address; // @[fifo.scala 27:33]
  reg  memReg_54_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_54_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_55_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_55_address; // @[fifo.scala 27:33]
  reg  memReg_55_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_55_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_56_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_56_address; // @[fifo.scala 27:33]
  reg  memReg_56_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_56_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_57_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_57_address; // @[fifo.scala 27:33]
  reg  memReg_57_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_57_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_58_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_58_address; // @[fifo.scala 27:33]
  reg  memReg_58_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_58_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_59_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_59_address; // @[fifo.scala 27:33]
  reg  memReg_59_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_59_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_60_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_60_address; // @[fifo.scala 27:33]
  reg  memReg_60_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_60_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_61_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_61_address; // @[fifo.scala 27:33]
  reg  memReg_61_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_61_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_62_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_62_address; // @[fifo.scala 27:33]
  reg  memReg_62_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_62_branch_mask; // @[fifo.scala 27:33]
  reg  memReg_63_valid; // @[fifo.scala 27:33]
  reg [31:0] memReg_63_address; // @[fifo.scala 27:33]
  reg  memReg_63_branch_valid; // @[fifo.scala 27:33]
  reg [4:0] memReg_63_branch_mask; // @[fifo.scala 27:33]
  reg [5:0] readPtr; // @[fifo.scala 33:25]
  wire [5:0] _nextVal_T_2 = readPtr + 6'h1; // @[fifo.scala 34:60]
  wire [5:0] nextRead = readPtr == 6'h3f ? 6'h0 : _nextVal_T_2; // @[fifo.scala 34:22]
  wire [1:0] op = {write_data_valid,read_ready}; // @[fifo.scala 46:29]
  reg  emptyReg; // @[fifo.scala 43:25]
  wire  _T_2 = ~emptyReg; // @[fifo.scala 52:12]
  wire  _GEN_21 = 2'h2 == op ? 1'h0 : 2'h3 == op & _T_2; // @[fifo.scala 49:14]
  wire  _GEN_24 = 2'h1 == op ? _T_2 : _GEN_21; // @[fifo.scala 49:14]
  wire  incrRead = 2'h0 == op ? 1'h0 : _GEN_24; // @[fifo.scala 49:14]
  reg [5:0] writePtr; // @[fifo.scala 33:25]
  wire [5:0] _nextVal_T_5 = writePtr + 6'h1; // @[fifo.scala 34:60]
  wire [5:0] nextWrite = writePtr == 6'h3f ? 6'h0 : _nextVal_T_5; // @[fifo.scala 34:22]
  reg  fullReg; // @[fifo.scala 44:34]
  wire  _T_4 = ~fullReg; // @[fifo.scala 59:12]
  wire  _GEN_18 = 2'h2 == op ? _T_4 : 2'h3 == op & _T_4; // @[fifo.scala 49:14]
  wire  _GEN_25 = 2'h1 == op ? 1'h0 : _GEN_18; // @[fifo.scala 49:14]
  wire  incrWrite = 2'h0 == op ? 1'h0 : _GEN_25; // @[fifo.scala 49:14]
  wire  _GEN_3 = ~emptyReg ? nextRead == writePtr : emptyReg; // @[fifo.scala 52:23 54:18 43:25]
  wire  _GEN_6 = ~fullReg ? 1'h0 : emptyReg; // @[fifo.scala 59:22 61:18 43:25]
  wire  _GEN_7 = ~fullReg ? nextWrite == readPtr : fullReg; // @[fifo.scala 59:22 62:17 44:34]
  wire  _fullReg_T_2 = emptyReg ? 1'h0 : nextWrite == nextRead; // @[fifo.scala 70:23]
  wire  _GEN_10 = _T_4 ? _fullReg_T_2 : fullReg; // @[fifo.scala 67:22 70:17 44:34]
  wire  _emptyReg_T_2 = fullReg ? 1'h0 : nextRead == nextWrite; // @[fifo.scala 75:24]
  wire  _GEN_11 = _T_2 ? 1'h0 : _GEN_10; // @[fifo.scala 73:23 74:17]
  wire  _GEN_12 = _T_2 ? _emptyReg_T_2 : _GEN_6; // @[fifo.scala 73:23 75:18]
  wire  _GEN_15 = 2'h3 == op ? _GEN_12 : emptyReg; // @[fifo.scala 49:14 43:25]
  wire  _GEN_16 = 2'h3 == op ? _GEN_11 : fullReg; // @[fifo.scala 49:14 44:34]
  wire  _GEN_19 = 2'h2 == op ? _GEN_6 : _GEN_15; // @[fifo.scala 49:14]
  wire  _GEN_23 = 2'h1 == op ? _GEN_3 : _GEN_19; // @[fifo.scala 49:14]
  wire  _GEN_27 = 2'h0 == op ? emptyReg : _GEN_23; // @[fifo.scala 49:14 43:25]
  wire  _GEN_30 = 6'h0 == writePtr ? write_data_valid : memReg_0_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_31 = 6'h1 == writePtr ? write_data_valid : memReg_1_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_32 = 6'h2 == writePtr ? write_data_valid : memReg_2_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_33 = 6'h3 == writePtr ? write_data_valid : memReg_3_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_34 = 6'h4 == writePtr ? write_data_valid : memReg_4_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_35 = 6'h5 == writePtr ? write_data_valid : memReg_5_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_36 = 6'h6 == writePtr ? write_data_valid : memReg_6_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_37 = 6'h7 == writePtr ? write_data_valid : memReg_7_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_38 = 6'h8 == writePtr ? write_data_valid : memReg_8_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_39 = 6'h9 == writePtr ? write_data_valid : memReg_9_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_40 = 6'ha == writePtr ? write_data_valid : memReg_10_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_41 = 6'hb == writePtr ? write_data_valid : memReg_11_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_42 = 6'hc == writePtr ? write_data_valid : memReg_12_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_43 = 6'hd == writePtr ? write_data_valid : memReg_13_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_44 = 6'he == writePtr ? write_data_valid : memReg_14_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_45 = 6'hf == writePtr ? write_data_valid : memReg_15_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_46 = 6'h10 == writePtr ? write_data_valid : memReg_16_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_47 = 6'h11 == writePtr ? write_data_valid : memReg_17_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_48 = 6'h12 == writePtr ? write_data_valid : memReg_18_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_49 = 6'h13 == writePtr ? write_data_valid : memReg_19_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_50 = 6'h14 == writePtr ? write_data_valid : memReg_20_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_51 = 6'h15 == writePtr ? write_data_valid : memReg_21_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_52 = 6'h16 == writePtr ? write_data_valid : memReg_22_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_53 = 6'h17 == writePtr ? write_data_valid : memReg_23_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_54 = 6'h18 == writePtr ? write_data_valid : memReg_24_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_55 = 6'h19 == writePtr ? write_data_valid : memReg_25_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_56 = 6'h1a == writePtr ? write_data_valid : memReg_26_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_57 = 6'h1b == writePtr ? write_data_valid : memReg_27_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_58 = 6'h1c == writePtr ? write_data_valid : memReg_28_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_59 = 6'h1d == writePtr ? write_data_valid : memReg_29_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_60 = 6'h1e == writePtr ? write_data_valid : memReg_30_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_61 = 6'h1f == writePtr ? write_data_valid : memReg_31_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_62 = 6'h20 == writePtr ? write_data_valid : memReg_32_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_63 = 6'h21 == writePtr ? write_data_valid : memReg_33_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_64 = 6'h22 == writePtr ? write_data_valid : memReg_34_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_65 = 6'h23 == writePtr ? write_data_valid : memReg_35_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_66 = 6'h24 == writePtr ? write_data_valid : memReg_36_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_67 = 6'h25 == writePtr ? write_data_valid : memReg_37_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_68 = 6'h26 == writePtr ? write_data_valid : memReg_38_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_69 = 6'h27 == writePtr ? write_data_valid : memReg_39_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_70 = 6'h28 == writePtr ? write_data_valid : memReg_40_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_71 = 6'h29 == writePtr ? write_data_valid : memReg_41_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_72 = 6'h2a == writePtr ? write_data_valid : memReg_42_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_73 = 6'h2b == writePtr ? write_data_valid : memReg_43_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_74 = 6'h2c == writePtr ? write_data_valid : memReg_44_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_75 = 6'h2d == writePtr ? write_data_valid : memReg_45_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_76 = 6'h2e == writePtr ? write_data_valid : memReg_46_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_77 = 6'h2f == writePtr ? write_data_valid : memReg_47_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_78 = 6'h30 == writePtr ? write_data_valid : memReg_48_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_79 = 6'h31 == writePtr ? write_data_valid : memReg_49_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_80 = 6'h32 == writePtr ? write_data_valid : memReg_50_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_81 = 6'h33 == writePtr ? write_data_valid : memReg_51_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_82 = 6'h34 == writePtr ? write_data_valid : memReg_52_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_83 = 6'h35 == writePtr ? write_data_valid : memReg_53_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_84 = 6'h36 == writePtr ? write_data_valid : memReg_54_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_85 = 6'h37 == writePtr ? write_data_valid : memReg_55_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_86 = 6'h38 == writePtr ? write_data_valid : memReg_56_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_87 = 6'h39 == writePtr ? write_data_valid : memReg_57_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_88 = 6'h3a == writePtr ? write_data_valid : memReg_58_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_89 = 6'h3b == writePtr ? write_data_valid : memReg_59_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_90 = 6'h3c == writePtr ? write_data_valid : memReg_60_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_91 = 6'h3d == writePtr ? write_data_valid : memReg_61_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_92 = 6'h3e == writePtr ? write_data_valid : memReg_62_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_93 = 6'h3f == writePtr ? write_data_valid : memReg_63_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_350 = 6'h0 == writePtr ? write_data_branch_valid : memReg_0_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_351 = 6'h1 == writePtr ? write_data_branch_valid : memReg_1_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_352 = 6'h2 == writePtr ? write_data_branch_valid : memReg_2_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_353 = 6'h3 == writePtr ? write_data_branch_valid : memReg_3_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_354 = 6'h4 == writePtr ? write_data_branch_valid : memReg_4_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_355 = 6'h5 == writePtr ? write_data_branch_valid : memReg_5_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_356 = 6'h6 == writePtr ? write_data_branch_valid : memReg_6_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_357 = 6'h7 == writePtr ? write_data_branch_valid : memReg_7_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_358 = 6'h8 == writePtr ? write_data_branch_valid : memReg_8_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_359 = 6'h9 == writePtr ? write_data_branch_valid : memReg_9_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_360 = 6'ha == writePtr ? write_data_branch_valid : memReg_10_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_361 = 6'hb == writePtr ? write_data_branch_valid : memReg_11_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_362 = 6'hc == writePtr ? write_data_branch_valid : memReg_12_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_363 = 6'hd == writePtr ? write_data_branch_valid : memReg_13_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_364 = 6'he == writePtr ? write_data_branch_valid : memReg_14_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_365 = 6'hf == writePtr ? write_data_branch_valid : memReg_15_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_366 = 6'h10 == writePtr ? write_data_branch_valid : memReg_16_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_367 = 6'h11 == writePtr ? write_data_branch_valid : memReg_17_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_368 = 6'h12 == writePtr ? write_data_branch_valid : memReg_18_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_369 = 6'h13 == writePtr ? write_data_branch_valid : memReg_19_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_370 = 6'h14 == writePtr ? write_data_branch_valid : memReg_20_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_371 = 6'h15 == writePtr ? write_data_branch_valid : memReg_21_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_372 = 6'h16 == writePtr ? write_data_branch_valid : memReg_22_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_373 = 6'h17 == writePtr ? write_data_branch_valid : memReg_23_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_374 = 6'h18 == writePtr ? write_data_branch_valid : memReg_24_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_375 = 6'h19 == writePtr ? write_data_branch_valid : memReg_25_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_376 = 6'h1a == writePtr ? write_data_branch_valid : memReg_26_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_377 = 6'h1b == writePtr ? write_data_branch_valid : memReg_27_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_378 = 6'h1c == writePtr ? write_data_branch_valid : memReg_28_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_379 = 6'h1d == writePtr ? write_data_branch_valid : memReg_29_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_380 = 6'h1e == writePtr ? write_data_branch_valid : memReg_30_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_381 = 6'h1f == writePtr ? write_data_branch_valid : memReg_31_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_382 = 6'h20 == writePtr ? write_data_branch_valid : memReg_32_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_383 = 6'h21 == writePtr ? write_data_branch_valid : memReg_33_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_384 = 6'h22 == writePtr ? write_data_branch_valid : memReg_34_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_385 = 6'h23 == writePtr ? write_data_branch_valid : memReg_35_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_386 = 6'h24 == writePtr ? write_data_branch_valid : memReg_36_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_387 = 6'h25 == writePtr ? write_data_branch_valid : memReg_37_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_388 = 6'h26 == writePtr ? write_data_branch_valid : memReg_38_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_389 = 6'h27 == writePtr ? write_data_branch_valid : memReg_39_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_390 = 6'h28 == writePtr ? write_data_branch_valid : memReg_40_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_391 = 6'h29 == writePtr ? write_data_branch_valid : memReg_41_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_392 = 6'h2a == writePtr ? write_data_branch_valid : memReg_42_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_393 = 6'h2b == writePtr ? write_data_branch_valid : memReg_43_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_394 = 6'h2c == writePtr ? write_data_branch_valid : memReg_44_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_395 = 6'h2d == writePtr ? write_data_branch_valid : memReg_45_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_396 = 6'h2e == writePtr ? write_data_branch_valid : memReg_46_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_397 = 6'h2f == writePtr ? write_data_branch_valid : memReg_47_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_398 = 6'h30 == writePtr ? write_data_branch_valid : memReg_48_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_399 = 6'h31 == writePtr ? write_data_branch_valid : memReg_49_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_400 = 6'h32 == writePtr ? write_data_branch_valid : memReg_50_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_401 = 6'h33 == writePtr ? write_data_branch_valid : memReg_51_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_402 = 6'h34 == writePtr ? write_data_branch_valid : memReg_52_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_403 = 6'h35 == writePtr ? write_data_branch_valid : memReg_53_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_404 = 6'h36 == writePtr ? write_data_branch_valid : memReg_54_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_405 = 6'h37 == writePtr ? write_data_branch_valid : memReg_55_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_406 = 6'h38 == writePtr ? write_data_branch_valid : memReg_56_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_407 = 6'h39 == writePtr ? write_data_branch_valid : memReg_57_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_408 = 6'h3a == writePtr ? write_data_branch_valid : memReg_58_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_409 = 6'h3b == writePtr ? write_data_branch_valid : memReg_59_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_410 = 6'h3c == writePtr ? write_data_branch_valid : memReg_60_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_411 = 6'h3d == writePtr ? write_data_branch_valid : memReg_61_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_412 = 6'h3e == writePtr ? write_data_branch_valid : memReg_62_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_413 = 6'h3f == writePtr ? write_data_branch_valid : memReg_63_branch_valid; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_414 = 6'h0 == writePtr ? write_data_branch_mask : memReg_0_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_415 = 6'h1 == writePtr ? write_data_branch_mask : memReg_1_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_416 = 6'h2 == writePtr ? write_data_branch_mask : memReg_2_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_417 = 6'h3 == writePtr ? write_data_branch_mask : memReg_3_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_418 = 6'h4 == writePtr ? write_data_branch_mask : memReg_4_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_419 = 6'h5 == writePtr ? write_data_branch_mask : memReg_5_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_420 = 6'h6 == writePtr ? write_data_branch_mask : memReg_6_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_421 = 6'h7 == writePtr ? write_data_branch_mask : memReg_7_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_422 = 6'h8 == writePtr ? write_data_branch_mask : memReg_8_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_423 = 6'h9 == writePtr ? write_data_branch_mask : memReg_9_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_424 = 6'ha == writePtr ? write_data_branch_mask : memReg_10_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_425 = 6'hb == writePtr ? write_data_branch_mask : memReg_11_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_426 = 6'hc == writePtr ? write_data_branch_mask : memReg_12_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_427 = 6'hd == writePtr ? write_data_branch_mask : memReg_13_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_428 = 6'he == writePtr ? write_data_branch_mask : memReg_14_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_429 = 6'hf == writePtr ? write_data_branch_mask : memReg_15_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_430 = 6'h10 == writePtr ? write_data_branch_mask : memReg_16_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_431 = 6'h11 == writePtr ? write_data_branch_mask : memReg_17_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_432 = 6'h12 == writePtr ? write_data_branch_mask : memReg_18_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_433 = 6'h13 == writePtr ? write_data_branch_mask : memReg_19_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_434 = 6'h14 == writePtr ? write_data_branch_mask : memReg_20_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_435 = 6'h15 == writePtr ? write_data_branch_mask : memReg_21_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_436 = 6'h16 == writePtr ? write_data_branch_mask : memReg_22_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_437 = 6'h17 == writePtr ? write_data_branch_mask : memReg_23_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_438 = 6'h18 == writePtr ? write_data_branch_mask : memReg_24_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_439 = 6'h19 == writePtr ? write_data_branch_mask : memReg_25_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_440 = 6'h1a == writePtr ? write_data_branch_mask : memReg_26_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_441 = 6'h1b == writePtr ? write_data_branch_mask : memReg_27_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_442 = 6'h1c == writePtr ? write_data_branch_mask : memReg_28_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_443 = 6'h1d == writePtr ? write_data_branch_mask : memReg_29_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_444 = 6'h1e == writePtr ? write_data_branch_mask : memReg_30_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_445 = 6'h1f == writePtr ? write_data_branch_mask : memReg_31_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_446 = 6'h20 == writePtr ? write_data_branch_mask : memReg_32_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_447 = 6'h21 == writePtr ? write_data_branch_mask : memReg_33_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_448 = 6'h22 == writePtr ? write_data_branch_mask : memReg_34_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_449 = 6'h23 == writePtr ? write_data_branch_mask : memReg_35_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_450 = 6'h24 == writePtr ? write_data_branch_mask : memReg_36_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_451 = 6'h25 == writePtr ? write_data_branch_mask : memReg_37_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_452 = 6'h26 == writePtr ? write_data_branch_mask : memReg_38_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_453 = 6'h27 == writePtr ? write_data_branch_mask : memReg_39_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_454 = 6'h28 == writePtr ? write_data_branch_mask : memReg_40_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_455 = 6'h29 == writePtr ? write_data_branch_mask : memReg_41_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_456 = 6'h2a == writePtr ? write_data_branch_mask : memReg_42_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_457 = 6'h2b == writePtr ? write_data_branch_mask : memReg_43_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_458 = 6'h2c == writePtr ? write_data_branch_mask : memReg_44_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_459 = 6'h2d == writePtr ? write_data_branch_mask : memReg_45_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_460 = 6'h2e == writePtr ? write_data_branch_mask : memReg_46_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_461 = 6'h2f == writePtr ? write_data_branch_mask : memReg_47_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_462 = 6'h30 == writePtr ? write_data_branch_mask : memReg_48_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_463 = 6'h31 == writePtr ? write_data_branch_mask : memReg_49_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_464 = 6'h32 == writePtr ? write_data_branch_mask : memReg_50_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_465 = 6'h33 == writePtr ? write_data_branch_mask : memReg_51_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_466 = 6'h34 == writePtr ? write_data_branch_mask : memReg_52_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_467 = 6'h35 == writePtr ? write_data_branch_mask : memReg_53_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_468 = 6'h36 == writePtr ? write_data_branch_mask : memReg_54_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_469 = 6'h37 == writePtr ? write_data_branch_mask : memReg_55_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_470 = 6'h38 == writePtr ? write_data_branch_mask : memReg_56_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_471 = 6'h39 == writePtr ? write_data_branch_mask : memReg_57_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_472 = 6'h3a == writePtr ? write_data_branch_mask : memReg_58_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_473 = 6'h3b == writePtr ? write_data_branch_mask : memReg_59_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_474 = 6'h3c == writePtr ? write_data_branch_mask : memReg_60_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_475 = 6'h3d == writePtr ? write_data_branch_mask : memReg_61_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_476 = 6'h3e == writePtr ? write_data_branch_mask : memReg_62_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire [4:0] _GEN_477 = 6'h3f == writePtr ? write_data_branch_mask : memReg_63_branch_mask; // @[fifo.scala 82:{22,22} 27:33]
  wire  _GEN_798 = incrWrite ? _GEN_30 : memReg_0_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_799 = incrWrite ? _GEN_31 : memReg_1_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_800 = incrWrite ? _GEN_32 : memReg_2_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_801 = incrWrite ? _GEN_33 : memReg_3_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_802 = incrWrite ? _GEN_34 : memReg_4_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_803 = incrWrite ? _GEN_35 : memReg_5_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_804 = incrWrite ? _GEN_36 : memReg_6_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_805 = incrWrite ? _GEN_37 : memReg_7_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_806 = incrWrite ? _GEN_38 : memReg_8_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_807 = incrWrite ? _GEN_39 : memReg_9_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_808 = incrWrite ? _GEN_40 : memReg_10_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_809 = incrWrite ? _GEN_41 : memReg_11_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_810 = incrWrite ? _GEN_42 : memReg_12_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_811 = incrWrite ? _GEN_43 : memReg_13_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_812 = incrWrite ? _GEN_44 : memReg_14_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_813 = incrWrite ? _GEN_45 : memReg_15_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_814 = incrWrite ? _GEN_46 : memReg_16_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_815 = incrWrite ? _GEN_47 : memReg_17_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_816 = incrWrite ? _GEN_48 : memReg_18_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_817 = incrWrite ? _GEN_49 : memReg_19_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_818 = incrWrite ? _GEN_50 : memReg_20_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_819 = incrWrite ? _GEN_51 : memReg_21_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_820 = incrWrite ? _GEN_52 : memReg_22_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_821 = incrWrite ? _GEN_53 : memReg_23_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_822 = incrWrite ? _GEN_54 : memReg_24_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_823 = incrWrite ? _GEN_55 : memReg_25_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_824 = incrWrite ? _GEN_56 : memReg_26_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_825 = incrWrite ? _GEN_57 : memReg_27_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_826 = incrWrite ? _GEN_58 : memReg_28_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_827 = incrWrite ? _GEN_59 : memReg_29_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_828 = incrWrite ? _GEN_60 : memReg_30_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_829 = incrWrite ? _GEN_61 : memReg_31_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_830 = incrWrite ? _GEN_62 : memReg_32_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_831 = incrWrite ? _GEN_63 : memReg_33_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_832 = incrWrite ? _GEN_64 : memReg_34_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_833 = incrWrite ? _GEN_65 : memReg_35_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_834 = incrWrite ? _GEN_66 : memReg_36_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_835 = incrWrite ? _GEN_67 : memReg_37_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_836 = incrWrite ? _GEN_68 : memReg_38_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_837 = incrWrite ? _GEN_69 : memReg_39_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_838 = incrWrite ? _GEN_70 : memReg_40_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_839 = incrWrite ? _GEN_71 : memReg_41_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_840 = incrWrite ? _GEN_72 : memReg_42_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_841 = incrWrite ? _GEN_73 : memReg_43_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_842 = incrWrite ? _GEN_74 : memReg_44_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_843 = incrWrite ? _GEN_75 : memReg_45_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_844 = incrWrite ? _GEN_76 : memReg_46_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_845 = incrWrite ? _GEN_77 : memReg_47_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_846 = incrWrite ? _GEN_78 : memReg_48_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_847 = incrWrite ? _GEN_79 : memReg_49_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_848 = incrWrite ? _GEN_80 : memReg_50_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_849 = incrWrite ? _GEN_81 : memReg_51_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_850 = incrWrite ? _GEN_82 : memReg_52_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_851 = incrWrite ? _GEN_83 : memReg_53_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_852 = incrWrite ? _GEN_84 : memReg_54_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_853 = incrWrite ? _GEN_85 : memReg_55_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_854 = incrWrite ? _GEN_86 : memReg_56_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_855 = incrWrite ? _GEN_87 : memReg_57_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_856 = incrWrite ? _GEN_88 : memReg_58_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_857 = incrWrite ? _GEN_89 : memReg_59_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_858 = incrWrite ? _GEN_90 : memReg_60_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_859 = incrWrite ? _GEN_91 : memReg_61_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_860 = incrWrite ? _GEN_92 : memReg_62_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_861 = incrWrite ? _GEN_93 : memReg_63_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1118 = incrWrite ? _GEN_350 : memReg_0_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1119 = incrWrite ? _GEN_351 : memReg_1_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1120 = incrWrite ? _GEN_352 : memReg_2_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1121 = incrWrite ? _GEN_353 : memReg_3_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1122 = incrWrite ? _GEN_354 : memReg_4_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1123 = incrWrite ? _GEN_355 : memReg_5_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1124 = incrWrite ? _GEN_356 : memReg_6_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1125 = incrWrite ? _GEN_357 : memReg_7_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1126 = incrWrite ? _GEN_358 : memReg_8_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1127 = incrWrite ? _GEN_359 : memReg_9_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1128 = incrWrite ? _GEN_360 : memReg_10_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1129 = incrWrite ? _GEN_361 : memReg_11_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1130 = incrWrite ? _GEN_362 : memReg_12_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1131 = incrWrite ? _GEN_363 : memReg_13_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1132 = incrWrite ? _GEN_364 : memReg_14_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1133 = incrWrite ? _GEN_365 : memReg_15_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1134 = incrWrite ? _GEN_366 : memReg_16_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1135 = incrWrite ? _GEN_367 : memReg_17_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1136 = incrWrite ? _GEN_368 : memReg_18_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1137 = incrWrite ? _GEN_369 : memReg_19_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1138 = incrWrite ? _GEN_370 : memReg_20_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1139 = incrWrite ? _GEN_371 : memReg_21_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1140 = incrWrite ? _GEN_372 : memReg_22_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1141 = incrWrite ? _GEN_373 : memReg_23_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1142 = incrWrite ? _GEN_374 : memReg_24_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1143 = incrWrite ? _GEN_375 : memReg_25_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1144 = incrWrite ? _GEN_376 : memReg_26_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1145 = incrWrite ? _GEN_377 : memReg_27_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1146 = incrWrite ? _GEN_378 : memReg_28_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1147 = incrWrite ? _GEN_379 : memReg_29_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1148 = incrWrite ? _GEN_380 : memReg_30_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1149 = incrWrite ? _GEN_381 : memReg_31_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1150 = incrWrite ? _GEN_382 : memReg_32_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1151 = incrWrite ? _GEN_383 : memReg_33_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1152 = incrWrite ? _GEN_384 : memReg_34_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1153 = incrWrite ? _GEN_385 : memReg_35_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1154 = incrWrite ? _GEN_386 : memReg_36_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1155 = incrWrite ? _GEN_387 : memReg_37_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1156 = incrWrite ? _GEN_388 : memReg_38_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1157 = incrWrite ? _GEN_389 : memReg_39_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1158 = incrWrite ? _GEN_390 : memReg_40_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1159 = incrWrite ? _GEN_391 : memReg_41_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1160 = incrWrite ? _GEN_392 : memReg_42_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1161 = incrWrite ? _GEN_393 : memReg_43_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1162 = incrWrite ? _GEN_394 : memReg_44_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1163 = incrWrite ? _GEN_395 : memReg_45_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1164 = incrWrite ? _GEN_396 : memReg_46_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1165 = incrWrite ? _GEN_397 : memReg_47_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1166 = incrWrite ? _GEN_398 : memReg_48_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1167 = incrWrite ? _GEN_399 : memReg_49_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1168 = incrWrite ? _GEN_400 : memReg_50_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1169 = incrWrite ? _GEN_401 : memReg_51_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1170 = incrWrite ? _GEN_402 : memReg_52_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1171 = incrWrite ? _GEN_403 : memReg_53_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1172 = incrWrite ? _GEN_404 : memReg_54_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1173 = incrWrite ? _GEN_405 : memReg_55_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1174 = incrWrite ? _GEN_406 : memReg_56_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1175 = incrWrite ? _GEN_407 : memReg_57_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1176 = incrWrite ? _GEN_408 : memReg_58_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1177 = incrWrite ? _GEN_409 : memReg_59_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1178 = incrWrite ? _GEN_410 : memReg_60_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1179 = incrWrite ? _GEN_411 : memReg_61_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1180 = incrWrite ? _GEN_412 : memReg_62_branch_valid; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1181 = incrWrite ? _GEN_413 : memReg_63_branch_valid; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1182 = incrWrite ? _GEN_414 : memReg_0_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1183 = incrWrite ? _GEN_415 : memReg_1_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1184 = incrWrite ? _GEN_416 : memReg_2_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1185 = incrWrite ? _GEN_417 : memReg_3_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1186 = incrWrite ? _GEN_418 : memReg_4_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1187 = incrWrite ? _GEN_419 : memReg_5_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1188 = incrWrite ? _GEN_420 : memReg_6_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1189 = incrWrite ? _GEN_421 : memReg_7_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1190 = incrWrite ? _GEN_422 : memReg_8_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1191 = incrWrite ? _GEN_423 : memReg_9_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1192 = incrWrite ? _GEN_424 : memReg_10_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1193 = incrWrite ? _GEN_425 : memReg_11_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1194 = incrWrite ? _GEN_426 : memReg_12_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1195 = incrWrite ? _GEN_427 : memReg_13_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1196 = incrWrite ? _GEN_428 : memReg_14_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1197 = incrWrite ? _GEN_429 : memReg_15_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1198 = incrWrite ? _GEN_430 : memReg_16_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1199 = incrWrite ? _GEN_431 : memReg_17_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1200 = incrWrite ? _GEN_432 : memReg_18_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1201 = incrWrite ? _GEN_433 : memReg_19_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1202 = incrWrite ? _GEN_434 : memReg_20_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1203 = incrWrite ? _GEN_435 : memReg_21_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1204 = incrWrite ? _GEN_436 : memReg_22_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1205 = incrWrite ? _GEN_437 : memReg_23_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1206 = incrWrite ? _GEN_438 : memReg_24_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1207 = incrWrite ? _GEN_439 : memReg_25_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1208 = incrWrite ? _GEN_440 : memReg_26_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1209 = incrWrite ? _GEN_441 : memReg_27_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1210 = incrWrite ? _GEN_442 : memReg_28_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1211 = incrWrite ? _GEN_443 : memReg_29_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1212 = incrWrite ? _GEN_444 : memReg_30_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1213 = incrWrite ? _GEN_445 : memReg_31_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1214 = incrWrite ? _GEN_446 : memReg_32_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1215 = incrWrite ? _GEN_447 : memReg_33_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1216 = incrWrite ? _GEN_448 : memReg_34_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1217 = incrWrite ? _GEN_449 : memReg_35_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1218 = incrWrite ? _GEN_450 : memReg_36_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1219 = incrWrite ? _GEN_451 : memReg_37_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1220 = incrWrite ? _GEN_452 : memReg_38_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1221 = incrWrite ? _GEN_453 : memReg_39_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1222 = incrWrite ? _GEN_454 : memReg_40_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1223 = incrWrite ? _GEN_455 : memReg_41_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1224 = incrWrite ? _GEN_456 : memReg_42_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1225 = incrWrite ? _GEN_457 : memReg_43_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1226 = incrWrite ? _GEN_458 : memReg_44_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1227 = incrWrite ? _GEN_459 : memReg_45_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1228 = incrWrite ? _GEN_460 : memReg_46_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1229 = incrWrite ? _GEN_461 : memReg_47_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1230 = incrWrite ? _GEN_462 : memReg_48_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1231 = incrWrite ? _GEN_463 : memReg_49_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1232 = incrWrite ? _GEN_464 : memReg_50_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1233 = incrWrite ? _GEN_465 : memReg_51_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1234 = incrWrite ? _GEN_466 : memReg_52_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1235 = incrWrite ? _GEN_467 : memReg_53_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1236 = incrWrite ? _GEN_468 : memReg_54_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1237 = incrWrite ? _GEN_469 : memReg_55_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1238 = incrWrite ? _GEN_470 : memReg_56_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1239 = incrWrite ? _GEN_471 : memReg_57_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1240 = incrWrite ? _GEN_472 : memReg_58_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1241 = incrWrite ? _GEN_473 : memReg_59_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1242 = incrWrite ? _GEN_474 : memReg_60_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1243 = incrWrite ? _GEN_475 : memReg_61_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1244 = incrWrite ? _GEN_476 : memReg_62_branch_mask; // @[fifo.scala 81:17 27:33]
  wire [4:0] _GEN_1245 = incrWrite ? _GEN_477 : memReg_63_branch_mask; // @[fifo.scala 81:17 27:33]
  wire  _GEN_1567 = 6'h1 == readPtr ? memReg_1_valid : memReg_0_valid; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1568 = 6'h2 == readPtr ? memReg_2_valid : _GEN_1567; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1569 = 6'h3 == readPtr ? memReg_3_valid : _GEN_1568; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1570 = 6'h4 == readPtr ? memReg_4_valid : _GEN_1569; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1571 = 6'h5 == readPtr ? memReg_5_valid : _GEN_1570; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1572 = 6'h6 == readPtr ? memReg_6_valid : _GEN_1571; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1573 = 6'h7 == readPtr ? memReg_7_valid : _GEN_1572; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1574 = 6'h8 == readPtr ? memReg_8_valid : _GEN_1573; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1575 = 6'h9 == readPtr ? memReg_9_valid : _GEN_1574; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1576 = 6'ha == readPtr ? memReg_10_valid : _GEN_1575; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1577 = 6'hb == readPtr ? memReg_11_valid : _GEN_1576; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1578 = 6'hc == readPtr ? memReg_12_valid : _GEN_1577; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1579 = 6'hd == readPtr ? memReg_13_valid : _GEN_1578; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1580 = 6'he == readPtr ? memReg_14_valid : _GEN_1579; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1581 = 6'hf == readPtr ? memReg_15_valid : _GEN_1580; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1582 = 6'h10 == readPtr ? memReg_16_valid : _GEN_1581; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1583 = 6'h11 == readPtr ? memReg_17_valid : _GEN_1582; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1584 = 6'h12 == readPtr ? memReg_18_valid : _GEN_1583; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1585 = 6'h13 == readPtr ? memReg_19_valid : _GEN_1584; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1586 = 6'h14 == readPtr ? memReg_20_valid : _GEN_1585; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1587 = 6'h15 == readPtr ? memReg_21_valid : _GEN_1586; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1588 = 6'h16 == readPtr ? memReg_22_valid : _GEN_1587; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1589 = 6'h17 == readPtr ? memReg_23_valid : _GEN_1588; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1590 = 6'h18 == readPtr ? memReg_24_valid : _GEN_1589; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1591 = 6'h19 == readPtr ? memReg_25_valid : _GEN_1590; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1592 = 6'h1a == readPtr ? memReg_26_valid : _GEN_1591; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1593 = 6'h1b == readPtr ? memReg_27_valid : _GEN_1592; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1594 = 6'h1c == readPtr ? memReg_28_valid : _GEN_1593; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1595 = 6'h1d == readPtr ? memReg_29_valid : _GEN_1594; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1596 = 6'h1e == readPtr ? memReg_30_valid : _GEN_1595; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1597 = 6'h1f == readPtr ? memReg_31_valid : _GEN_1596; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1598 = 6'h20 == readPtr ? memReg_32_valid : _GEN_1597; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1599 = 6'h21 == readPtr ? memReg_33_valid : _GEN_1598; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1600 = 6'h22 == readPtr ? memReg_34_valid : _GEN_1599; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1601 = 6'h23 == readPtr ? memReg_35_valid : _GEN_1600; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1602 = 6'h24 == readPtr ? memReg_36_valid : _GEN_1601; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1603 = 6'h25 == readPtr ? memReg_37_valid : _GEN_1602; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1604 = 6'h26 == readPtr ? memReg_38_valid : _GEN_1603; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1605 = 6'h27 == readPtr ? memReg_39_valid : _GEN_1604; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1606 = 6'h28 == readPtr ? memReg_40_valid : _GEN_1605; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1607 = 6'h29 == readPtr ? memReg_41_valid : _GEN_1606; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1608 = 6'h2a == readPtr ? memReg_42_valid : _GEN_1607; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1609 = 6'h2b == readPtr ? memReg_43_valid : _GEN_1608; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1610 = 6'h2c == readPtr ? memReg_44_valid : _GEN_1609; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1611 = 6'h2d == readPtr ? memReg_45_valid : _GEN_1610; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1612 = 6'h2e == readPtr ? memReg_46_valid : _GEN_1611; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1613 = 6'h2f == readPtr ? memReg_47_valid : _GEN_1612; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1614 = 6'h30 == readPtr ? memReg_48_valid : _GEN_1613; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1615 = 6'h31 == readPtr ? memReg_49_valid : _GEN_1614; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1616 = 6'h32 == readPtr ? memReg_50_valid : _GEN_1615; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1617 = 6'h33 == readPtr ? memReg_51_valid : _GEN_1616; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1618 = 6'h34 == readPtr ? memReg_52_valid : _GEN_1617; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1619 = 6'h35 == readPtr ? memReg_53_valid : _GEN_1618; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1620 = 6'h36 == readPtr ? memReg_54_valid : _GEN_1619; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1621 = 6'h37 == readPtr ? memReg_55_valid : _GEN_1620; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1622 = 6'h38 == readPtr ? memReg_56_valid : _GEN_1621; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1623 = 6'h39 == readPtr ? memReg_57_valid : _GEN_1622; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1624 = 6'h3a == readPtr ? memReg_58_valid : _GEN_1623; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1625 = 6'h3b == readPtr ? memReg_59_valid : _GEN_1624; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1626 = 6'h3c == readPtr ? memReg_60_valid : _GEN_1625; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1627 = 6'h3d == readPtr ? memReg_61_valid : _GEN_1626; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1628 = 6'h3e == readPtr ? memReg_62_valid : _GEN_1627; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1629 = 6'h3f == readPtr ? memReg_63_valid : _GEN_1628; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1887 = 6'h1 == readPtr ? memReg_1_branch_valid : memReg_0_branch_valid; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1888 = 6'h2 == readPtr ? memReg_2_branch_valid : _GEN_1887; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1889 = 6'h3 == readPtr ? memReg_3_branch_valid : _GEN_1888; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1890 = 6'h4 == readPtr ? memReg_4_branch_valid : _GEN_1889; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1891 = 6'h5 == readPtr ? memReg_5_branch_valid : _GEN_1890; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1892 = 6'h6 == readPtr ? memReg_6_branch_valid : _GEN_1891; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1893 = 6'h7 == readPtr ? memReg_7_branch_valid : _GEN_1892; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1894 = 6'h8 == readPtr ? memReg_8_branch_valid : _GEN_1893; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1895 = 6'h9 == readPtr ? memReg_9_branch_valid : _GEN_1894; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1896 = 6'ha == readPtr ? memReg_10_branch_valid : _GEN_1895; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1897 = 6'hb == readPtr ? memReg_11_branch_valid : _GEN_1896; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1898 = 6'hc == readPtr ? memReg_12_branch_valid : _GEN_1897; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1899 = 6'hd == readPtr ? memReg_13_branch_valid : _GEN_1898; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1900 = 6'he == readPtr ? memReg_14_branch_valid : _GEN_1899; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1901 = 6'hf == readPtr ? memReg_15_branch_valid : _GEN_1900; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1902 = 6'h10 == readPtr ? memReg_16_branch_valid : _GEN_1901; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1903 = 6'h11 == readPtr ? memReg_17_branch_valid : _GEN_1902; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1904 = 6'h12 == readPtr ? memReg_18_branch_valid : _GEN_1903; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1905 = 6'h13 == readPtr ? memReg_19_branch_valid : _GEN_1904; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1906 = 6'h14 == readPtr ? memReg_20_branch_valid : _GEN_1905; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1907 = 6'h15 == readPtr ? memReg_21_branch_valid : _GEN_1906; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1908 = 6'h16 == readPtr ? memReg_22_branch_valid : _GEN_1907; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1909 = 6'h17 == readPtr ? memReg_23_branch_valid : _GEN_1908; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1910 = 6'h18 == readPtr ? memReg_24_branch_valid : _GEN_1909; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1911 = 6'h19 == readPtr ? memReg_25_branch_valid : _GEN_1910; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1912 = 6'h1a == readPtr ? memReg_26_branch_valid : _GEN_1911; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1913 = 6'h1b == readPtr ? memReg_27_branch_valid : _GEN_1912; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1914 = 6'h1c == readPtr ? memReg_28_branch_valid : _GEN_1913; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1915 = 6'h1d == readPtr ? memReg_29_branch_valid : _GEN_1914; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1916 = 6'h1e == readPtr ? memReg_30_branch_valid : _GEN_1915; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1917 = 6'h1f == readPtr ? memReg_31_branch_valid : _GEN_1916; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1918 = 6'h20 == readPtr ? memReg_32_branch_valid : _GEN_1917; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1919 = 6'h21 == readPtr ? memReg_33_branch_valid : _GEN_1918; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1920 = 6'h22 == readPtr ? memReg_34_branch_valid : _GEN_1919; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1921 = 6'h23 == readPtr ? memReg_35_branch_valid : _GEN_1920; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1922 = 6'h24 == readPtr ? memReg_36_branch_valid : _GEN_1921; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1923 = 6'h25 == readPtr ? memReg_37_branch_valid : _GEN_1922; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1924 = 6'h26 == readPtr ? memReg_38_branch_valid : _GEN_1923; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1925 = 6'h27 == readPtr ? memReg_39_branch_valid : _GEN_1924; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1926 = 6'h28 == readPtr ? memReg_40_branch_valid : _GEN_1925; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1927 = 6'h29 == readPtr ? memReg_41_branch_valid : _GEN_1926; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1928 = 6'h2a == readPtr ? memReg_42_branch_valid : _GEN_1927; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1929 = 6'h2b == readPtr ? memReg_43_branch_valid : _GEN_1928; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1930 = 6'h2c == readPtr ? memReg_44_branch_valid : _GEN_1929; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1931 = 6'h2d == readPtr ? memReg_45_branch_valid : _GEN_1930; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1932 = 6'h2e == readPtr ? memReg_46_branch_valid : _GEN_1931; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1933 = 6'h2f == readPtr ? memReg_47_branch_valid : _GEN_1932; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1934 = 6'h30 == readPtr ? memReg_48_branch_valid : _GEN_1933; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1935 = 6'h31 == readPtr ? memReg_49_branch_valid : _GEN_1934; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1936 = 6'h32 == readPtr ? memReg_50_branch_valid : _GEN_1935; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1937 = 6'h33 == readPtr ? memReg_51_branch_valid : _GEN_1936; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1938 = 6'h34 == readPtr ? memReg_52_branch_valid : _GEN_1937; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1939 = 6'h35 == readPtr ? memReg_53_branch_valid : _GEN_1938; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1940 = 6'h36 == readPtr ? memReg_54_branch_valid : _GEN_1939; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1941 = 6'h37 == readPtr ? memReg_55_branch_valid : _GEN_1940; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1942 = 6'h38 == readPtr ? memReg_56_branch_valid : _GEN_1941; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1943 = 6'h39 == readPtr ? memReg_57_branch_valid : _GEN_1942; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1944 = 6'h3a == readPtr ? memReg_58_branch_valid : _GEN_1943; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1945 = 6'h3b == readPtr ? memReg_59_branch_valid : _GEN_1944; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1946 = 6'h3c == readPtr ? memReg_60_branch_valid : _GEN_1945; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1947 = 6'h3d == readPtr ? memReg_61_branch_valid : _GEN_1946; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1948 = 6'h3e == readPtr ? memReg_62_branch_valid : _GEN_1947; // @[fifo.scala 86:{13,13}]
  wire  _GEN_1949 = 6'h3f == readPtr ? memReg_63_branch_valid : _GEN_1948; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1951 = 6'h1 == readPtr ? memReg_1_branch_mask : memReg_0_branch_mask; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1952 = 6'h2 == readPtr ? memReg_2_branch_mask : _GEN_1951; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1953 = 6'h3 == readPtr ? memReg_3_branch_mask : _GEN_1952; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1954 = 6'h4 == readPtr ? memReg_4_branch_mask : _GEN_1953; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1955 = 6'h5 == readPtr ? memReg_5_branch_mask : _GEN_1954; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1956 = 6'h6 == readPtr ? memReg_6_branch_mask : _GEN_1955; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1957 = 6'h7 == readPtr ? memReg_7_branch_mask : _GEN_1956; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1958 = 6'h8 == readPtr ? memReg_8_branch_mask : _GEN_1957; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1959 = 6'h9 == readPtr ? memReg_9_branch_mask : _GEN_1958; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1960 = 6'ha == readPtr ? memReg_10_branch_mask : _GEN_1959; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1961 = 6'hb == readPtr ? memReg_11_branch_mask : _GEN_1960; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1962 = 6'hc == readPtr ? memReg_12_branch_mask : _GEN_1961; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1963 = 6'hd == readPtr ? memReg_13_branch_mask : _GEN_1962; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1964 = 6'he == readPtr ? memReg_14_branch_mask : _GEN_1963; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1965 = 6'hf == readPtr ? memReg_15_branch_mask : _GEN_1964; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1966 = 6'h10 == readPtr ? memReg_16_branch_mask : _GEN_1965; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1967 = 6'h11 == readPtr ? memReg_17_branch_mask : _GEN_1966; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1968 = 6'h12 == readPtr ? memReg_18_branch_mask : _GEN_1967; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1969 = 6'h13 == readPtr ? memReg_19_branch_mask : _GEN_1968; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1970 = 6'h14 == readPtr ? memReg_20_branch_mask : _GEN_1969; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1971 = 6'h15 == readPtr ? memReg_21_branch_mask : _GEN_1970; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1972 = 6'h16 == readPtr ? memReg_22_branch_mask : _GEN_1971; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1973 = 6'h17 == readPtr ? memReg_23_branch_mask : _GEN_1972; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1974 = 6'h18 == readPtr ? memReg_24_branch_mask : _GEN_1973; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1975 = 6'h19 == readPtr ? memReg_25_branch_mask : _GEN_1974; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1976 = 6'h1a == readPtr ? memReg_26_branch_mask : _GEN_1975; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1977 = 6'h1b == readPtr ? memReg_27_branch_mask : _GEN_1976; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1978 = 6'h1c == readPtr ? memReg_28_branch_mask : _GEN_1977; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1979 = 6'h1d == readPtr ? memReg_29_branch_mask : _GEN_1978; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1980 = 6'h1e == readPtr ? memReg_30_branch_mask : _GEN_1979; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1981 = 6'h1f == readPtr ? memReg_31_branch_mask : _GEN_1980; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1982 = 6'h20 == readPtr ? memReg_32_branch_mask : _GEN_1981; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1983 = 6'h21 == readPtr ? memReg_33_branch_mask : _GEN_1982; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1984 = 6'h22 == readPtr ? memReg_34_branch_mask : _GEN_1983; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1985 = 6'h23 == readPtr ? memReg_35_branch_mask : _GEN_1984; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1986 = 6'h24 == readPtr ? memReg_36_branch_mask : _GEN_1985; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1987 = 6'h25 == readPtr ? memReg_37_branch_mask : _GEN_1986; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1988 = 6'h26 == readPtr ? memReg_38_branch_mask : _GEN_1987; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1989 = 6'h27 == readPtr ? memReg_39_branch_mask : _GEN_1988; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1990 = 6'h28 == readPtr ? memReg_40_branch_mask : _GEN_1989; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1991 = 6'h29 == readPtr ? memReg_41_branch_mask : _GEN_1990; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1992 = 6'h2a == readPtr ? memReg_42_branch_mask : _GEN_1991; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1993 = 6'h2b == readPtr ? memReg_43_branch_mask : _GEN_1992; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1994 = 6'h2c == readPtr ? memReg_44_branch_mask : _GEN_1993; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1995 = 6'h2d == readPtr ? memReg_45_branch_mask : _GEN_1994; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1996 = 6'h2e == readPtr ? memReg_46_branch_mask : _GEN_1995; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1997 = 6'h2f == readPtr ? memReg_47_branch_mask : _GEN_1996; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1998 = 6'h30 == readPtr ? memReg_48_branch_mask : _GEN_1997; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_1999 = 6'h31 == readPtr ? memReg_49_branch_mask : _GEN_1998; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_2000 = 6'h32 == readPtr ? memReg_50_branch_mask : _GEN_1999; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_2001 = 6'h33 == readPtr ? memReg_51_branch_mask : _GEN_2000; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_2002 = 6'h34 == readPtr ? memReg_52_branch_mask : _GEN_2001; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_2003 = 6'h35 == readPtr ? memReg_53_branch_mask : _GEN_2002; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_2004 = 6'h36 == readPtr ? memReg_54_branch_mask : _GEN_2003; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_2005 = 6'h37 == readPtr ? memReg_55_branch_mask : _GEN_2004; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_2006 = 6'h38 == readPtr ? memReg_56_branch_mask : _GEN_2005; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_2007 = 6'h39 == readPtr ? memReg_57_branch_mask : _GEN_2006; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_2008 = 6'h3a == readPtr ? memReg_58_branch_mask : _GEN_2007; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_2009 = 6'h3b == readPtr ? memReg_59_branch_mask : _GEN_2008; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_2010 = 6'h3c == readPtr ? memReg_60_branch_mask : _GEN_2009; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_2011 = 6'h3d == readPtr ? memReg_61_branch_mask : _GEN_2010; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_2012 = 6'h3e == readPtr ? memReg_62_branch_mask : _GEN_2011; // @[fifo.scala 86:{13,13}]
  wire [4:0] _GEN_2013 = 6'h3f == readPtr ? memReg_63_branch_mask : _GEN_2012; // @[fifo.scala 86:{13,13}]
  wire [4:0] _T_8 = write_data_branch_mask & branchOps_branchMask; // @[utils.scala 62:31]
  wire  _T_9 = |_T_8; // @[utils.scala 62:55]
  wire [4:0] _memReg_branch_mask_T = write_data_branch_mask ^ branchOps_branchMask; // @[utils.scala 63:42]
  wire [4:0] _GEN_2334 = 6'h0 == writePtr ? _memReg_branch_mask_T : _GEN_1182; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2335 = 6'h1 == writePtr ? _memReg_branch_mask_T : _GEN_1183; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2336 = 6'h2 == writePtr ? _memReg_branch_mask_T : _GEN_1184; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2337 = 6'h3 == writePtr ? _memReg_branch_mask_T : _GEN_1185; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2338 = 6'h4 == writePtr ? _memReg_branch_mask_T : _GEN_1186; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2339 = 6'h5 == writePtr ? _memReg_branch_mask_T : _GEN_1187; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2340 = 6'h6 == writePtr ? _memReg_branch_mask_T : _GEN_1188; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2341 = 6'h7 == writePtr ? _memReg_branch_mask_T : _GEN_1189; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2342 = 6'h8 == writePtr ? _memReg_branch_mask_T : _GEN_1190; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2343 = 6'h9 == writePtr ? _memReg_branch_mask_T : _GEN_1191; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2344 = 6'ha == writePtr ? _memReg_branch_mask_T : _GEN_1192; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2345 = 6'hb == writePtr ? _memReg_branch_mask_T : _GEN_1193; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2346 = 6'hc == writePtr ? _memReg_branch_mask_T : _GEN_1194; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2347 = 6'hd == writePtr ? _memReg_branch_mask_T : _GEN_1195; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2348 = 6'he == writePtr ? _memReg_branch_mask_T : _GEN_1196; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2349 = 6'hf == writePtr ? _memReg_branch_mask_T : _GEN_1197; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2350 = 6'h10 == writePtr ? _memReg_branch_mask_T : _GEN_1198; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2351 = 6'h11 == writePtr ? _memReg_branch_mask_T : _GEN_1199; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2352 = 6'h12 == writePtr ? _memReg_branch_mask_T : _GEN_1200; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2353 = 6'h13 == writePtr ? _memReg_branch_mask_T : _GEN_1201; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2354 = 6'h14 == writePtr ? _memReg_branch_mask_T : _GEN_1202; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2355 = 6'h15 == writePtr ? _memReg_branch_mask_T : _GEN_1203; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2356 = 6'h16 == writePtr ? _memReg_branch_mask_T : _GEN_1204; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2357 = 6'h17 == writePtr ? _memReg_branch_mask_T : _GEN_1205; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2358 = 6'h18 == writePtr ? _memReg_branch_mask_T : _GEN_1206; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2359 = 6'h19 == writePtr ? _memReg_branch_mask_T : _GEN_1207; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2360 = 6'h1a == writePtr ? _memReg_branch_mask_T : _GEN_1208; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2361 = 6'h1b == writePtr ? _memReg_branch_mask_T : _GEN_1209; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2362 = 6'h1c == writePtr ? _memReg_branch_mask_T : _GEN_1210; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2363 = 6'h1d == writePtr ? _memReg_branch_mask_T : _GEN_1211; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2364 = 6'h1e == writePtr ? _memReg_branch_mask_T : _GEN_1212; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2365 = 6'h1f == writePtr ? _memReg_branch_mask_T : _GEN_1213; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2366 = 6'h20 == writePtr ? _memReg_branch_mask_T : _GEN_1214; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2367 = 6'h21 == writePtr ? _memReg_branch_mask_T : _GEN_1215; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2368 = 6'h22 == writePtr ? _memReg_branch_mask_T : _GEN_1216; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2369 = 6'h23 == writePtr ? _memReg_branch_mask_T : _GEN_1217; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2370 = 6'h24 == writePtr ? _memReg_branch_mask_T : _GEN_1218; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2371 = 6'h25 == writePtr ? _memReg_branch_mask_T : _GEN_1219; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2372 = 6'h26 == writePtr ? _memReg_branch_mask_T : _GEN_1220; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2373 = 6'h27 == writePtr ? _memReg_branch_mask_T : _GEN_1221; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2374 = 6'h28 == writePtr ? _memReg_branch_mask_T : _GEN_1222; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2375 = 6'h29 == writePtr ? _memReg_branch_mask_T : _GEN_1223; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2376 = 6'h2a == writePtr ? _memReg_branch_mask_T : _GEN_1224; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2377 = 6'h2b == writePtr ? _memReg_branch_mask_T : _GEN_1225; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2378 = 6'h2c == writePtr ? _memReg_branch_mask_T : _GEN_1226; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2379 = 6'h2d == writePtr ? _memReg_branch_mask_T : _GEN_1227; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2380 = 6'h2e == writePtr ? _memReg_branch_mask_T : _GEN_1228; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2381 = 6'h2f == writePtr ? _memReg_branch_mask_T : _GEN_1229; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2382 = 6'h30 == writePtr ? _memReg_branch_mask_T : _GEN_1230; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2383 = 6'h31 == writePtr ? _memReg_branch_mask_T : _GEN_1231; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2384 = 6'h32 == writePtr ? _memReg_branch_mask_T : _GEN_1232; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2385 = 6'h33 == writePtr ? _memReg_branch_mask_T : _GEN_1233; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2386 = 6'h34 == writePtr ? _memReg_branch_mask_T : _GEN_1234; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2387 = 6'h35 == writePtr ? _memReg_branch_mask_T : _GEN_1235; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2388 = 6'h36 == writePtr ? _memReg_branch_mask_T : _GEN_1236; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2389 = 6'h37 == writePtr ? _memReg_branch_mask_T : _GEN_1237; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2390 = 6'h38 == writePtr ? _memReg_branch_mask_T : _GEN_1238; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2391 = 6'h39 == writePtr ? _memReg_branch_mask_T : _GEN_1239; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2392 = 6'h3a == writePtr ? _memReg_branch_mask_T : _GEN_1240; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2393 = 6'h3b == writePtr ? _memReg_branch_mask_T : _GEN_1241; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2394 = 6'h3c == writePtr ? _memReg_branch_mask_T : _GEN_1242; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2395 = 6'h3d == writePtr ? _memReg_branch_mask_T : _GEN_1243; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2396 = 6'h3e == writePtr ? _memReg_branch_mask_T : _GEN_1244; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2397 = 6'h3f == writePtr ? _memReg_branch_mask_T : _GEN_1245; // @[utils.scala 63:{23,23}]
  wire [4:0] _GEN_2398 = 6'h0 == writePtr ? write_data_branch_mask : _GEN_1182; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2399 = 6'h1 == writePtr ? write_data_branch_mask : _GEN_1183; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2400 = 6'h2 == writePtr ? write_data_branch_mask : _GEN_1184; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2401 = 6'h3 == writePtr ? write_data_branch_mask : _GEN_1185; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2402 = 6'h4 == writePtr ? write_data_branch_mask : _GEN_1186; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2403 = 6'h5 == writePtr ? write_data_branch_mask : _GEN_1187; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2404 = 6'h6 == writePtr ? write_data_branch_mask : _GEN_1188; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2405 = 6'h7 == writePtr ? write_data_branch_mask : _GEN_1189; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2406 = 6'h8 == writePtr ? write_data_branch_mask : _GEN_1190; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2407 = 6'h9 == writePtr ? write_data_branch_mask : _GEN_1191; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2408 = 6'ha == writePtr ? write_data_branch_mask : _GEN_1192; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2409 = 6'hb == writePtr ? write_data_branch_mask : _GEN_1193; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2410 = 6'hc == writePtr ? write_data_branch_mask : _GEN_1194; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2411 = 6'hd == writePtr ? write_data_branch_mask : _GEN_1195; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2412 = 6'he == writePtr ? write_data_branch_mask : _GEN_1196; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2413 = 6'hf == writePtr ? write_data_branch_mask : _GEN_1197; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2414 = 6'h10 == writePtr ? write_data_branch_mask : _GEN_1198; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2415 = 6'h11 == writePtr ? write_data_branch_mask : _GEN_1199; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2416 = 6'h12 == writePtr ? write_data_branch_mask : _GEN_1200; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2417 = 6'h13 == writePtr ? write_data_branch_mask : _GEN_1201; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2418 = 6'h14 == writePtr ? write_data_branch_mask : _GEN_1202; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2419 = 6'h15 == writePtr ? write_data_branch_mask : _GEN_1203; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2420 = 6'h16 == writePtr ? write_data_branch_mask : _GEN_1204; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2421 = 6'h17 == writePtr ? write_data_branch_mask : _GEN_1205; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2422 = 6'h18 == writePtr ? write_data_branch_mask : _GEN_1206; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2423 = 6'h19 == writePtr ? write_data_branch_mask : _GEN_1207; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2424 = 6'h1a == writePtr ? write_data_branch_mask : _GEN_1208; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2425 = 6'h1b == writePtr ? write_data_branch_mask : _GEN_1209; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2426 = 6'h1c == writePtr ? write_data_branch_mask : _GEN_1210; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2427 = 6'h1d == writePtr ? write_data_branch_mask : _GEN_1211; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2428 = 6'h1e == writePtr ? write_data_branch_mask : _GEN_1212; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2429 = 6'h1f == writePtr ? write_data_branch_mask : _GEN_1213; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2430 = 6'h20 == writePtr ? write_data_branch_mask : _GEN_1214; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2431 = 6'h21 == writePtr ? write_data_branch_mask : _GEN_1215; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2432 = 6'h22 == writePtr ? write_data_branch_mask : _GEN_1216; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2433 = 6'h23 == writePtr ? write_data_branch_mask : _GEN_1217; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2434 = 6'h24 == writePtr ? write_data_branch_mask : _GEN_1218; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2435 = 6'h25 == writePtr ? write_data_branch_mask : _GEN_1219; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2436 = 6'h26 == writePtr ? write_data_branch_mask : _GEN_1220; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2437 = 6'h27 == writePtr ? write_data_branch_mask : _GEN_1221; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2438 = 6'h28 == writePtr ? write_data_branch_mask : _GEN_1222; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2439 = 6'h29 == writePtr ? write_data_branch_mask : _GEN_1223; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2440 = 6'h2a == writePtr ? write_data_branch_mask : _GEN_1224; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2441 = 6'h2b == writePtr ? write_data_branch_mask : _GEN_1225; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2442 = 6'h2c == writePtr ? write_data_branch_mask : _GEN_1226; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2443 = 6'h2d == writePtr ? write_data_branch_mask : _GEN_1227; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2444 = 6'h2e == writePtr ? write_data_branch_mask : _GEN_1228; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2445 = 6'h2f == writePtr ? write_data_branch_mask : _GEN_1229; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2446 = 6'h30 == writePtr ? write_data_branch_mask : _GEN_1230; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2447 = 6'h31 == writePtr ? write_data_branch_mask : _GEN_1231; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2448 = 6'h32 == writePtr ? write_data_branch_mask : _GEN_1232; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2449 = 6'h33 == writePtr ? write_data_branch_mask : _GEN_1233; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2450 = 6'h34 == writePtr ? write_data_branch_mask : _GEN_1234; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2451 = 6'h35 == writePtr ? write_data_branch_mask : _GEN_1235; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2452 = 6'h36 == writePtr ? write_data_branch_mask : _GEN_1236; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2453 = 6'h37 == writePtr ? write_data_branch_mask : _GEN_1237; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2454 = 6'h38 == writePtr ? write_data_branch_mask : _GEN_1238; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2455 = 6'h39 == writePtr ? write_data_branch_mask : _GEN_1239; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2456 = 6'h3a == writePtr ? write_data_branch_mask : _GEN_1240; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2457 = 6'h3b == writePtr ? write_data_branch_mask : _GEN_1241; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2458 = 6'h3c == writePtr ? write_data_branch_mask : _GEN_1242; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2459 = 6'h3d == writePtr ? write_data_branch_mask : _GEN_1243; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2460 = 6'h3e == writePtr ? write_data_branch_mask : _GEN_1244; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2461 = 6'h3f == writePtr ? write_data_branch_mask : _GEN_1245; // @[utils.scala 65:{23,23}]
  wire [4:0] _GEN_2462 = |_T_8 ? _GEN_2334 : _GEN_2398; // @[utils.scala 62:60]
  wire [4:0] _GEN_2463 = |_T_8 ? _GEN_2335 : _GEN_2399; // @[utils.scala 62:60]
  wire [4:0] _GEN_2464 = |_T_8 ? _GEN_2336 : _GEN_2400; // @[utils.scala 62:60]
  wire [4:0] _GEN_2465 = |_T_8 ? _GEN_2337 : _GEN_2401; // @[utils.scala 62:60]
  wire [4:0] _GEN_2466 = |_T_8 ? _GEN_2338 : _GEN_2402; // @[utils.scala 62:60]
  wire [4:0] _GEN_2467 = |_T_8 ? _GEN_2339 : _GEN_2403; // @[utils.scala 62:60]
  wire [4:0] _GEN_2468 = |_T_8 ? _GEN_2340 : _GEN_2404; // @[utils.scala 62:60]
  wire [4:0] _GEN_2469 = |_T_8 ? _GEN_2341 : _GEN_2405; // @[utils.scala 62:60]
  wire [4:0] _GEN_2470 = |_T_8 ? _GEN_2342 : _GEN_2406; // @[utils.scala 62:60]
  wire [4:0] _GEN_2471 = |_T_8 ? _GEN_2343 : _GEN_2407; // @[utils.scala 62:60]
  wire [4:0] _GEN_2472 = |_T_8 ? _GEN_2344 : _GEN_2408; // @[utils.scala 62:60]
  wire [4:0] _GEN_2473 = |_T_8 ? _GEN_2345 : _GEN_2409; // @[utils.scala 62:60]
  wire [4:0] _GEN_2474 = |_T_8 ? _GEN_2346 : _GEN_2410; // @[utils.scala 62:60]
  wire [4:0] _GEN_2475 = |_T_8 ? _GEN_2347 : _GEN_2411; // @[utils.scala 62:60]
  wire [4:0] _GEN_2476 = |_T_8 ? _GEN_2348 : _GEN_2412; // @[utils.scala 62:60]
  wire [4:0] _GEN_2477 = |_T_8 ? _GEN_2349 : _GEN_2413; // @[utils.scala 62:60]
  wire [4:0] _GEN_2478 = |_T_8 ? _GEN_2350 : _GEN_2414; // @[utils.scala 62:60]
  wire [4:0] _GEN_2479 = |_T_8 ? _GEN_2351 : _GEN_2415; // @[utils.scala 62:60]
  wire [4:0] _GEN_2480 = |_T_8 ? _GEN_2352 : _GEN_2416; // @[utils.scala 62:60]
  wire [4:0] _GEN_2481 = |_T_8 ? _GEN_2353 : _GEN_2417; // @[utils.scala 62:60]
  wire [4:0] _GEN_2482 = |_T_8 ? _GEN_2354 : _GEN_2418; // @[utils.scala 62:60]
  wire [4:0] _GEN_2483 = |_T_8 ? _GEN_2355 : _GEN_2419; // @[utils.scala 62:60]
  wire [4:0] _GEN_2484 = |_T_8 ? _GEN_2356 : _GEN_2420; // @[utils.scala 62:60]
  wire [4:0] _GEN_2485 = |_T_8 ? _GEN_2357 : _GEN_2421; // @[utils.scala 62:60]
  wire [4:0] _GEN_2486 = |_T_8 ? _GEN_2358 : _GEN_2422; // @[utils.scala 62:60]
  wire [4:0] _GEN_2487 = |_T_8 ? _GEN_2359 : _GEN_2423; // @[utils.scala 62:60]
  wire [4:0] _GEN_2488 = |_T_8 ? _GEN_2360 : _GEN_2424; // @[utils.scala 62:60]
  wire [4:0] _GEN_2489 = |_T_8 ? _GEN_2361 : _GEN_2425; // @[utils.scala 62:60]
  wire [4:0] _GEN_2490 = |_T_8 ? _GEN_2362 : _GEN_2426; // @[utils.scala 62:60]
  wire [4:0] _GEN_2491 = |_T_8 ? _GEN_2363 : _GEN_2427; // @[utils.scala 62:60]
  wire [4:0] _GEN_2492 = |_T_8 ? _GEN_2364 : _GEN_2428; // @[utils.scala 62:60]
  wire [4:0] _GEN_2493 = |_T_8 ? _GEN_2365 : _GEN_2429; // @[utils.scala 62:60]
  wire [4:0] _GEN_2494 = |_T_8 ? _GEN_2366 : _GEN_2430; // @[utils.scala 62:60]
  wire [4:0] _GEN_2495 = |_T_8 ? _GEN_2367 : _GEN_2431; // @[utils.scala 62:60]
  wire [4:0] _GEN_2496 = |_T_8 ? _GEN_2368 : _GEN_2432; // @[utils.scala 62:60]
  wire [4:0] _GEN_2497 = |_T_8 ? _GEN_2369 : _GEN_2433; // @[utils.scala 62:60]
  wire [4:0] _GEN_2498 = |_T_8 ? _GEN_2370 : _GEN_2434; // @[utils.scala 62:60]
  wire [4:0] _GEN_2499 = |_T_8 ? _GEN_2371 : _GEN_2435; // @[utils.scala 62:60]
  wire [4:0] _GEN_2500 = |_T_8 ? _GEN_2372 : _GEN_2436; // @[utils.scala 62:60]
  wire [4:0] _GEN_2501 = |_T_8 ? _GEN_2373 : _GEN_2437; // @[utils.scala 62:60]
  wire [4:0] _GEN_2502 = |_T_8 ? _GEN_2374 : _GEN_2438; // @[utils.scala 62:60]
  wire [4:0] _GEN_2503 = |_T_8 ? _GEN_2375 : _GEN_2439; // @[utils.scala 62:60]
  wire [4:0] _GEN_2504 = |_T_8 ? _GEN_2376 : _GEN_2440; // @[utils.scala 62:60]
  wire [4:0] _GEN_2505 = |_T_8 ? _GEN_2377 : _GEN_2441; // @[utils.scala 62:60]
  wire [4:0] _GEN_2506 = |_T_8 ? _GEN_2378 : _GEN_2442; // @[utils.scala 62:60]
  wire [4:0] _GEN_2507 = |_T_8 ? _GEN_2379 : _GEN_2443; // @[utils.scala 62:60]
  wire [4:0] _GEN_2508 = |_T_8 ? _GEN_2380 : _GEN_2444; // @[utils.scala 62:60]
  wire [4:0] _GEN_2509 = |_T_8 ? _GEN_2381 : _GEN_2445; // @[utils.scala 62:60]
  wire [4:0] _GEN_2510 = |_T_8 ? _GEN_2382 : _GEN_2446; // @[utils.scala 62:60]
  wire [4:0] _GEN_2511 = |_T_8 ? _GEN_2383 : _GEN_2447; // @[utils.scala 62:60]
  wire [4:0] _GEN_2512 = |_T_8 ? _GEN_2384 : _GEN_2448; // @[utils.scala 62:60]
  wire [4:0] _GEN_2513 = |_T_8 ? _GEN_2385 : _GEN_2449; // @[utils.scala 62:60]
  wire [4:0] _GEN_2514 = |_T_8 ? _GEN_2386 : _GEN_2450; // @[utils.scala 62:60]
  wire [4:0] _GEN_2515 = |_T_8 ? _GEN_2387 : _GEN_2451; // @[utils.scala 62:60]
  wire [4:0] _GEN_2516 = |_T_8 ? _GEN_2388 : _GEN_2452; // @[utils.scala 62:60]
  wire [4:0] _GEN_2517 = |_T_8 ? _GEN_2389 : _GEN_2453; // @[utils.scala 62:60]
  wire [4:0] _GEN_2518 = |_T_8 ? _GEN_2390 : _GEN_2454; // @[utils.scala 62:60]
  wire [4:0] _GEN_2519 = |_T_8 ? _GEN_2391 : _GEN_2455; // @[utils.scala 62:60]
  wire [4:0] _GEN_2520 = |_T_8 ? _GEN_2392 : _GEN_2456; // @[utils.scala 62:60]
  wire [4:0] _GEN_2521 = |_T_8 ? _GEN_2393 : _GEN_2457; // @[utils.scala 62:60]
  wire [4:0] _GEN_2522 = |_T_8 ? _GEN_2394 : _GEN_2458; // @[utils.scala 62:60]
  wire [4:0] _GEN_2523 = |_T_8 ? _GEN_2395 : _GEN_2459; // @[utils.scala 62:60]
  wire [4:0] _GEN_2524 = |_T_8 ? _GEN_2396 : _GEN_2460; // @[utils.scala 62:60]
  wire [4:0] _GEN_2525 = |_T_8 ? _GEN_2397 : _GEN_2461; // @[utils.scala 62:60]
  wire  _GEN_2526 = 6'h0 == writePtr ? write_data_branch_valid : _GEN_1118; // @[utils.scala 67:{22,22}]
  wire  _GEN_2527 = 6'h1 == writePtr ? write_data_branch_valid : _GEN_1119; // @[utils.scala 67:{22,22}]
  wire  _GEN_2528 = 6'h2 == writePtr ? write_data_branch_valid : _GEN_1120; // @[utils.scala 67:{22,22}]
  wire  _GEN_2529 = 6'h3 == writePtr ? write_data_branch_valid : _GEN_1121; // @[utils.scala 67:{22,22}]
  wire  _GEN_2530 = 6'h4 == writePtr ? write_data_branch_valid : _GEN_1122; // @[utils.scala 67:{22,22}]
  wire  _GEN_2531 = 6'h5 == writePtr ? write_data_branch_valid : _GEN_1123; // @[utils.scala 67:{22,22}]
  wire  _GEN_2532 = 6'h6 == writePtr ? write_data_branch_valid : _GEN_1124; // @[utils.scala 67:{22,22}]
  wire  _GEN_2533 = 6'h7 == writePtr ? write_data_branch_valid : _GEN_1125; // @[utils.scala 67:{22,22}]
  wire  _GEN_2534 = 6'h8 == writePtr ? write_data_branch_valid : _GEN_1126; // @[utils.scala 67:{22,22}]
  wire  _GEN_2535 = 6'h9 == writePtr ? write_data_branch_valid : _GEN_1127; // @[utils.scala 67:{22,22}]
  wire  _GEN_2536 = 6'ha == writePtr ? write_data_branch_valid : _GEN_1128; // @[utils.scala 67:{22,22}]
  wire  _GEN_2537 = 6'hb == writePtr ? write_data_branch_valid : _GEN_1129; // @[utils.scala 67:{22,22}]
  wire  _GEN_2538 = 6'hc == writePtr ? write_data_branch_valid : _GEN_1130; // @[utils.scala 67:{22,22}]
  wire  _GEN_2539 = 6'hd == writePtr ? write_data_branch_valid : _GEN_1131; // @[utils.scala 67:{22,22}]
  wire  _GEN_2540 = 6'he == writePtr ? write_data_branch_valid : _GEN_1132; // @[utils.scala 67:{22,22}]
  wire  _GEN_2541 = 6'hf == writePtr ? write_data_branch_valid : _GEN_1133; // @[utils.scala 67:{22,22}]
  wire  _GEN_2542 = 6'h10 == writePtr ? write_data_branch_valid : _GEN_1134; // @[utils.scala 67:{22,22}]
  wire  _GEN_2543 = 6'h11 == writePtr ? write_data_branch_valid : _GEN_1135; // @[utils.scala 67:{22,22}]
  wire  _GEN_2544 = 6'h12 == writePtr ? write_data_branch_valid : _GEN_1136; // @[utils.scala 67:{22,22}]
  wire  _GEN_2545 = 6'h13 == writePtr ? write_data_branch_valid : _GEN_1137; // @[utils.scala 67:{22,22}]
  wire  _GEN_2546 = 6'h14 == writePtr ? write_data_branch_valid : _GEN_1138; // @[utils.scala 67:{22,22}]
  wire  _GEN_2547 = 6'h15 == writePtr ? write_data_branch_valid : _GEN_1139; // @[utils.scala 67:{22,22}]
  wire  _GEN_2548 = 6'h16 == writePtr ? write_data_branch_valid : _GEN_1140; // @[utils.scala 67:{22,22}]
  wire  _GEN_2549 = 6'h17 == writePtr ? write_data_branch_valid : _GEN_1141; // @[utils.scala 67:{22,22}]
  wire  _GEN_2550 = 6'h18 == writePtr ? write_data_branch_valid : _GEN_1142; // @[utils.scala 67:{22,22}]
  wire  _GEN_2551 = 6'h19 == writePtr ? write_data_branch_valid : _GEN_1143; // @[utils.scala 67:{22,22}]
  wire  _GEN_2552 = 6'h1a == writePtr ? write_data_branch_valid : _GEN_1144; // @[utils.scala 67:{22,22}]
  wire  _GEN_2553 = 6'h1b == writePtr ? write_data_branch_valid : _GEN_1145; // @[utils.scala 67:{22,22}]
  wire  _GEN_2554 = 6'h1c == writePtr ? write_data_branch_valid : _GEN_1146; // @[utils.scala 67:{22,22}]
  wire  _GEN_2555 = 6'h1d == writePtr ? write_data_branch_valid : _GEN_1147; // @[utils.scala 67:{22,22}]
  wire  _GEN_2556 = 6'h1e == writePtr ? write_data_branch_valid : _GEN_1148; // @[utils.scala 67:{22,22}]
  wire  _GEN_2557 = 6'h1f == writePtr ? write_data_branch_valid : _GEN_1149; // @[utils.scala 67:{22,22}]
  wire  _GEN_2558 = 6'h20 == writePtr ? write_data_branch_valid : _GEN_1150; // @[utils.scala 67:{22,22}]
  wire  _GEN_2559 = 6'h21 == writePtr ? write_data_branch_valid : _GEN_1151; // @[utils.scala 67:{22,22}]
  wire  _GEN_2560 = 6'h22 == writePtr ? write_data_branch_valid : _GEN_1152; // @[utils.scala 67:{22,22}]
  wire  _GEN_2561 = 6'h23 == writePtr ? write_data_branch_valid : _GEN_1153; // @[utils.scala 67:{22,22}]
  wire  _GEN_2562 = 6'h24 == writePtr ? write_data_branch_valid : _GEN_1154; // @[utils.scala 67:{22,22}]
  wire  _GEN_2563 = 6'h25 == writePtr ? write_data_branch_valid : _GEN_1155; // @[utils.scala 67:{22,22}]
  wire  _GEN_2564 = 6'h26 == writePtr ? write_data_branch_valid : _GEN_1156; // @[utils.scala 67:{22,22}]
  wire  _GEN_2565 = 6'h27 == writePtr ? write_data_branch_valid : _GEN_1157; // @[utils.scala 67:{22,22}]
  wire  _GEN_2566 = 6'h28 == writePtr ? write_data_branch_valid : _GEN_1158; // @[utils.scala 67:{22,22}]
  wire  _GEN_2567 = 6'h29 == writePtr ? write_data_branch_valid : _GEN_1159; // @[utils.scala 67:{22,22}]
  wire  _GEN_2568 = 6'h2a == writePtr ? write_data_branch_valid : _GEN_1160; // @[utils.scala 67:{22,22}]
  wire  _GEN_2569 = 6'h2b == writePtr ? write_data_branch_valid : _GEN_1161; // @[utils.scala 67:{22,22}]
  wire  _GEN_2570 = 6'h2c == writePtr ? write_data_branch_valid : _GEN_1162; // @[utils.scala 67:{22,22}]
  wire  _GEN_2571 = 6'h2d == writePtr ? write_data_branch_valid : _GEN_1163; // @[utils.scala 67:{22,22}]
  wire  _GEN_2572 = 6'h2e == writePtr ? write_data_branch_valid : _GEN_1164; // @[utils.scala 67:{22,22}]
  wire  _GEN_2573 = 6'h2f == writePtr ? write_data_branch_valid : _GEN_1165; // @[utils.scala 67:{22,22}]
  wire  _GEN_2574 = 6'h30 == writePtr ? write_data_branch_valid : _GEN_1166; // @[utils.scala 67:{22,22}]
  wire  _GEN_2575 = 6'h31 == writePtr ? write_data_branch_valid : _GEN_1167; // @[utils.scala 67:{22,22}]
  wire  _GEN_2576 = 6'h32 == writePtr ? write_data_branch_valid : _GEN_1168; // @[utils.scala 67:{22,22}]
  wire  _GEN_2577 = 6'h33 == writePtr ? write_data_branch_valid : _GEN_1169; // @[utils.scala 67:{22,22}]
  wire  _GEN_2578 = 6'h34 == writePtr ? write_data_branch_valid : _GEN_1170; // @[utils.scala 67:{22,22}]
  wire  _GEN_2579 = 6'h35 == writePtr ? write_data_branch_valid : _GEN_1171; // @[utils.scala 67:{22,22}]
  wire  _GEN_2580 = 6'h36 == writePtr ? write_data_branch_valid : _GEN_1172; // @[utils.scala 67:{22,22}]
  wire  _GEN_2581 = 6'h37 == writePtr ? write_data_branch_valid : _GEN_1173; // @[utils.scala 67:{22,22}]
  wire  _GEN_2582 = 6'h38 == writePtr ? write_data_branch_valid : _GEN_1174; // @[utils.scala 67:{22,22}]
  wire  _GEN_2583 = 6'h39 == writePtr ? write_data_branch_valid : _GEN_1175; // @[utils.scala 67:{22,22}]
  wire  _GEN_2584 = 6'h3a == writePtr ? write_data_branch_valid : _GEN_1176; // @[utils.scala 67:{22,22}]
  wire  _GEN_2585 = 6'h3b == writePtr ? write_data_branch_valid : _GEN_1177; // @[utils.scala 67:{22,22}]
  wire  _GEN_2586 = 6'h3c == writePtr ? write_data_branch_valid : _GEN_1178; // @[utils.scala 67:{22,22}]
  wire  _GEN_2587 = 6'h3d == writePtr ? write_data_branch_valid : _GEN_1179; // @[utils.scala 67:{22,22}]
  wire  _GEN_2588 = 6'h3e == writePtr ? write_data_branch_valid : _GEN_1180; // @[utils.scala 67:{22,22}]
  wire  _GEN_2589 = 6'h3f == writePtr ? write_data_branch_valid : _GEN_1181; // @[utils.scala 67:{22,22}]
  wire  _GEN_2590 = 6'h0 == writePtr ? 1'h0 : _GEN_1118; // @[utils.scala 71:{24,24}]
  wire  _GEN_2591 = 6'h1 == writePtr ? 1'h0 : _GEN_1119; // @[utils.scala 71:{24,24}]
  wire  _GEN_2592 = 6'h2 == writePtr ? 1'h0 : _GEN_1120; // @[utils.scala 71:{24,24}]
  wire  _GEN_2593 = 6'h3 == writePtr ? 1'h0 : _GEN_1121; // @[utils.scala 71:{24,24}]
  wire  _GEN_2594 = 6'h4 == writePtr ? 1'h0 : _GEN_1122; // @[utils.scala 71:{24,24}]
  wire  _GEN_2595 = 6'h5 == writePtr ? 1'h0 : _GEN_1123; // @[utils.scala 71:{24,24}]
  wire  _GEN_2596 = 6'h6 == writePtr ? 1'h0 : _GEN_1124; // @[utils.scala 71:{24,24}]
  wire  _GEN_2597 = 6'h7 == writePtr ? 1'h0 : _GEN_1125; // @[utils.scala 71:{24,24}]
  wire  _GEN_2598 = 6'h8 == writePtr ? 1'h0 : _GEN_1126; // @[utils.scala 71:{24,24}]
  wire  _GEN_2599 = 6'h9 == writePtr ? 1'h0 : _GEN_1127; // @[utils.scala 71:{24,24}]
  wire  _GEN_2600 = 6'ha == writePtr ? 1'h0 : _GEN_1128; // @[utils.scala 71:{24,24}]
  wire  _GEN_2601 = 6'hb == writePtr ? 1'h0 : _GEN_1129; // @[utils.scala 71:{24,24}]
  wire  _GEN_2602 = 6'hc == writePtr ? 1'h0 : _GEN_1130; // @[utils.scala 71:{24,24}]
  wire  _GEN_2603 = 6'hd == writePtr ? 1'h0 : _GEN_1131; // @[utils.scala 71:{24,24}]
  wire  _GEN_2604 = 6'he == writePtr ? 1'h0 : _GEN_1132; // @[utils.scala 71:{24,24}]
  wire  _GEN_2605 = 6'hf == writePtr ? 1'h0 : _GEN_1133; // @[utils.scala 71:{24,24}]
  wire  _GEN_2606 = 6'h10 == writePtr ? 1'h0 : _GEN_1134; // @[utils.scala 71:{24,24}]
  wire  _GEN_2607 = 6'h11 == writePtr ? 1'h0 : _GEN_1135; // @[utils.scala 71:{24,24}]
  wire  _GEN_2608 = 6'h12 == writePtr ? 1'h0 : _GEN_1136; // @[utils.scala 71:{24,24}]
  wire  _GEN_2609 = 6'h13 == writePtr ? 1'h0 : _GEN_1137; // @[utils.scala 71:{24,24}]
  wire  _GEN_2610 = 6'h14 == writePtr ? 1'h0 : _GEN_1138; // @[utils.scala 71:{24,24}]
  wire  _GEN_2611 = 6'h15 == writePtr ? 1'h0 : _GEN_1139; // @[utils.scala 71:{24,24}]
  wire  _GEN_2612 = 6'h16 == writePtr ? 1'h0 : _GEN_1140; // @[utils.scala 71:{24,24}]
  wire  _GEN_2613 = 6'h17 == writePtr ? 1'h0 : _GEN_1141; // @[utils.scala 71:{24,24}]
  wire  _GEN_2614 = 6'h18 == writePtr ? 1'h0 : _GEN_1142; // @[utils.scala 71:{24,24}]
  wire  _GEN_2615 = 6'h19 == writePtr ? 1'h0 : _GEN_1143; // @[utils.scala 71:{24,24}]
  wire  _GEN_2616 = 6'h1a == writePtr ? 1'h0 : _GEN_1144; // @[utils.scala 71:{24,24}]
  wire  _GEN_2617 = 6'h1b == writePtr ? 1'h0 : _GEN_1145; // @[utils.scala 71:{24,24}]
  wire  _GEN_2618 = 6'h1c == writePtr ? 1'h0 : _GEN_1146; // @[utils.scala 71:{24,24}]
  wire  _GEN_2619 = 6'h1d == writePtr ? 1'h0 : _GEN_1147; // @[utils.scala 71:{24,24}]
  wire  _GEN_2620 = 6'h1e == writePtr ? 1'h0 : _GEN_1148; // @[utils.scala 71:{24,24}]
  wire  _GEN_2621 = 6'h1f == writePtr ? 1'h0 : _GEN_1149; // @[utils.scala 71:{24,24}]
  wire  _GEN_2622 = 6'h20 == writePtr ? 1'h0 : _GEN_1150; // @[utils.scala 71:{24,24}]
  wire  _GEN_2623 = 6'h21 == writePtr ? 1'h0 : _GEN_1151; // @[utils.scala 71:{24,24}]
  wire  _GEN_2624 = 6'h22 == writePtr ? 1'h0 : _GEN_1152; // @[utils.scala 71:{24,24}]
  wire  _GEN_2625 = 6'h23 == writePtr ? 1'h0 : _GEN_1153; // @[utils.scala 71:{24,24}]
  wire  _GEN_2626 = 6'h24 == writePtr ? 1'h0 : _GEN_1154; // @[utils.scala 71:{24,24}]
  wire  _GEN_2627 = 6'h25 == writePtr ? 1'h0 : _GEN_1155; // @[utils.scala 71:{24,24}]
  wire  _GEN_2628 = 6'h26 == writePtr ? 1'h0 : _GEN_1156; // @[utils.scala 71:{24,24}]
  wire  _GEN_2629 = 6'h27 == writePtr ? 1'h0 : _GEN_1157; // @[utils.scala 71:{24,24}]
  wire  _GEN_2630 = 6'h28 == writePtr ? 1'h0 : _GEN_1158; // @[utils.scala 71:{24,24}]
  wire  _GEN_2631 = 6'h29 == writePtr ? 1'h0 : _GEN_1159; // @[utils.scala 71:{24,24}]
  wire  _GEN_2632 = 6'h2a == writePtr ? 1'h0 : _GEN_1160; // @[utils.scala 71:{24,24}]
  wire  _GEN_2633 = 6'h2b == writePtr ? 1'h0 : _GEN_1161; // @[utils.scala 71:{24,24}]
  wire  _GEN_2634 = 6'h2c == writePtr ? 1'h0 : _GEN_1162; // @[utils.scala 71:{24,24}]
  wire  _GEN_2635 = 6'h2d == writePtr ? 1'h0 : _GEN_1163; // @[utils.scala 71:{24,24}]
  wire  _GEN_2636 = 6'h2e == writePtr ? 1'h0 : _GEN_1164; // @[utils.scala 71:{24,24}]
  wire  _GEN_2637 = 6'h2f == writePtr ? 1'h0 : _GEN_1165; // @[utils.scala 71:{24,24}]
  wire  _GEN_2638 = 6'h30 == writePtr ? 1'h0 : _GEN_1166; // @[utils.scala 71:{24,24}]
  wire  _GEN_2639 = 6'h31 == writePtr ? 1'h0 : _GEN_1167; // @[utils.scala 71:{24,24}]
  wire  _GEN_2640 = 6'h32 == writePtr ? 1'h0 : _GEN_1168; // @[utils.scala 71:{24,24}]
  wire  _GEN_2641 = 6'h33 == writePtr ? 1'h0 : _GEN_1169; // @[utils.scala 71:{24,24}]
  wire  _GEN_2642 = 6'h34 == writePtr ? 1'h0 : _GEN_1170; // @[utils.scala 71:{24,24}]
  wire  _GEN_2643 = 6'h35 == writePtr ? 1'h0 : _GEN_1171; // @[utils.scala 71:{24,24}]
  wire  _GEN_2644 = 6'h36 == writePtr ? 1'h0 : _GEN_1172; // @[utils.scala 71:{24,24}]
  wire  _GEN_2645 = 6'h37 == writePtr ? 1'h0 : _GEN_1173; // @[utils.scala 71:{24,24}]
  wire  _GEN_2646 = 6'h38 == writePtr ? 1'h0 : _GEN_1174; // @[utils.scala 71:{24,24}]
  wire  _GEN_2647 = 6'h39 == writePtr ? 1'h0 : _GEN_1175; // @[utils.scala 71:{24,24}]
  wire  _GEN_2648 = 6'h3a == writePtr ? 1'h0 : _GEN_1176; // @[utils.scala 71:{24,24}]
  wire  _GEN_2649 = 6'h3b == writePtr ? 1'h0 : _GEN_1177; // @[utils.scala 71:{24,24}]
  wire  _GEN_2650 = 6'h3c == writePtr ? 1'h0 : _GEN_1178; // @[utils.scala 71:{24,24}]
  wire  _GEN_2651 = 6'h3d == writePtr ? 1'h0 : _GEN_1179; // @[utils.scala 71:{24,24}]
  wire  _GEN_2652 = 6'h3e == writePtr ? 1'h0 : _GEN_1180; // @[utils.scala 71:{24,24}]
  wire  _GEN_2653 = 6'h3f == writePtr ? 1'h0 : _GEN_1181; // @[utils.scala 71:{24,24}]
  wire [4:0] _GEN_2654 = 6'h0 == writePtr ? 5'h0 : _GEN_1182; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2655 = 6'h1 == writePtr ? 5'h0 : _GEN_1183; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2656 = 6'h2 == writePtr ? 5'h0 : _GEN_1184; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2657 = 6'h3 == writePtr ? 5'h0 : _GEN_1185; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2658 = 6'h4 == writePtr ? 5'h0 : _GEN_1186; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2659 = 6'h5 == writePtr ? 5'h0 : _GEN_1187; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2660 = 6'h6 == writePtr ? 5'h0 : _GEN_1188; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2661 = 6'h7 == writePtr ? 5'h0 : _GEN_1189; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2662 = 6'h8 == writePtr ? 5'h0 : _GEN_1190; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2663 = 6'h9 == writePtr ? 5'h0 : _GEN_1191; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2664 = 6'ha == writePtr ? 5'h0 : _GEN_1192; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2665 = 6'hb == writePtr ? 5'h0 : _GEN_1193; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2666 = 6'hc == writePtr ? 5'h0 : _GEN_1194; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2667 = 6'hd == writePtr ? 5'h0 : _GEN_1195; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2668 = 6'he == writePtr ? 5'h0 : _GEN_1196; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2669 = 6'hf == writePtr ? 5'h0 : _GEN_1197; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2670 = 6'h10 == writePtr ? 5'h0 : _GEN_1198; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2671 = 6'h11 == writePtr ? 5'h0 : _GEN_1199; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2672 = 6'h12 == writePtr ? 5'h0 : _GEN_1200; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2673 = 6'h13 == writePtr ? 5'h0 : _GEN_1201; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2674 = 6'h14 == writePtr ? 5'h0 : _GEN_1202; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2675 = 6'h15 == writePtr ? 5'h0 : _GEN_1203; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2676 = 6'h16 == writePtr ? 5'h0 : _GEN_1204; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2677 = 6'h17 == writePtr ? 5'h0 : _GEN_1205; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2678 = 6'h18 == writePtr ? 5'h0 : _GEN_1206; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2679 = 6'h19 == writePtr ? 5'h0 : _GEN_1207; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2680 = 6'h1a == writePtr ? 5'h0 : _GEN_1208; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2681 = 6'h1b == writePtr ? 5'h0 : _GEN_1209; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2682 = 6'h1c == writePtr ? 5'h0 : _GEN_1210; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2683 = 6'h1d == writePtr ? 5'h0 : _GEN_1211; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2684 = 6'h1e == writePtr ? 5'h0 : _GEN_1212; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2685 = 6'h1f == writePtr ? 5'h0 : _GEN_1213; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2686 = 6'h20 == writePtr ? 5'h0 : _GEN_1214; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2687 = 6'h21 == writePtr ? 5'h0 : _GEN_1215; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2688 = 6'h22 == writePtr ? 5'h0 : _GEN_1216; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2689 = 6'h23 == writePtr ? 5'h0 : _GEN_1217; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2690 = 6'h24 == writePtr ? 5'h0 : _GEN_1218; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2691 = 6'h25 == writePtr ? 5'h0 : _GEN_1219; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2692 = 6'h26 == writePtr ? 5'h0 : _GEN_1220; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2693 = 6'h27 == writePtr ? 5'h0 : _GEN_1221; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2694 = 6'h28 == writePtr ? 5'h0 : _GEN_1222; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2695 = 6'h29 == writePtr ? 5'h0 : _GEN_1223; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2696 = 6'h2a == writePtr ? 5'h0 : _GEN_1224; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2697 = 6'h2b == writePtr ? 5'h0 : _GEN_1225; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2698 = 6'h2c == writePtr ? 5'h0 : _GEN_1226; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2699 = 6'h2d == writePtr ? 5'h0 : _GEN_1227; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2700 = 6'h2e == writePtr ? 5'h0 : _GEN_1228; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2701 = 6'h2f == writePtr ? 5'h0 : _GEN_1229; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2702 = 6'h30 == writePtr ? 5'h0 : _GEN_1230; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2703 = 6'h31 == writePtr ? 5'h0 : _GEN_1231; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2704 = 6'h32 == writePtr ? 5'h0 : _GEN_1232; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2705 = 6'h33 == writePtr ? 5'h0 : _GEN_1233; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2706 = 6'h34 == writePtr ? 5'h0 : _GEN_1234; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2707 = 6'h35 == writePtr ? 5'h0 : _GEN_1235; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2708 = 6'h36 == writePtr ? 5'h0 : _GEN_1236; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2709 = 6'h37 == writePtr ? 5'h0 : _GEN_1237; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2710 = 6'h38 == writePtr ? 5'h0 : _GEN_1238; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2711 = 6'h39 == writePtr ? 5'h0 : _GEN_1239; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2712 = 6'h3a == writePtr ? 5'h0 : _GEN_1240; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2713 = 6'h3b == writePtr ? 5'h0 : _GEN_1241; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2714 = 6'h3c == writePtr ? 5'h0 : _GEN_1242; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2715 = 6'h3d == writePtr ? 5'h0 : _GEN_1243; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2716 = 6'h3e == writePtr ? 5'h0 : _GEN_1244; // @[utils.scala 72:{23,23}]
  wire [4:0] _GEN_2717 = 6'h3f == writePtr ? 5'h0 : _GEN_1245; // @[utils.scala 72:{23,23}]
  wire  _GEN_2846 = _T_9 ? _GEN_2590 : _GEN_2526; // @[utils.scala 70:60]
  wire  _GEN_2847 = _T_9 ? _GEN_2591 : _GEN_2527; // @[utils.scala 70:60]
  wire  _GEN_2848 = _T_9 ? _GEN_2592 : _GEN_2528; // @[utils.scala 70:60]
  wire  _GEN_2849 = _T_9 ? _GEN_2593 : _GEN_2529; // @[utils.scala 70:60]
  wire  _GEN_2850 = _T_9 ? _GEN_2594 : _GEN_2530; // @[utils.scala 70:60]
  wire  _GEN_2851 = _T_9 ? _GEN_2595 : _GEN_2531; // @[utils.scala 70:60]
  wire  _GEN_2852 = _T_9 ? _GEN_2596 : _GEN_2532; // @[utils.scala 70:60]
  wire  _GEN_2853 = _T_9 ? _GEN_2597 : _GEN_2533; // @[utils.scala 70:60]
  wire  _GEN_2854 = _T_9 ? _GEN_2598 : _GEN_2534; // @[utils.scala 70:60]
  wire  _GEN_2855 = _T_9 ? _GEN_2599 : _GEN_2535; // @[utils.scala 70:60]
  wire  _GEN_2856 = _T_9 ? _GEN_2600 : _GEN_2536; // @[utils.scala 70:60]
  wire  _GEN_2857 = _T_9 ? _GEN_2601 : _GEN_2537; // @[utils.scala 70:60]
  wire  _GEN_2858 = _T_9 ? _GEN_2602 : _GEN_2538; // @[utils.scala 70:60]
  wire  _GEN_2859 = _T_9 ? _GEN_2603 : _GEN_2539; // @[utils.scala 70:60]
  wire  _GEN_2860 = _T_9 ? _GEN_2604 : _GEN_2540; // @[utils.scala 70:60]
  wire  _GEN_2861 = _T_9 ? _GEN_2605 : _GEN_2541; // @[utils.scala 70:60]
  wire  _GEN_2862 = _T_9 ? _GEN_2606 : _GEN_2542; // @[utils.scala 70:60]
  wire  _GEN_2863 = _T_9 ? _GEN_2607 : _GEN_2543; // @[utils.scala 70:60]
  wire  _GEN_2864 = _T_9 ? _GEN_2608 : _GEN_2544; // @[utils.scala 70:60]
  wire  _GEN_2865 = _T_9 ? _GEN_2609 : _GEN_2545; // @[utils.scala 70:60]
  wire  _GEN_2866 = _T_9 ? _GEN_2610 : _GEN_2546; // @[utils.scala 70:60]
  wire  _GEN_2867 = _T_9 ? _GEN_2611 : _GEN_2547; // @[utils.scala 70:60]
  wire  _GEN_2868 = _T_9 ? _GEN_2612 : _GEN_2548; // @[utils.scala 70:60]
  wire  _GEN_2869 = _T_9 ? _GEN_2613 : _GEN_2549; // @[utils.scala 70:60]
  wire  _GEN_2870 = _T_9 ? _GEN_2614 : _GEN_2550; // @[utils.scala 70:60]
  wire  _GEN_2871 = _T_9 ? _GEN_2615 : _GEN_2551; // @[utils.scala 70:60]
  wire  _GEN_2872 = _T_9 ? _GEN_2616 : _GEN_2552; // @[utils.scala 70:60]
  wire  _GEN_2873 = _T_9 ? _GEN_2617 : _GEN_2553; // @[utils.scala 70:60]
  wire  _GEN_2874 = _T_9 ? _GEN_2618 : _GEN_2554; // @[utils.scala 70:60]
  wire  _GEN_2875 = _T_9 ? _GEN_2619 : _GEN_2555; // @[utils.scala 70:60]
  wire  _GEN_2876 = _T_9 ? _GEN_2620 : _GEN_2556; // @[utils.scala 70:60]
  wire  _GEN_2877 = _T_9 ? _GEN_2621 : _GEN_2557; // @[utils.scala 70:60]
  wire  _GEN_2878 = _T_9 ? _GEN_2622 : _GEN_2558; // @[utils.scala 70:60]
  wire  _GEN_2879 = _T_9 ? _GEN_2623 : _GEN_2559; // @[utils.scala 70:60]
  wire  _GEN_2880 = _T_9 ? _GEN_2624 : _GEN_2560; // @[utils.scala 70:60]
  wire  _GEN_2881 = _T_9 ? _GEN_2625 : _GEN_2561; // @[utils.scala 70:60]
  wire  _GEN_2882 = _T_9 ? _GEN_2626 : _GEN_2562; // @[utils.scala 70:60]
  wire  _GEN_2883 = _T_9 ? _GEN_2627 : _GEN_2563; // @[utils.scala 70:60]
  wire  _GEN_2884 = _T_9 ? _GEN_2628 : _GEN_2564; // @[utils.scala 70:60]
  wire  _GEN_2885 = _T_9 ? _GEN_2629 : _GEN_2565; // @[utils.scala 70:60]
  wire  _GEN_2886 = _T_9 ? _GEN_2630 : _GEN_2566; // @[utils.scala 70:60]
  wire  _GEN_2887 = _T_9 ? _GEN_2631 : _GEN_2567; // @[utils.scala 70:60]
  wire  _GEN_2888 = _T_9 ? _GEN_2632 : _GEN_2568; // @[utils.scala 70:60]
  wire  _GEN_2889 = _T_9 ? _GEN_2633 : _GEN_2569; // @[utils.scala 70:60]
  wire  _GEN_2890 = _T_9 ? _GEN_2634 : _GEN_2570; // @[utils.scala 70:60]
  wire  _GEN_2891 = _T_9 ? _GEN_2635 : _GEN_2571; // @[utils.scala 70:60]
  wire  _GEN_2892 = _T_9 ? _GEN_2636 : _GEN_2572; // @[utils.scala 70:60]
  wire  _GEN_2893 = _T_9 ? _GEN_2637 : _GEN_2573; // @[utils.scala 70:60]
  wire  _GEN_2894 = _T_9 ? _GEN_2638 : _GEN_2574; // @[utils.scala 70:60]
  wire  _GEN_2895 = _T_9 ? _GEN_2639 : _GEN_2575; // @[utils.scala 70:60]
  wire  _GEN_2896 = _T_9 ? _GEN_2640 : _GEN_2576; // @[utils.scala 70:60]
  wire  _GEN_2897 = _T_9 ? _GEN_2641 : _GEN_2577; // @[utils.scala 70:60]
  wire  _GEN_2898 = _T_9 ? _GEN_2642 : _GEN_2578; // @[utils.scala 70:60]
  wire  _GEN_2899 = _T_9 ? _GEN_2643 : _GEN_2579; // @[utils.scala 70:60]
  wire  _GEN_2900 = _T_9 ? _GEN_2644 : _GEN_2580; // @[utils.scala 70:60]
  wire  _GEN_2901 = _T_9 ? _GEN_2645 : _GEN_2581; // @[utils.scala 70:60]
  wire  _GEN_2902 = _T_9 ? _GEN_2646 : _GEN_2582; // @[utils.scala 70:60]
  wire  _GEN_2903 = _T_9 ? _GEN_2647 : _GEN_2583; // @[utils.scala 70:60]
  wire  _GEN_2904 = _T_9 ? _GEN_2648 : _GEN_2584; // @[utils.scala 70:60]
  wire  _GEN_2905 = _T_9 ? _GEN_2649 : _GEN_2585; // @[utils.scala 70:60]
  wire  _GEN_2906 = _T_9 ? _GEN_2650 : _GEN_2586; // @[utils.scala 70:60]
  wire  _GEN_2907 = _T_9 ? _GEN_2651 : _GEN_2587; // @[utils.scala 70:60]
  wire  _GEN_2908 = _T_9 ? _GEN_2652 : _GEN_2588; // @[utils.scala 70:60]
  wire  _GEN_2909 = _T_9 ? _GEN_2653 : _GEN_2589; // @[utils.scala 70:60]
  wire [4:0] _GEN_2910 = _T_9 ? _GEN_2654 : _GEN_2398; // @[utils.scala 70:60]
  wire [4:0] _GEN_2911 = _T_9 ? _GEN_2655 : _GEN_2399; // @[utils.scala 70:60]
  wire [4:0] _GEN_2912 = _T_9 ? _GEN_2656 : _GEN_2400; // @[utils.scala 70:60]
  wire [4:0] _GEN_2913 = _T_9 ? _GEN_2657 : _GEN_2401; // @[utils.scala 70:60]
  wire [4:0] _GEN_2914 = _T_9 ? _GEN_2658 : _GEN_2402; // @[utils.scala 70:60]
  wire [4:0] _GEN_2915 = _T_9 ? _GEN_2659 : _GEN_2403; // @[utils.scala 70:60]
  wire [4:0] _GEN_2916 = _T_9 ? _GEN_2660 : _GEN_2404; // @[utils.scala 70:60]
  wire [4:0] _GEN_2917 = _T_9 ? _GEN_2661 : _GEN_2405; // @[utils.scala 70:60]
  wire [4:0] _GEN_2918 = _T_9 ? _GEN_2662 : _GEN_2406; // @[utils.scala 70:60]
  wire [4:0] _GEN_2919 = _T_9 ? _GEN_2663 : _GEN_2407; // @[utils.scala 70:60]
  wire [4:0] _GEN_2920 = _T_9 ? _GEN_2664 : _GEN_2408; // @[utils.scala 70:60]
  wire [4:0] _GEN_2921 = _T_9 ? _GEN_2665 : _GEN_2409; // @[utils.scala 70:60]
  wire [4:0] _GEN_2922 = _T_9 ? _GEN_2666 : _GEN_2410; // @[utils.scala 70:60]
  wire [4:0] _GEN_2923 = _T_9 ? _GEN_2667 : _GEN_2411; // @[utils.scala 70:60]
  wire [4:0] _GEN_2924 = _T_9 ? _GEN_2668 : _GEN_2412; // @[utils.scala 70:60]
  wire [4:0] _GEN_2925 = _T_9 ? _GEN_2669 : _GEN_2413; // @[utils.scala 70:60]
  wire [4:0] _GEN_2926 = _T_9 ? _GEN_2670 : _GEN_2414; // @[utils.scala 70:60]
  wire [4:0] _GEN_2927 = _T_9 ? _GEN_2671 : _GEN_2415; // @[utils.scala 70:60]
  wire [4:0] _GEN_2928 = _T_9 ? _GEN_2672 : _GEN_2416; // @[utils.scala 70:60]
  wire [4:0] _GEN_2929 = _T_9 ? _GEN_2673 : _GEN_2417; // @[utils.scala 70:60]
  wire [4:0] _GEN_2930 = _T_9 ? _GEN_2674 : _GEN_2418; // @[utils.scala 70:60]
  wire [4:0] _GEN_2931 = _T_9 ? _GEN_2675 : _GEN_2419; // @[utils.scala 70:60]
  wire [4:0] _GEN_2932 = _T_9 ? _GEN_2676 : _GEN_2420; // @[utils.scala 70:60]
  wire [4:0] _GEN_2933 = _T_9 ? _GEN_2677 : _GEN_2421; // @[utils.scala 70:60]
  wire [4:0] _GEN_2934 = _T_9 ? _GEN_2678 : _GEN_2422; // @[utils.scala 70:60]
  wire [4:0] _GEN_2935 = _T_9 ? _GEN_2679 : _GEN_2423; // @[utils.scala 70:60]
  wire [4:0] _GEN_2936 = _T_9 ? _GEN_2680 : _GEN_2424; // @[utils.scala 70:60]
  wire [4:0] _GEN_2937 = _T_9 ? _GEN_2681 : _GEN_2425; // @[utils.scala 70:60]
  wire [4:0] _GEN_2938 = _T_9 ? _GEN_2682 : _GEN_2426; // @[utils.scala 70:60]
  wire [4:0] _GEN_2939 = _T_9 ? _GEN_2683 : _GEN_2427; // @[utils.scala 70:60]
  wire [4:0] _GEN_2940 = _T_9 ? _GEN_2684 : _GEN_2428; // @[utils.scala 70:60]
  wire [4:0] _GEN_2941 = _T_9 ? _GEN_2685 : _GEN_2429; // @[utils.scala 70:60]
  wire [4:0] _GEN_2942 = _T_9 ? _GEN_2686 : _GEN_2430; // @[utils.scala 70:60]
  wire [4:0] _GEN_2943 = _T_9 ? _GEN_2687 : _GEN_2431; // @[utils.scala 70:60]
  wire [4:0] _GEN_2944 = _T_9 ? _GEN_2688 : _GEN_2432; // @[utils.scala 70:60]
  wire [4:0] _GEN_2945 = _T_9 ? _GEN_2689 : _GEN_2433; // @[utils.scala 70:60]
  wire [4:0] _GEN_2946 = _T_9 ? _GEN_2690 : _GEN_2434; // @[utils.scala 70:60]
  wire [4:0] _GEN_2947 = _T_9 ? _GEN_2691 : _GEN_2435; // @[utils.scala 70:60]
  wire [4:0] _GEN_2948 = _T_9 ? _GEN_2692 : _GEN_2436; // @[utils.scala 70:60]
  wire [4:0] _GEN_2949 = _T_9 ? _GEN_2693 : _GEN_2437; // @[utils.scala 70:60]
  wire [4:0] _GEN_2950 = _T_9 ? _GEN_2694 : _GEN_2438; // @[utils.scala 70:60]
  wire [4:0] _GEN_2951 = _T_9 ? _GEN_2695 : _GEN_2439; // @[utils.scala 70:60]
  wire [4:0] _GEN_2952 = _T_9 ? _GEN_2696 : _GEN_2440; // @[utils.scala 70:60]
  wire [4:0] _GEN_2953 = _T_9 ? _GEN_2697 : _GEN_2441; // @[utils.scala 70:60]
  wire [4:0] _GEN_2954 = _T_9 ? _GEN_2698 : _GEN_2442; // @[utils.scala 70:60]
  wire [4:0] _GEN_2955 = _T_9 ? _GEN_2699 : _GEN_2443; // @[utils.scala 70:60]
  wire [4:0] _GEN_2956 = _T_9 ? _GEN_2700 : _GEN_2444; // @[utils.scala 70:60]
  wire [4:0] _GEN_2957 = _T_9 ? _GEN_2701 : _GEN_2445; // @[utils.scala 70:60]
  wire [4:0] _GEN_2958 = _T_9 ? _GEN_2702 : _GEN_2446; // @[utils.scala 70:60]
  wire [4:0] _GEN_2959 = _T_9 ? _GEN_2703 : _GEN_2447; // @[utils.scala 70:60]
  wire [4:0] _GEN_2960 = _T_9 ? _GEN_2704 : _GEN_2448; // @[utils.scala 70:60]
  wire [4:0] _GEN_2961 = _T_9 ? _GEN_2705 : _GEN_2449; // @[utils.scala 70:60]
  wire [4:0] _GEN_2962 = _T_9 ? _GEN_2706 : _GEN_2450; // @[utils.scala 70:60]
  wire [4:0] _GEN_2963 = _T_9 ? _GEN_2707 : _GEN_2451; // @[utils.scala 70:60]
  wire [4:0] _GEN_2964 = _T_9 ? _GEN_2708 : _GEN_2452; // @[utils.scala 70:60]
  wire [4:0] _GEN_2965 = _T_9 ? _GEN_2709 : _GEN_2453; // @[utils.scala 70:60]
  wire [4:0] _GEN_2966 = _T_9 ? _GEN_2710 : _GEN_2454; // @[utils.scala 70:60]
  wire [4:0] _GEN_2967 = _T_9 ? _GEN_2711 : _GEN_2455; // @[utils.scala 70:60]
  wire [4:0] _GEN_2968 = _T_9 ? _GEN_2712 : _GEN_2456; // @[utils.scala 70:60]
  wire [4:0] _GEN_2969 = _T_9 ? _GEN_2713 : _GEN_2457; // @[utils.scala 70:60]
  wire [4:0] _GEN_2970 = _T_9 ? _GEN_2714 : _GEN_2458; // @[utils.scala 70:60]
  wire [4:0] _GEN_2971 = _T_9 ? _GEN_2715 : _GEN_2459; // @[utils.scala 70:60]
  wire [4:0] _GEN_2972 = _T_9 ? _GEN_2716 : _GEN_2460; // @[utils.scala 70:60]
  wire [4:0] _GEN_2973 = _T_9 ? _GEN_2717 : _GEN_2461; // @[utils.scala 70:60]
  wire [4:0] _GEN_2974 = branchOps_passed ? _GEN_2462 : _GEN_2910; // @[utils.scala 60:30]
  wire [4:0] _GEN_2975 = branchOps_passed ? _GEN_2463 : _GEN_2911; // @[utils.scala 60:30]
  wire [4:0] _GEN_2976 = branchOps_passed ? _GEN_2464 : _GEN_2912; // @[utils.scala 60:30]
  wire [4:0] _GEN_2977 = branchOps_passed ? _GEN_2465 : _GEN_2913; // @[utils.scala 60:30]
  wire [4:0] _GEN_2978 = branchOps_passed ? _GEN_2466 : _GEN_2914; // @[utils.scala 60:30]
  wire [4:0] _GEN_2979 = branchOps_passed ? _GEN_2467 : _GEN_2915; // @[utils.scala 60:30]
  wire [4:0] _GEN_2980 = branchOps_passed ? _GEN_2468 : _GEN_2916; // @[utils.scala 60:30]
  wire [4:0] _GEN_2981 = branchOps_passed ? _GEN_2469 : _GEN_2917; // @[utils.scala 60:30]
  wire [4:0] _GEN_2982 = branchOps_passed ? _GEN_2470 : _GEN_2918; // @[utils.scala 60:30]
  wire [4:0] _GEN_2983 = branchOps_passed ? _GEN_2471 : _GEN_2919; // @[utils.scala 60:30]
  wire [4:0] _GEN_2984 = branchOps_passed ? _GEN_2472 : _GEN_2920; // @[utils.scala 60:30]
  wire [4:0] _GEN_2985 = branchOps_passed ? _GEN_2473 : _GEN_2921; // @[utils.scala 60:30]
  wire [4:0] _GEN_2986 = branchOps_passed ? _GEN_2474 : _GEN_2922; // @[utils.scala 60:30]
  wire [4:0] _GEN_2987 = branchOps_passed ? _GEN_2475 : _GEN_2923; // @[utils.scala 60:30]
  wire [4:0] _GEN_2988 = branchOps_passed ? _GEN_2476 : _GEN_2924; // @[utils.scala 60:30]
  wire [4:0] _GEN_2989 = branchOps_passed ? _GEN_2477 : _GEN_2925; // @[utils.scala 60:30]
  wire [4:0] _GEN_2990 = branchOps_passed ? _GEN_2478 : _GEN_2926; // @[utils.scala 60:30]
  wire [4:0] _GEN_2991 = branchOps_passed ? _GEN_2479 : _GEN_2927; // @[utils.scala 60:30]
  wire [4:0] _GEN_2992 = branchOps_passed ? _GEN_2480 : _GEN_2928; // @[utils.scala 60:30]
  wire [4:0] _GEN_2993 = branchOps_passed ? _GEN_2481 : _GEN_2929; // @[utils.scala 60:30]
  wire [4:0] _GEN_2994 = branchOps_passed ? _GEN_2482 : _GEN_2930; // @[utils.scala 60:30]
  wire [4:0] _GEN_2995 = branchOps_passed ? _GEN_2483 : _GEN_2931; // @[utils.scala 60:30]
  wire [4:0] _GEN_2996 = branchOps_passed ? _GEN_2484 : _GEN_2932; // @[utils.scala 60:30]
  wire [4:0] _GEN_2997 = branchOps_passed ? _GEN_2485 : _GEN_2933; // @[utils.scala 60:30]
  wire [4:0] _GEN_2998 = branchOps_passed ? _GEN_2486 : _GEN_2934; // @[utils.scala 60:30]
  wire [4:0] _GEN_2999 = branchOps_passed ? _GEN_2487 : _GEN_2935; // @[utils.scala 60:30]
  wire [4:0] _GEN_3000 = branchOps_passed ? _GEN_2488 : _GEN_2936; // @[utils.scala 60:30]
  wire [4:0] _GEN_3001 = branchOps_passed ? _GEN_2489 : _GEN_2937; // @[utils.scala 60:30]
  wire [4:0] _GEN_3002 = branchOps_passed ? _GEN_2490 : _GEN_2938; // @[utils.scala 60:30]
  wire [4:0] _GEN_3003 = branchOps_passed ? _GEN_2491 : _GEN_2939; // @[utils.scala 60:30]
  wire [4:0] _GEN_3004 = branchOps_passed ? _GEN_2492 : _GEN_2940; // @[utils.scala 60:30]
  wire [4:0] _GEN_3005 = branchOps_passed ? _GEN_2493 : _GEN_2941; // @[utils.scala 60:30]
  wire [4:0] _GEN_3006 = branchOps_passed ? _GEN_2494 : _GEN_2942; // @[utils.scala 60:30]
  wire [4:0] _GEN_3007 = branchOps_passed ? _GEN_2495 : _GEN_2943; // @[utils.scala 60:30]
  wire [4:0] _GEN_3008 = branchOps_passed ? _GEN_2496 : _GEN_2944; // @[utils.scala 60:30]
  wire [4:0] _GEN_3009 = branchOps_passed ? _GEN_2497 : _GEN_2945; // @[utils.scala 60:30]
  wire [4:0] _GEN_3010 = branchOps_passed ? _GEN_2498 : _GEN_2946; // @[utils.scala 60:30]
  wire [4:0] _GEN_3011 = branchOps_passed ? _GEN_2499 : _GEN_2947; // @[utils.scala 60:30]
  wire [4:0] _GEN_3012 = branchOps_passed ? _GEN_2500 : _GEN_2948; // @[utils.scala 60:30]
  wire [4:0] _GEN_3013 = branchOps_passed ? _GEN_2501 : _GEN_2949; // @[utils.scala 60:30]
  wire [4:0] _GEN_3014 = branchOps_passed ? _GEN_2502 : _GEN_2950; // @[utils.scala 60:30]
  wire [4:0] _GEN_3015 = branchOps_passed ? _GEN_2503 : _GEN_2951; // @[utils.scala 60:30]
  wire [4:0] _GEN_3016 = branchOps_passed ? _GEN_2504 : _GEN_2952; // @[utils.scala 60:30]
  wire [4:0] _GEN_3017 = branchOps_passed ? _GEN_2505 : _GEN_2953; // @[utils.scala 60:30]
  wire [4:0] _GEN_3018 = branchOps_passed ? _GEN_2506 : _GEN_2954; // @[utils.scala 60:30]
  wire [4:0] _GEN_3019 = branchOps_passed ? _GEN_2507 : _GEN_2955; // @[utils.scala 60:30]
  wire [4:0] _GEN_3020 = branchOps_passed ? _GEN_2508 : _GEN_2956; // @[utils.scala 60:30]
  wire [4:0] _GEN_3021 = branchOps_passed ? _GEN_2509 : _GEN_2957; // @[utils.scala 60:30]
  wire [4:0] _GEN_3022 = branchOps_passed ? _GEN_2510 : _GEN_2958; // @[utils.scala 60:30]
  wire [4:0] _GEN_3023 = branchOps_passed ? _GEN_2511 : _GEN_2959; // @[utils.scala 60:30]
  wire [4:0] _GEN_3024 = branchOps_passed ? _GEN_2512 : _GEN_2960; // @[utils.scala 60:30]
  wire [4:0] _GEN_3025 = branchOps_passed ? _GEN_2513 : _GEN_2961; // @[utils.scala 60:30]
  wire [4:0] _GEN_3026 = branchOps_passed ? _GEN_2514 : _GEN_2962; // @[utils.scala 60:30]
  wire [4:0] _GEN_3027 = branchOps_passed ? _GEN_2515 : _GEN_2963; // @[utils.scala 60:30]
  wire [4:0] _GEN_3028 = branchOps_passed ? _GEN_2516 : _GEN_2964; // @[utils.scala 60:30]
  wire [4:0] _GEN_3029 = branchOps_passed ? _GEN_2517 : _GEN_2965; // @[utils.scala 60:30]
  wire [4:0] _GEN_3030 = branchOps_passed ? _GEN_2518 : _GEN_2966; // @[utils.scala 60:30]
  wire [4:0] _GEN_3031 = branchOps_passed ? _GEN_2519 : _GEN_2967; // @[utils.scala 60:30]
  wire [4:0] _GEN_3032 = branchOps_passed ? _GEN_2520 : _GEN_2968; // @[utils.scala 60:30]
  wire [4:0] _GEN_3033 = branchOps_passed ? _GEN_2521 : _GEN_2969; // @[utils.scala 60:30]
  wire [4:0] _GEN_3034 = branchOps_passed ? _GEN_2522 : _GEN_2970; // @[utils.scala 60:30]
  wire [4:0] _GEN_3035 = branchOps_passed ? _GEN_2523 : _GEN_2971; // @[utils.scala 60:30]
  wire [4:0] _GEN_3036 = branchOps_passed ? _GEN_2524 : _GEN_2972; // @[utils.scala 60:30]
  wire [4:0] _GEN_3037 = branchOps_passed ? _GEN_2525 : _GEN_2973; // @[utils.scala 60:30]
  wire  _GEN_3038 = branchOps_passed ? _GEN_2526 : _GEN_2846; // @[utils.scala 60:30]
  wire  _GEN_3039 = branchOps_passed ? _GEN_2527 : _GEN_2847; // @[utils.scala 60:30]
  wire  _GEN_3040 = branchOps_passed ? _GEN_2528 : _GEN_2848; // @[utils.scala 60:30]
  wire  _GEN_3041 = branchOps_passed ? _GEN_2529 : _GEN_2849; // @[utils.scala 60:30]
  wire  _GEN_3042 = branchOps_passed ? _GEN_2530 : _GEN_2850; // @[utils.scala 60:30]
  wire  _GEN_3043 = branchOps_passed ? _GEN_2531 : _GEN_2851; // @[utils.scala 60:30]
  wire  _GEN_3044 = branchOps_passed ? _GEN_2532 : _GEN_2852; // @[utils.scala 60:30]
  wire  _GEN_3045 = branchOps_passed ? _GEN_2533 : _GEN_2853; // @[utils.scala 60:30]
  wire  _GEN_3046 = branchOps_passed ? _GEN_2534 : _GEN_2854; // @[utils.scala 60:30]
  wire  _GEN_3047 = branchOps_passed ? _GEN_2535 : _GEN_2855; // @[utils.scala 60:30]
  wire  _GEN_3048 = branchOps_passed ? _GEN_2536 : _GEN_2856; // @[utils.scala 60:30]
  wire  _GEN_3049 = branchOps_passed ? _GEN_2537 : _GEN_2857; // @[utils.scala 60:30]
  wire  _GEN_3050 = branchOps_passed ? _GEN_2538 : _GEN_2858; // @[utils.scala 60:30]
  wire  _GEN_3051 = branchOps_passed ? _GEN_2539 : _GEN_2859; // @[utils.scala 60:30]
  wire  _GEN_3052 = branchOps_passed ? _GEN_2540 : _GEN_2860; // @[utils.scala 60:30]
  wire  _GEN_3053 = branchOps_passed ? _GEN_2541 : _GEN_2861; // @[utils.scala 60:30]
  wire  _GEN_3054 = branchOps_passed ? _GEN_2542 : _GEN_2862; // @[utils.scala 60:30]
  wire  _GEN_3055 = branchOps_passed ? _GEN_2543 : _GEN_2863; // @[utils.scala 60:30]
  wire  _GEN_3056 = branchOps_passed ? _GEN_2544 : _GEN_2864; // @[utils.scala 60:30]
  wire  _GEN_3057 = branchOps_passed ? _GEN_2545 : _GEN_2865; // @[utils.scala 60:30]
  wire  _GEN_3058 = branchOps_passed ? _GEN_2546 : _GEN_2866; // @[utils.scala 60:30]
  wire  _GEN_3059 = branchOps_passed ? _GEN_2547 : _GEN_2867; // @[utils.scala 60:30]
  wire  _GEN_3060 = branchOps_passed ? _GEN_2548 : _GEN_2868; // @[utils.scala 60:30]
  wire  _GEN_3061 = branchOps_passed ? _GEN_2549 : _GEN_2869; // @[utils.scala 60:30]
  wire  _GEN_3062 = branchOps_passed ? _GEN_2550 : _GEN_2870; // @[utils.scala 60:30]
  wire  _GEN_3063 = branchOps_passed ? _GEN_2551 : _GEN_2871; // @[utils.scala 60:30]
  wire  _GEN_3064 = branchOps_passed ? _GEN_2552 : _GEN_2872; // @[utils.scala 60:30]
  wire  _GEN_3065 = branchOps_passed ? _GEN_2553 : _GEN_2873; // @[utils.scala 60:30]
  wire  _GEN_3066 = branchOps_passed ? _GEN_2554 : _GEN_2874; // @[utils.scala 60:30]
  wire  _GEN_3067 = branchOps_passed ? _GEN_2555 : _GEN_2875; // @[utils.scala 60:30]
  wire  _GEN_3068 = branchOps_passed ? _GEN_2556 : _GEN_2876; // @[utils.scala 60:30]
  wire  _GEN_3069 = branchOps_passed ? _GEN_2557 : _GEN_2877; // @[utils.scala 60:30]
  wire  _GEN_3070 = branchOps_passed ? _GEN_2558 : _GEN_2878; // @[utils.scala 60:30]
  wire  _GEN_3071 = branchOps_passed ? _GEN_2559 : _GEN_2879; // @[utils.scala 60:30]
  wire  _GEN_3072 = branchOps_passed ? _GEN_2560 : _GEN_2880; // @[utils.scala 60:30]
  wire  _GEN_3073 = branchOps_passed ? _GEN_2561 : _GEN_2881; // @[utils.scala 60:30]
  wire  _GEN_3074 = branchOps_passed ? _GEN_2562 : _GEN_2882; // @[utils.scala 60:30]
  wire  _GEN_3075 = branchOps_passed ? _GEN_2563 : _GEN_2883; // @[utils.scala 60:30]
  wire  _GEN_3076 = branchOps_passed ? _GEN_2564 : _GEN_2884; // @[utils.scala 60:30]
  wire  _GEN_3077 = branchOps_passed ? _GEN_2565 : _GEN_2885; // @[utils.scala 60:30]
  wire  _GEN_3078 = branchOps_passed ? _GEN_2566 : _GEN_2886; // @[utils.scala 60:30]
  wire  _GEN_3079 = branchOps_passed ? _GEN_2567 : _GEN_2887; // @[utils.scala 60:30]
  wire  _GEN_3080 = branchOps_passed ? _GEN_2568 : _GEN_2888; // @[utils.scala 60:30]
  wire  _GEN_3081 = branchOps_passed ? _GEN_2569 : _GEN_2889; // @[utils.scala 60:30]
  wire  _GEN_3082 = branchOps_passed ? _GEN_2570 : _GEN_2890; // @[utils.scala 60:30]
  wire  _GEN_3083 = branchOps_passed ? _GEN_2571 : _GEN_2891; // @[utils.scala 60:30]
  wire  _GEN_3084 = branchOps_passed ? _GEN_2572 : _GEN_2892; // @[utils.scala 60:30]
  wire  _GEN_3085 = branchOps_passed ? _GEN_2573 : _GEN_2893; // @[utils.scala 60:30]
  wire  _GEN_3086 = branchOps_passed ? _GEN_2574 : _GEN_2894; // @[utils.scala 60:30]
  wire  _GEN_3087 = branchOps_passed ? _GEN_2575 : _GEN_2895; // @[utils.scala 60:30]
  wire  _GEN_3088 = branchOps_passed ? _GEN_2576 : _GEN_2896; // @[utils.scala 60:30]
  wire  _GEN_3089 = branchOps_passed ? _GEN_2577 : _GEN_2897; // @[utils.scala 60:30]
  wire  _GEN_3090 = branchOps_passed ? _GEN_2578 : _GEN_2898; // @[utils.scala 60:30]
  wire  _GEN_3091 = branchOps_passed ? _GEN_2579 : _GEN_2899; // @[utils.scala 60:30]
  wire  _GEN_3092 = branchOps_passed ? _GEN_2580 : _GEN_2900; // @[utils.scala 60:30]
  wire  _GEN_3093 = branchOps_passed ? _GEN_2581 : _GEN_2901; // @[utils.scala 60:30]
  wire  _GEN_3094 = branchOps_passed ? _GEN_2582 : _GEN_2902; // @[utils.scala 60:30]
  wire  _GEN_3095 = branchOps_passed ? _GEN_2583 : _GEN_2903; // @[utils.scala 60:30]
  wire  _GEN_3096 = branchOps_passed ? _GEN_2584 : _GEN_2904; // @[utils.scala 60:30]
  wire  _GEN_3097 = branchOps_passed ? _GEN_2585 : _GEN_2905; // @[utils.scala 60:30]
  wire  _GEN_3098 = branchOps_passed ? _GEN_2586 : _GEN_2906; // @[utils.scala 60:30]
  wire  _GEN_3099 = branchOps_passed ? _GEN_2587 : _GEN_2907; // @[utils.scala 60:30]
  wire  _GEN_3100 = branchOps_passed ? _GEN_2588 : _GEN_2908; // @[utils.scala 60:30]
  wire  _GEN_3101 = branchOps_passed ? _GEN_2589 : _GEN_2909; // @[utils.scala 60:30]
  wire [4:0] _GEN_3230 = branchOps_valid ? _GEN_2974 : _GEN_2398; // @[utils.scala 59:26]
  wire [4:0] _GEN_3231 = branchOps_valid ? _GEN_2975 : _GEN_2399; // @[utils.scala 59:26]
  wire [4:0] _GEN_3232 = branchOps_valid ? _GEN_2976 : _GEN_2400; // @[utils.scala 59:26]
  wire [4:0] _GEN_3233 = branchOps_valid ? _GEN_2977 : _GEN_2401; // @[utils.scala 59:26]
  wire [4:0] _GEN_3234 = branchOps_valid ? _GEN_2978 : _GEN_2402; // @[utils.scala 59:26]
  wire [4:0] _GEN_3235 = branchOps_valid ? _GEN_2979 : _GEN_2403; // @[utils.scala 59:26]
  wire [4:0] _GEN_3236 = branchOps_valid ? _GEN_2980 : _GEN_2404; // @[utils.scala 59:26]
  wire [4:0] _GEN_3237 = branchOps_valid ? _GEN_2981 : _GEN_2405; // @[utils.scala 59:26]
  wire [4:0] _GEN_3238 = branchOps_valid ? _GEN_2982 : _GEN_2406; // @[utils.scala 59:26]
  wire [4:0] _GEN_3239 = branchOps_valid ? _GEN_2983 : _GEN_2407; // @[utils.scala 59:26]
  wire [4:0] _GEN_3240 = branchOps_valid ? _GEN_2984 : _GEN_2408; // @[utils.scala 59:26]
  wire [4:0] _GEN_3241 = branchOps_valid ? _GEN_2985 : _GEN_2409; // @[utils.scala 59:26]
  wire [4:0] _GEN_3242 = branchOps_valid ? _GEN_2986 : _GEN_2410; // @[utils.scala 59:26]
  wire [4:0] _GEN_3243 = branchOps_valid ? _GEN_2987 : _GEN_2411; // @[utils.scala 59:26]
  wire [4:0] _GEN_3244 = branchOps_valid ? _GEN_2988 : _GEN_2412; // @[utils.scala 59:26]
  wire [4:0] _GEN_3245 = branchOps_valid ? _GEN_2989 : _GEN_2413; // @[utils.scala 59:26]
  wire [4:0] _GEN_3246 = branchOps_valid ? _GEN_2990 : _GEN_2414; // @[utils.scala 59:26]
  wire [4:0] _GEN_3247 = branchOps_valid ? _GEN_2991 : _GEN_2415; // @[utils.scala 59:26]
  wire [4:0] _GEN_3248 = branchOps_valid ? _GEN_2992 : _GEN_2416; // @[utils.scala 59:26]
  wire [4:0] _GEN_3249 = branchOps_valid ? _GEN_2993 : _GEN_2417; // @[utils.scala 59:26]
  wire [4:0] _GEN_3250 = branchOps_valid ? _GEN_2994 : _GEN_2418; // @[utils.scala 59:26]
  wire [4:0] _GEN_3251 = branchOps_valid ? _GEN_2995 : _GEN_2419; // @[utils.scala 59:26]
  wire [4:0] _GEN_3252 = branchOps_valid ? _GEN_2996 : _GEN_2420; // @[utils.scala 59:26]
  wire [4:0] _GEN_3253 = branchOps_valid ? _GEN_2997 : _GEN_2421; // @[utils.scala 59:26]
  wire [4:0] _GEN_3254 = branchOps_valid ? _GEN_2998 : _GEN_2422; // @[utils.scala 59:26]
  wire [4:0] _GEN_3255 = branchOps_valid ? _GEN_2999 : _GEN_2423; // @[utils.scala 59:26]
  wire [4:0] _GEN_3256 = branchOps_valid ? _GEN_3000 : _GEN_2424; // @[utils.scala 59:26]
  wire [4:0] _GEN_3257 = branchOps_valid ? _GEN_3001 : _GEN_2425; // @[utils.scala 59:26]
  wire [4:0] _GEN_3258 = branchOps_valid ? _GEN_3002 : _GEN_2426; // @[utils.scala 59:26]
  wire [4:0] _GEN_3259 = branchOps_valid ? _GEN_3003 : _GEN_2427; // @[utils.scala 59:26]
  wire [4:0] _GEN_3260 = branchOps_valid ? _GEN_3004 : _GEN_2428; // @[utils.scala 59:26]
  wire [4:0] _GEN_3261 = branchOps_valid ? _GEN_3005 : _GEN_2429; // @[utils.scala 59:26]
  wire [4:0] _GEN_3262 = branchOps_valid ? _GEN_3006 : _GEN_2430; // @[utils.scala 59:26]
  wire [4:0] _GEN_3263 = branchOps_valid ? _GEN_3007 : _GEN_2431; // @[utils.scala 59:26]
  wire [4:0] _GEN_3264 = branchOps_valid ? _GEN_3008 : _GEN_2432; // @[utils.scala 59:26]
  wire [4:0] _GEN_3265 = branchOps_valid ? _GEN_3009 : _GEN_2433; // @[utils.scala 59:26]
  wire [4:0] _GEN_3266 = branchOps_valid ? _GEN_3010 : _GEN_2434; // @[utils.scala 59:26]
  wire [4:0] _GEN_3267 = branchOps_valid ? _GEN_3011 : _GEN_2435; // @[utils.scala 59:26]
  wire [4:0] _GEN_3268 = branchOps_valid ? _GEN_3012 : _GEN_2436; // @[utils.scala 59:26]
  wire [4:0] _GEN_3269 = branchOps_valid ? _GEN_3013 : _GEN_2437; // @[utils.scala 59:26]
  wire [4:0] _GEN_3270 = branchOps_valid ? _GEN_3014 : _GEN_2438; // @[utils.scala 59:26]
  wire [4:0] _GEN_3271 = branchOps_valid ? _GEN_3015 : _GEN_2439; // @[utils.scala 59:26]
  wire [4:0] _GEN_3272 = branchOps_valid ? _GEN_3016 : _GEN_2440; // @[utils.scala 59:26]
  wire [4:0] _GEN_3273 = branchOps_valid ? _GEN_3017 : _GEN_2441; // @[utils.scala 59:26]
  wire [4:0] _GEN_3274 = branchOps_valid ? _GEN_3018 : _GEN_2442; // @[utils.scala 59:26]
  wire [4:0] _GEN_3275 = branchOps_valid ? _GEN_3019 : _GEN_2443; // @[utils.scala 59:26]
  wire [4:0] _GEN_3276 = branchOps_valid ? _GEN_3020 : _GEN_2444; // @[utils.scala 59:26]
  wire [4:0] _GEN_3277 = branchOps_valid ? _GEN_3021 : _GEN_2445; // @[utils.scala 59:26]
  wire [4:0] _GEN_3278 = branchOps_valid ? _GEN_3022 : _GEN_2446; // @[utils.scala 59:26]
  wire [4:0] _GEN_3279 = branchOps_valid ? _GEN_3023 : _GEN_2447; // @[utils.scala 59:26]
  wire [4:0] _GEN_3280 = branchOps_valid ? _GEN_3024 : _GEN_2448; // @[utils.scala 59:26]
  wire [4:0] _GEN_3281 = branchOps_valid ? _GEN_3025 : _GEN_2449; // @[utils.scala 59:26]
  wire [4:0] _GEN_3282 = branchOps_valid ? _GEN_3026 : _GEN_2450; // @[utils.scala 59:26]
  wire [4:0] _GEN_3283 = branchOps_valid ? _GEN_3027 : _GEN_2451; // @[utils.scala 59:26]
  wire [4:0] _GEN_3284 = branchOps_valid ? _GEN_3028 : _GEN_2452; // @[utils.scala 59:26]
  wire [4:0] _GEN_3285 = branchOps_valid ? _GEN_3029 : _GEN_2453; // @[utils.scala 59:26]
  wire [4:0] _GEN_3286 = branchOps_valid ? _GEN_3030 : _GEN_2454; // @[utils.scala 59:26]
  wire [4:0] _GEN_3287 = branchOps_valid ? _GEN_3031 : _GEN_2455; // @[utils.scala 59:26]
  wire [4:0] _GEN_3288 = branchOps_valid ? _GEN_3032 : _GEN_2456; // @[utils.scala 59:26]
  wire [4:0] _GEN_3289 = branchOps_valid ? _GEN_3033 : _GEN_2457; // @[utils.scala 59:26]
  wire [4:0] _GEN_3290 = branchOps_valid ? _GEN_3034 : _GEN_2458; // @[utils.scala 59:26]
  wire [4:0] _GEN_3291 = branchOps_valid ? _GEN_3035 : _GEN_2459; // @[utils.scala 59:26]
  wire [4:0] _GEN_3292 = branchOps_valid ? _GEN_3036 : _GEN_2460; // @[utils.scala 59:26]
  wire [4:0] _GEN_3293 = branchOps_valid ? _GEN_3037 : _GEN_2461; // @[utils.scala 59:26]
  wire  _GEN_3294 = branchOps_valid ? _GEN_3038 : _GEN_2526; // @[utils.scala 59:26]
  wire  _GEN_3295 = branchOps_valid ? _GEN_3039 : _GEN_2527; // @[utils.scala 59:26]
  wire  _GEN_3296 = branchOps_valid ? _GEN_3040 : _GEN_2528; // @[utils.scala 59:26]
  wire  _GEN_3297 = branchOps_valid ? _GEN_3041 : _GEN_2529; // @[utils.scala 59:26]
  wire  _GEN_3298 = branchOps_valid ? _GEN_3042 : _GEN_2530; // @[utils.scala 59:26]
  wire  _GEN_3299 = branchOps_valid ? _GEN_3043 : _GEN_2531; // @[utils.scala 59:26]
  wire  _GEN_3300 = branchOps_valid ? _GEN_3044 : _GEN_2532; // @[utils.scala 59:26]
  wire  _GEN_3301 = branchOps_valid ? _GEN_3045 : _GEN_2533; // @[utils.scala 59:26]
  wire  _GEN_3302 = branchOps_valid ? _GEN_3046 : _GEN_2534; // @[utils.scala 59:26]
  wire  _GEN_3303 = branchOps_valid ? _GEN_3047 : _GEN_2535; // @[utils.scala 59:26]
  wire  _GEN_3304 = branchOps_valid ? _GEN_3048 : _GEN_2536; // @[utils.scala 59:26]
  wire  _GEN_3305 = branchOps_valid ? _GEN_3049 : _GEN_2537; // @[utils.scala 59:26]
  wire  _GEN_3306 = branchOps_valid ? _GEN_3050 : _GEN_2538; // @[utils.scala 59:26]
  wire  _GEN_3307 = branchOps_valid ? _GEN_3051 : _GEN_2539; // @[utils.scala 59:26]
  wire  _GEN_3308 = branchOps_valid ? _GEN_3052 : _GEN_2540; // @[utils.scala 59:26]
  wire  _GEN_3309 = branchOps_valid ? _GEN_3053 : _GEN_2541; // @[utils.scala 59:26]
  wire  _GEN_3310 = branchOps_valid ? _GEN_3054 : _GEN_2542; // @[utils.scala 59:26]
  wire  _GEN_3311 = branchOps_valid ? _GEN_3055 : _GEN_2543; // @[utils.scala 59:26]
  wire  _GEN_3312 = branchOps_valid ? _GEN_3056 : _GEN_2544; // @[utils.scala 59:26]
  wire  _GEN_3313 = branchOps_valid ? _GEN_3057 : _GEN_2545; // @[utils.scala 59:26]
  wire  _GEN_3314 = branchOps_valid ? _GEN_3058 : _GEN_2546; // @[utils.scala 59:26]
  wire  _GEN_3315 = branchOps_valid ? _GEN_3059 : _GEN_2547; // @[utils.scala 59:26]
  wire  _GEN_3316 = branchOps_valid ? _GEN_3060 : _GEN_2548; // @[utils.scala 59:26]
  wire  _GEN_3317 = branchOps_valid ? _GEN_3061 : _GEN_2549; // @[utils.scala 59:26]
  wire  _GEN_3318 = branchOps_valid ? _GEN_3062 : _GEN_2550; // @[utils.scala 59:26]
  wire  _GEN_3319 = branchOps_valid ? _GEN_3063 : _GEN_2551; // @[utils.scala 59:26]
  wire  _GEN_3320 = branchOps_valid ? _GEN_3064 : _GEN_2552; // @[utils.scala 59:26]
  wire  _GEN_3321 = branchOps_valid ? _GEN_3065 : _GEN_2553; // @[utils.scala 59:26]
  wire  _GEN_3322 = branchOps_valid ? _GEN_3066 : _GEN_2554; // @[utils.scala 59:26]
  wire  _GEN_3323 = branchOps_valid ? _GEN_3067 : _GEN_2555; // @[utils.scala 59:26]
  wire  _GEN_3324 = branchOps_valid ? _GEN_3068 : _GEN_2556; // @[utils.scala 59:26]
  wire  _GEN_3325 = branchOps_valid ? _GEN_3069 : _GEN_2557; // @[utils.scala 59:26]
  wire  _GEN_3326 = branchOps_valid ? _GEN_3070 : _GEN_2558; // @[utils.scala 59:26]
  wire  _GEN_3327 = branchOps_valid ? _GEN_3071 : _GEN_2559; // @[utils.scala 59:26]
  wire  _GEN_3328 = branchOps_valid ? _GEN_3072 : _GEN_2560; // @[utils.scala 59:26]
  wire  _GEN_3329 = branchOps_valid ? _GEN_3073 : _GEN_2561; // @[utils.scala 59:26]
  wire  _GEN_3330 = branchOps_valid ? _GEN_3074 : _GEN_2562; // @[utils.scala 59:26]
  wire  _GEN_3331 = branchOps_valid ? _GEN_3075 : _GEN_2563; // @[utils.scala 59:26]
  wire  _GEN_3332 = branchOps_valid ? _GEN_3076 : _GEN_2564; // @[utils.scala 59:26]
  wire  _GEN_3333 = branchOps_valid ? _GEN_3077 : _GEN_2565; // @[utils.scala 59:26]
  wire  _GEN_3334 = branchOps_valid ? _GEN_3078 : _GEN_2566; // @[utils.scala 59:26]
  wire  _GEN_3335 = branchOps_valid ? _GEN_3079 : _GEN_2567; // @[utils.scala 59:26]
  wire  _GEN_3336 = branchOps_valid ? _GEN_3080 : _GEN_2568; // @[utils.scala 59:26]
  wire  _GEN_3337 = branchOps_valid ? _GEN_3081 : _GEN_2569; // @[utils.scala 59:26]
  wire  _GEN_3338 = branchOps_valid ? _GEN_3082 : _GEN_2570; // @[utils.scala 59:26]
  wire  _GEN_3339 = branchOps_valid ? _GEN_3083 : _GEN_2571; // @[utils.scala 59:26]
  wire  _GEN_3340 = branchOps_valid ? _GEN_3084 : _GEN_2572; // @[utils.scala 59:26]
  wire  _GEN_3341 = branchOps_valid ? _GEN_3085 : _GEN_2573; // @[utils.scala 59:26]
  wire  _GEN_3342 = branchOps_valid ? _GEN_3086 : _GEN_2574; // @[utils.scala 59:26]
  wire  _GEN_3343 = branchOps_valid ? _GEN_3087 : _GEN_2575; // @[utils.scala 59:26]
  wire  _GEN_3344 = branchOps_valid ? _GEN_3088 : _GEN_2576; // @[utils.scala 59:26]
  wire  _GEN_3345 = branchOps_valid ? _GEN_3089 : _GEN_2577; // @[utils.scala 59:26]
  wire  _GEN_3346 = branchOps_valid ? _GEN_3090 : _GEN_2578; // @[utils.scala 59:26]
  wire  _GEN_3347 = branchOps_valid ? _GEN_3091 : _GEN_2579; // @[utils.scala 59:26]
  wire  _GEN_3348 = branchOps_valid ? _GEN_3092 : _GEN_2580; // @[utils.scala 59:26]
  wire  _GEN_3349 = branchOps_valid ? _GEN_3093 : _GEN_2581; // @[utils.scala 59:26]
  wire  _GEN_3350 = branchOps_valid ? _GEN_3094 : _GEN_2582; // @[utils.scala 59:26]
  wire  _GEN_3351 = branchOps_valid ? _GEN_3095 : _GEN_2583; // @[utils.scala 59:26]
  wire  _GEN_3352 = branchOps_valid ? _GEN_3096 : _GEN_2584; // @[utils.scala 59:26]
  wire  _GEN_3353 = branchOps_valid ? _GEN_3097 : _GEN_2585; // @[utils.scala 59:26]
  wire  _GEN_3354 = branchOps_valid ? _GEN_3098 : _GEN_2586; // @[utils.scala 59:26]
  wire  _GEN_3355 = branchOps_valid ? _GEN_3099 : _GEN_2587; // @[utils.scala 59:26]
  wire  _GEN_3356 = branchOps_valid ? _GEN_3100 : _GEN_2588; // @[utils.scala 59:26]
  wire  _GEN_3357 = branchOps_valid ? _GEN_3101 : _GEN_2589; // @[utils.scala 59:26]
  wire [4:0] _GEN_3358 = incrWrite ? _GEN_3230 : _GEN_1182; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3359 = incrWrite ? _GEN_3231 : _GEN_1183; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3360 = incrWrite ? _GEN_3232 : _GEN_1184; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3361 = incrWrite ? _GEN_3233 : _GEN_1185; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3362 = incrWrite ? _GEN_3234 : _GEN_1186; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3363 = incrWrite ? _GEN_3235 : _GEN_1187; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3364 = incrWrite ? _GEN_3236 : _GEN_1188; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3365 = incrWrite ? _GEN_3237 : _GEN_1189; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3366 = incrWrite ? _GEN_3238 : _GEN_1190; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3367 = incrWrite ? _GEN_3239 : _GEN_1191; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3368 = incrWrite ? _GEN_3240 : _GEN_1192; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3369 = incrWrite ? _GEN_3241 : _GEN_1193; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3370 = incrWrite ? _GEN_3242 : _GEN_1194; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3371 = incrWrite ? _GEN_3243 : _GEN_1195; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3372 = incrWrite ? _GEN_3244 : _GEN_1196; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3373 = incrWrite ? _GEN_3245 : _GEN_1197; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3374 = incrWrite ? _GEN_3246 : _GEN_1198; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3375 = incrWrite ? _GEN_3247 : _GEN_1199; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3376 = incrWrite ? _GEN_3248 : _GEN_1200; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3377 = incrWrite ? _GEN_3249 : _GEN_1201; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3378 = incrWrite ? _GEN_3250 : _GEN_1202; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3379 = incrWrite ? _GEN_3251 : _GEN_1203; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3380 = incrWrite ? _GEN_3252 : _GEN_1204; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3381 = incrWrite ? _GEN_3253 : _GEN_1205; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3382 = incrWrite ? _GEN_3254 : _GEN_1206; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3383 = incrWrite ? _GEN_3255 : _GEN_1207; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3384 = incrWrite ? _GEN_3256 : _GEN_1208; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3385 = incrWrite ? _GEN_3257 : _GEN_1209; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3386 = incrWrite ? _GEN_3258 : _GEN_1210; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3387 = incrWrite ? _GEN_3259 : _GEN_1211; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3388 = incrWrite ? _GEN_3260 : _GEN_1212; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3389 = incrWrite ? _GEN_3261 : _GEN_1213; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3390 = incrWrite ? _GEN_3262 : _GEN_1214; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3391 = incrWrite ? _GEN_3263 : _GEN_1215; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3392 = incrWrite ? _GEN_3264 : _GEN_1216; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3393 = incrWrite ? _GEN_3265 : _GEN_1217; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3394 = incrWrite ? _GEN_3266 : _GEN_1218; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3395 = incrWrite ? _GEN_3267 : _GEN_1219; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3396 = incrWrite ? _GEN_3268 : _GEN_1220; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3397 = incrWrite ? _GEN_3269 : _GEN_1221; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3398 = incrWrite ? _GEN_3270 : _GEN_1222; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3399 = incrWrite ? _GEN_3271 : _GEN_1223; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3400 = incrWrite ? _GEN_3272 : _GEN_1224; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3401 = incrWrite ? _GEN_3273 : _GEN_1225; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3402 = incrWrite ? _GEN_3274 : _GEN_1226; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3403 = incrWrite ? _GEN_3275 : _GEN_1227; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3404 = incrWrite ? _GEN_3276 : _GEN_1228; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3405 = incrWrite ? _GEN_3277 : _GEN_1229; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3406 = incrWrite ? _GEN_3278 : _GEN_1230; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3407 = incrWrite ? _GEN_3279 : _GEN_1231; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3408 = incrWrite ? _GEN_3280 : _GEN_1232; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3409 = incrWrite ? _GEN_3281 : _GEN_1233; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3410 = incrWrite ? _GEN_3282 : _GEN_1234; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3411 = incrWrite ? _GEN_3283 : _GEN_1235; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3412 = incrWrite ? _GEN_3284 : _GEN_1236; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3413 = incrWrite ? _GEN_3285 : _GEN_1237; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3414 = incrWrite ? _GEN_3286 : _GEN_1238; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3415 = incrWrite ? _GEN_3287 : _GEN_1239; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3416 = incrWrite ? _GEN_3288 : _GEN_1240; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3417 = incrWrite ? _GEN_3289 : _GEN_1241; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3418 = incrWrite ? _GEN_3290 : _GEN_1242; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3419 = incrWrite ? _GEN_3291 : _GEN_1243; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3420 = incrWrite ? _GEN_3292 : _GEN_1244; // @[fifo.scala 97:16]
  wire [4:0] _GEN_3421 = incrWrite ? _GEN_3293 : _GEN_1245; // @[fifo.scala 97:16]
  wire  _GEN_3422 = incrWrite ? _GEN_3294 : _GEN_1118; // @[fifo.scala 97:16]
  wire  _GEN_3423 = incrWrite ? _GEN_3295 : _GEN_1119; // @[fifo.scala 97:16]
  wire  _GEN_3424 = incrWrite ? _GEN_3296 : _GEN_1120; // @[fifo.scala 97:16]
  wire  _GEN_3425 = incrWrite ? _GEN_3297 : _GEN_1121; // @[fifo.scala 97:16]
  wire  _GEN_3426 = incrWrite ? _GEN_3298 : _GEN_1122; // @[fifo.scala 97:16]
  wire  _GEN_3427 = incrWrite ? _GEN_3299 : _GEN_1123; // @[fifo.scala 97:16]
  wire  _GEN_3428 = incrWrite ? _GEN_3300 : _GEN_1124; // @[fifo.scala 97:16]
  wire  _GEN_3429 = incrWrite ? _GEN_3301 : _GEN_1125; // @[fifo.scala 97:16]
  wire  _GEN_3430 = incrWrite ? _GEN_3302 : _GEN_1126; // @[fifo.scala 97:16]
  wire  _GEN_3431 = incrWrite ? _GEN_3303 : _GEN_1127; // @[fifo.scala 97:16]
  wire  _GEN_3432 = incrWrite ? _GEN_3304 : _GEN_1128; // @[fifo.scala 97:16]
  wire  _GEN_3433 = incrWrite ? _GEN_3305 : _GEN_1129; // @[fifo.scala 97:16]
  wire  _GEN_3434 = incrWrite ? _GEN_3306 : _GEN_1130; // @[fifo.scala 97:16]
  wire  _GEN_3435 = incrWrite ? _GEN_3307 : _GEN_1131; // @[fifo.scala 97:16]
  wire  _GEN_3436 = incrWrite ? _GEN_3308 : _GEN_1132; // @[fifo.scala 97:16]
  wire  _GEN_3437 = incrWrite ? _GEN_3309 : _GEN_1133; // @[fifo.scala 97:16]
  wire  _GEN_3438 = incrWrite ? _GEN_3310 : _GEN_1134; // @[fifo.scala 97:16]
  wire  _GEN_3439 = incrWrite ? _GEN_3311 : _GEN_1135; // @[fifo.scala 97:16]
  wire  _GEN_3440 = incrWrite ? _GEN_3312 : _GEN_1136; // @[fifo.scala 97:16]
  wire  _GEN_3441 = incrWrite ? _GEN_3313 : _GEN_1137; // @[fifo.scala 97:16]
  wire  _GEN_3442 = incrWrite ? _GEN_3314 : _GEN_1138; // @[fifo.scala 97:16]
  wire  _GEN_3443 = incrWrite ? _GEN_3315 : _GEN_1139; // @[fifo.scala 97:16]
  wire  _GEN_3444 = incrWrite ? _GEN_3316 : _GEN_1140; // @[fifo.scala 97:16]
  wire  _GEN_3445 = incrWrite ? _GEN_3317 : _GEN_1141; // @[fifo.scala 97:16]
  wire  _GEN_3446 = incrWrite ? _GEN_3318 : _GEN_1142; // @[fifo.scala 97:16]
  wire  _GEN_3447 = incrWrite ? _GEN_3319 : _GEN_1143; // @[fifo.scala 97:16]
  wire  _GEN_3448 = incrWrite ? _GEN_3320 : _GEN_1144; // @[fifo.scala 97:16]
  wire  _GEN_3449 = incrWrite ? _GEN_3321 : _GEN_1145; // @[fifo.scala 97:16]
  wire  _GEN_3450 = incrWrite ? _GEN_3322 : _GEN_1146; // @[fifo.scala 97:16]
  wire  _GEN_3451 = incrWrite ? _GEN_3323 : _GEN_1147; // @[fifo.scala 97:16]
  wire  _GEN_3452 = incrWrite ? _GEN_3324 : _GEN_1148; // @[fifo.scala 97:16]
  wire  _GEN_3453 = incrWrite ? _GEN_3325 : _GEN_1149; // @[fifo.scala 97:16]
  wire  _GEN_3454 = incrWrite ? _GEN_3326 : _GEN_1150; // @[fifo.scala 97:16]
  wire  _GEN_3455 = incrWrite ? _GEN_3327 : _GEN_1151; // @[fifo.scala 97:16]
  wire  _GEN_3456 = incrWrite ? _GEN_3328 : _GEN_1152; // @[fifo.scala 97:16]
  wire  _GEN_3457 = incrWrite ? _GEN_3329 : _GEN_1153; // @[fifo.scala 97:16]
  wire  _GEN_3458 = incrWrite ? _GEN_3330 : _GEN_1154; // @[fifo.scala 97:16]
  wire  _GEN_3459 = incrWrite ? _GEN_3331 : _GEN_1155; // @[fifo.scala 97:16]
  wire  _GEN_3460 = incrWrite ? _GEN_3332 : _GEN_1156; // @[fifo.scala 97:16]
  wire  _GEN_3461 = incrWrite ? _GEN_3333 : _GEN_1157; // @[fifo.scala 97:16]
  wire  _GEN_3462 = incrWrite ? _GEN_3334 : _GEN_1158; // @[fifo.scala 97:16]
  wire  _GEN_3463 = incrWrite ? _GEN_3335 : _GEN_1159; // @[fifo.scala 97:16]
  wire  _GEN_3464 = incrWrite ? _GEN_3336 : _GEN_1160; // @[fifo.scala 97:16]
  wire  _GEN_3465 = incrWrite ? _GEN_3337 : _GEN_1161; // @[fifo.scala 97:16]
  wire  _GEN_3466 = incrWrite ? _GEN_3338 : _GEN_1162; // @[fifo.scala 97:16]
  wire  _GEN_3467 = incrWrite ? _GEN_3339 : _GEN_1163; // @[fifo.scala 97:16]
  wire  _GEN_3468 = incrWrite ? _GEN_3340 : _GEN_1164; // @[fifo.scala 97:16]
  wire  _GEN_3469 = incrWrite ? _GEN_3341 : _GEN_1165; // @[fifo.scala 97:16]
  wire  _GEN_3470 = incrWrite ? _GEN_3342 : _GEN_1166; // @[fifo.scala 97:16]
  wire  _GEN_3471 = incrWrite ? _GEN_3343 : _GEN_1167; // @[fifo.scala 97:16]
  wire  _GEN_3472 = incrWrite ? _GEN_3344 : _GEN_1168; // @[fifo.scala 97:16]
  wire  _GEN_3473 = incrWrite ? _GEN_3345 : _GEN_1169; // @[fifo.scala 97:16]
  wire  _GEN_3474 = incrWrite ? _GEN_3346 : _GEN_1170; // @[fifo.scala 97:16]
  wire  _GEN_3475 = incrWrite ? _GEN_3347 : _GEN_1171; // @[fifo.scala 97:16]
  wire  _GEN_3476 = incrWrite ? _GEN_3348 : _GEN_1172; // @[fifo.scala 97:16]
  wire  _GEN_3477 = incrWrite ? _GEN_3349 : _GEN_1173; // @[fifo.scala 97:16]
  wire  _GEN_3478 = incrWrite ? _GEN_3350 : _GEN_1174; // @[fifo.scala 97:16]
  wire  _GEN_3479 = incrWrite ? _GEN_3351 : _GEN_1175; // @[fifo.scala 97:16]
  wire  _GEN_3480 = incrWrite ? _GEN_3352 : _GEN_1176; // @[fifo.scala 97:16]
  wire  _GEN_3481 = incrWrite ? _GEN_3353 : _GEN_1177; // @[fifo.scala 97:16]
  wire  _GEN_3482 = incrWrite ? _GEN_3354 : _GEN_1178; // @[fifo.scala 97:16]
  wire  _GEN_3483 = incrWrite ? _GEN_3355 : _GEN_1179; // @[fifo.scala 97:16]
  wire  _GEN_3484 = incrWrite ? _GEN_3356 : _GEN_1180; // @[fifo.scala 97:16]
  wire  _GEN_3485 = incrWrite ? _GEN_3357 : _GEN_1181; // @[fifo.scala 97:16]
  wire [5:0] startPointer = read_ready ? _nextVal_T_2 : readPtr; // @[fifo.scala 102:25]
  wire [5:0] endPointer = writePtr - 6'h1; // @[fifo.scala 103:29]
  wire [4:0] _T_15 = memReg_0_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_16 = |_T_15; // @[fifo.scala 109:63]
  wire [4:0] _memReg_0_branch_mask_T = memReg_0_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _T_22 = memReg_1_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_23 = |_T_22; // @[fifo.scala 109:63]
  wire [4:0] _memReg_1_branch_mask_T = memReg_1_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3492 = |_T_22 ? _memReg_1_branch_mask_T : _GEN_3359; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3493 = _T_23 ? 1'h0 : _GEN_3423; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_29 = memReg_2_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_30 = |_T_29; // @[fifo.scala 109:63]
  wire [4:0] _memReg_2_branch_mask_T = memReg_2_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3498 = |_T_29 ? _memReg_2_branch_mask_T : _GEN_3360; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3499 = _T_30 ? 1'h0 : _GEN_3424; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_36 = memReg_3_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_37 = |_T_36; // @[fifo.scala 109:63]
  wire [4:0] _memReg_3_branch_mask_T = memReg_3_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3504 = |_T_36 ? _memReg_3_branch_mask_T : _GEN_3361; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3505 = _T_37 ? 1'h0 : _GEN_3425; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_43 = memReg_4_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_44 = |_T_43; // @[fifo.scala 109:63]
  wire [4:0] _memReg_4_branch_mask_T = memReg_4_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3510 = |_T_43 ? _memReg_4_branch_mask_T : _GEN_3362; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3511 = _T_44 ? 1'h0 : _GEN_3426; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_50 = memReg_5_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_51 = |_T_50; // @[fifo.scala 109:63]
  wire [4:0] _memReg_5_branch_mask_T = memReg_5_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3516 = |_T_50 ? _memReg_5_branch_mask_T : _GEN_3363; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3517 = _T_51 ? 1'h0 : _GEN_3427; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_57 = memReg_6_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_58 = |_T_57; // @[fifo.scala 109:63]
  wire [4:0] _memReg_6_branch_mask_T = memReg_6_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3522 = |_T_57 ? _memReg_6_branch_mask_T : _GEN_3364; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3523 = _T_58 ? 1'h0 : _GEN_3428; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_64 = memReg_7_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_65 = |_T_64; // @[fifo.scala 109:63]
  wire [4:0] _memReg_7_branch_mask_T = memReg_7_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3528 = |_T_64 ? _memReg_7_branch_mask_T : _GEN_3365; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3529 = _T_65 ? 1'h0 : _GEN_3429; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_71 = memReg_8_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_72 = |_T_71; // @[fifo.scala 109:63]
  wire [4:0] _memReg_8_branch_mask_T = memReg_8_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3534 = |_T_71 ? _memReg_8_branch_mask_T : _GEN_3366; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3535 = _T_72 ? 1'h0 : _GEN_3430; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_78 = memReg_9_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_79 = |_T_78; // @[fifo.scala 109:63]
  wire [4:0] _memReg_9_branch_mask_T = memReg_9_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3540 = |_T_78 ? _memReg_9_branch_mask_T : _GEN_3367; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3541 = _T_79 ? 1'h0 : _GEN_3431; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_85 = memReg_10_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_86 = |_T_85; // @[fifo.scala 109:63]
  wire [4:0] _memReg_10_branch_mask_T = memReg_10_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3546 = |_T_85 ? _memReg_10_branch_mask_T : _GEN_3368; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3547 = _T_86 ? 1'h0 : _GEN_3432; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_92 = memReg_11_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_93 = |_T_92; // @[fifo.scala 109:63]
  wire [4:0] _memReg_11_branch_mask_T = memReg_11_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3552 = |_T_92 ? _memReg_11_branch_mask_T : _GEN_3369; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3553 = _T_93 ? 1'h0 : _GEN_3433; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_99 = memReg_12_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_100 = |_T_99; // @[fifo.scala 109:63]
  wire [4:0] _memReg_12_branch_mask_T = memReg_12_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3558 = |_T_99 ? _memReg_12_branch_mask_T : _GEN_3370; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3559 = _T_100 ? 1'h0 : _GEN_3434; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_106 = memReg_13_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_107 = |_T_106; // @[fifo.scala 109:63]
  wire [4:0] _memReg_13_branch_mask_T = memReg_13_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3564 = |_T_106 ? _memReg_13_branch_mask_T : _GEN_3371; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3565 = _T_107 ? 1'h0 : _GEN_3435; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_113 = memReg_14_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_114 = |_T_113; // @[fifo.scala 109:63]
  wire [4:0] _memReg_14_branch_mask_T = memReg_14_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3570 = |_T_113 ? _memReg_14_branch_mask_T : _GEN_3372; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3571 = _T_114 ? 1'h0 : _GEN_3436; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_120 = memReg_15_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_121 = |_T_120; // @[fifo.scala 109:63]
  wire [4:0] _memReg_15_branch_mask_T = memReg_15_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3576 = |_T_120 ? _memReg_15_branch_mask_T : _GEN_3373; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3577 = _T_121 ? 1'h0 : _GEN_3437; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_127 = memReg_16_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_128 = |_T_127; // @[fifo.scala 109:63]
  wire [4:0] _memReg_16_branch_mask_T = memReg_16_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3582 = |_T_127 ? _memReg_16_branch_mask_T : _GEN_3374; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3583 = _T_128 ? 1'h0 : _GEN_3438; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_134 = memReg_17_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_135 = |_T_134; // @[fifo.scala 109:63]
  wire [4:0] _memReg_17_branch_mask_T = memReg_17_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3588 = |_T_134 ? _memReg_17_branch_mask_T : _GEN_3375; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3589 = _T_135 ? 1'h0 : _GEN_3439; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_141 = memReg_18_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_142 = |_T_141; // @[fifo.scala 109:63]
  wire [4:0] _memReg_18_branch_mask_T = memReg_18_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3594 = |_T_141 ? _memReg_18_branch_mask_T : _GEN_3376; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3595 = _T_142 ? 1'h0 : _GEN_3440; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_148 = memReg_19_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_149 = |_T_148; // @[fifo.scala 109:63]
  wire [4:0] _memReg_19_branch_mask_T = memReg_19_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3600 = |_T_148 ? _memReg_19_branch_mask_T : _GEN_3377; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3601 = _T_149 ? 1'h0 : _GEN_3441; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_155 = memReg_20_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_156 = |_T_155; // @[fifo.scala 109:63]
  wire [4:0] _memReg_20_branch_mask_T = memReg_20_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3606 = |_T_155 ? _memReg_20_branch_mask_T : _GEN_3378; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3607 = _T_156 ? 1'h0 : _GEN_3442; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_162 = memReg_21_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_163 = |_T_162; // @[fifo.scala 109:63]
  wire [4:0] _memReg_21_branch_mask_T = memReg_21_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3612 = |_T_162 ? _memReg_21_branch_mask_T : _GEN_3379; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3613 = _T_163 ? 1'h0 : _GEN_3443; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_169 = memReg_22_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_170 = |_T_169; // @[fifo.scala 109:63]
  wire [4:0] _memReg_22_branch_mask_T = memReg_22_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3618 = |_T_169 ? _memReg_22_branch_mask_T : _GEN_3380; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3619 = _T_170 ? 1'h0 : _GEN_3444; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_176 = memReg_23_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_177 = |_T_176; // @[fifo.scala 109:63]
  wire [4:0] _memReg_23_branch_mask_T = memReg_23_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3624 = |_T_176 ? _memReg_23_branch_mask_T : _GEN_3381; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3625 = _T_177 ? 1'h0 : _GEN_3445; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_183 = memReg_24_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_184 = |_T_183; // @[fifo.scala 109:63]
  wire [4:0] _memReg_24_branch_mask_T = memReg_24_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3630 = |_T_183 ? _memReg_24_branch_mask_T : _GEN_3382; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3631 = _T_184 ? 1'h0 : _GEN_3446; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_190 = memReg_25_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_191 = |_T_190; // @[fifo.scala 109:63]
  wire [4:0] _memReg_25_branch_mask_T = memReg_25_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3636 = |_T_190 ? _memReg_25_branch_mask_T : _GEN_3383; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3637 = _T_191 ? 1'h0 : _GEN_3447; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_197 = memReg_26_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_198 = |_T_197; // @[fifo.scala 109:63]
  wire [4:0] _memReg_26_branch_mask_T = memReg_26_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3642 = |_T_197 ? _memReg_26_branch_mask_T : _GEN_3384; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3643 = _T_198 ? 1'h0 : _GEN_3448; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_204 = memReg_27_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_205 = |_T_204; // @[fifo.scala 109:63]
  wire [4:0] _memReg_27_branch_mask_T = memReg_27_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3648 = |_T_204 ? _memReg_27_branch_mask_T : _GEN_3385; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3649 = _T_205 ? 1'h0 : _GEN_3449; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_211 = memReg_28_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_212 = |_T_211; // @[fifo.scala 109:63]
  wire [4:0] _memReg_28_branch_mask_T = memReg_28_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3654 = |_T_211 ? _memReg_28_branch_mask_T : _GEN_3386; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3655 = _T_212 ? 1'h0 : _GEN_3450; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_218 = memReg_29_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_219 = |_T_218; // @[fifo.scala 109:63]
  wire [4:0] _memReg_29_branch_mask_T = memReg_29_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3660 = |_T_218 ? _memReg_29_branch_mask_T : _GEN_3387; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3661 = _T_219 ? 1'h0 : _GEN_3451; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_225 = memReg_30_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_226 = |_T_225; // @[fifo.scala 109:63]
  wire [4:0] _memReg_30_branch_mask_T = memReg_30_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3666 = |_T_225 ? _memReg_30_branch_mask_T : _GEN_3388; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3667 = _T_226 ? 1'h0 : _GEN_3452; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_232 = memReg_31_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_233 = |_T_232; // @[fifo.scala 109:63]
  wire [4:0] _memReg_31_branch_mask_T = memReg_31_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3672 = |_T_232 ? _memReg_31_branch_mask_T : _GEN_3389; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3673 = _T_233 ? 1'h0 : _GEN_3453; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_239 = memReg_32_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_240 = |_T_239; // @[fifo.scala 109:63]
  wire [4:0] _memReg_32_branch_mask_T = memReg_32_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3678 = |_T_239 ? _memReg_32_branch_mask_T : _GEN_3390; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3679 = _T_240 ? 1'h0 : _GEN_3454; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_246 = memReg_33_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_247 = |_T_246; // @[fifo.scala 109:63]
  wire [4:0] _memReg_33_branch_mask_T = memReg_33_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3684 = |_T_246 ? _memReg_33_branch_mask_T : _GEN_3391; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3685 = _T_247 ? 1'h0 : _GEN_3455; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_253 = memReg_34_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_254 = |_T_253; // @[fifo.scala 109:63]
  wire [4:0] _memReg_34_branch_mask_T = memReg_34_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3690 = |_T_253 ? _memReg_34_branch_mask_T : _GEN_3392; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3691 = _T_254 ? 1'h0 : _GEN_3456; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_260 = memReg_35_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_261 = |_T_260; // @[fifo.scala 109:63]
  wire [4:0] _memReg_35_branch_mask_T = memReg_35_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3696 = |_T_260 ? _memReg_35_branch_mask_T : _GEN_3393; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3697 = _T_261 ? 1'h0 : _GEN_3457; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_267 = memReg_36_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_268 = |_T_267; // @[fifo.scala 109:63]
  wire [4:0] _memReg_36_branch_mask_T = memReg_36_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3702 = |_T_267 ? _memReg_36_branch_mask_T : _GEN_3394; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3703 = _T_268 ? 1'h0 : _GEN_3458; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_274 = memReg_37_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_275 = |_T_274; // @[fifo.scala 109:63]
  wire [4:0] _memReg_37_branch_mask_T = memReg_37_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3708 = |_T_274 ? _memReg_37_branch_mask_T : _GEN_3395; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3709 = _T_275 ? 1'h0 : _GEN_3459; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_281 = memReg_38_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_282 = |_T_281; // @[fifo.scala 109:63]
  wire [4:0] _memReg_38_branch_mask_T = memReg_38_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3714 = |_T_281 ? _memReg_38_branch_mask_T : _GEN_3396; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3715 = _T_282 ? 1'h0 : _GEN_3460; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_288 = memReg_39_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_289 = |_T_288; // @[fifo.scala 109:63]
  wire [4:0] _memReg_39_branch_mask_T = memReg_39_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3720 = |_T_288 ? _memReg_39_branch_mask_T : _GEN_3397; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3721 = _T_289 ? 1'h0 : _GEN_3461; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_295 = memReg_40_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_296 = |_T_295; // @[fifo.scala 109:63]
  wire [4:0] _memReg_40_branch_mask_T = memReg_40_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3726 = |_T_295 ? _memReg_40_branch_mask_T : _GEN_3398; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3727 = _T_296 ? 1'h0 : _GEN_3462; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_302 = memReg_41_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_303 = |_T_302; // @[fifo.scala 109:63]
  wire [4:0] _memReg_41_branch_mask_T = memReg_41_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3732 = |_T_302 ? _memReg_41_branch_mask_T : _GEN_3399; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3733 = _T_303 ? 1'h0 : _GEN_3463; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_309 = memReg_42_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_310 = |_T_309; // @[fifo.scala 109:63]
  wire [4:0] _memReg_42_branch_mask_T = memReg_42_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3738 = |_T_309 ? _memReg_42_branch_mask_T : _GEN_3400; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3739 = _T_310 ? 1'h0 : _GEN_3464; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_316 = memReg_43_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_317 = |_T_316; // @[fifo.scala 109:63]
  wire [4:0] _memReg_43_branch_mask_T = memReg_43_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3744 = |_T_316 ? _memReg_43_branch_mask_T : _GEN_3401; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3745 = _T_317 ? 1'h0 : _GEN_3465; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_323 = memReg_44_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_324 = |_T_323; // @[fifo.scala 109:63]
  wire [4:0] _memReg_44_branch_mask_T = memReg_44_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3750 = |_T_323 ? _memReg_44_branch_mask_T : _GEN_3402; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3751 = _T_324 ? 1'h0 : _GEN_3466; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_330 = memReg_45_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_331 = |_T_330; // @[fifo.scala 109:63]
  wire [4:0] _memReg_45_branch_mask_T = memReg_45_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3756 = |_T_330 ? _memReg_45_branch_mask_T : _GEN_3403; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3757 = _T_331 ? 1'h0 : _GEN_3467; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_337 = memReg_46_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_338 = |_T_337; // @[fifo.scala 109:63]
  wire [4:0] _memReg_46_branch_mask_T = memReg_46_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3762 = |_T_337 ? _memReg_46_branch_mask_T : _GEN_3404; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3763 = _T_338 ? 1'h0 : _GEN_3468; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_344 = memReg_47_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_345 = |_T_344; // @[fifo.scala 109:63]
  wire [4:0] _memReg_47_branch_mask_T = memReg_47_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3768 = |_T_344 ? _memReg_47_branch_mask_T : _GEN_3405; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3769 = _T_345 ? 1'h0 : _GEN_3469; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_351 = memReg_48_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_352 = |_T_351; // @[fifo.scala 109:63]
  wire [4:0] _memReg_48_branch_mask_T = memReg_48_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3774 = |_T_351 ? _memReg_48_branch_mask_T : _GEN_3406; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3775 = _T_352 ? 1'h0 : _GEN_3470; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_358 = memReg_49_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_359 = |_T_358; // @[fifo.scala 109:63]
  wire [4:0] _memReg_49_branch_mask_T = memReg_49_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3780 = |_T_358 ? _memReg_49_branch_mask_T : _GEN_3407; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3781 = _T_359 ? 1'h0 : _GEN_3471; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_365 = memReg_50_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_366 = |_T_365; // @[fifo.scala 109:63]
  wire [4:0] _memReg_50_branch_mask_T = memReg_50_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3786 = |_T_365 ? _memReg_50_branch_mask_T : _GEN_3408; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3787 = _T_366 ? 1'h0 : _GEN_3472; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_372 = memReg_51_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_373 = |_T_372; // @[fifo.scala 109:63]
  wire [4:0] _memReg_51_branch_mask_T = memReg_51_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3792 = |_T_372 ? _memReg_51_branch_mask_T : _GEN_3409; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3793 = _T_373 ? 1'h0 : _GEN_3473; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_379 = memReg_52_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_380 = |_T_379; // @[fifo.scala 109:63]
  wire [4:0] _memReg_52_branch_mask_T = memReg_52_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3798 = |_T_379 ? _memReg_52_branch_mask_T : _GEN_3410; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3799 = _T_380 ? 1'h0 : _GEN_3474; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_386 = memReg_53_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_387 = |_T_386; // @[fifo.scala 109:63]
  wire [4:0] _memReg_53_branch_mask_T = memReg_53_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3804 = |_T_386 ? _memReg_53_branch_mask_T : _GEN_3411; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3805 = _T_387 ? 1'h0 : _GEN_3475; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_393 = memReg_54_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_394 = |_T_393; // @[fifo.scala 109:63]
  wire [4:0] _memReg_54_branch_mask_T = memReg_54_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3810 = |_T_393 ? _memReg_54_branch_mask_T : _GEN_3412; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3811 = _T_394 ? 1'h0 : _GEN_3476; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_400 = memReg_55_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_401 = |_T_400; // @[fifo.scala 109:63]
  wire [4:0] _memReg_55_branch_mask_T = memReg_55_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3816 = |_T_400 ? _memReg_55_branch_mask_T : _GEN_3413; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3817 = _T_401 ? 1'h0 : _GEN_3477; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_407 = memReg_56_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_408 = |_T_407; // @[fifo.scala 109:63]
  wire [4:0] _memReg_56_branch_mask_T = memReg_56_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3822 = |_T_407 ? _memReg_56_branch_mask_T : _GEN_3414; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3823 = _T_408 ? 1'h0 : _GEN_3478; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_414 = memReg_57_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_415 = |_T_414; // @[fifo.scala 109:63]
  wire [4:0] _memReg_57_branch_mask_T = memReg_57_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3828 = |_T_414 ? _memReg_57_branch_mask_T : _GEN_3415; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3829 = _T_415 ? 1'h0 : _GEN_3479; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_421 = memReg_58_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_422 = |_T_421; // @[fifo.scala 109:63]
  wire [4:0] _memReg_58_branch_mask_T = memReg_58_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3834 = |_T_421 ? _memReg_58_branch_mask_T : _GEN_3416; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3835 = _T_422 ? 1'h0 : _GEN_3480; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_428 = memReg_59_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_429 = |_T_428; // @[fifo.scala 109:63]
  wire [4:0] _memReg_59_branch_mask_T = memReg_59_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3840 = |_T_428 ? _memReg_59_branch_mask_T : _GEN_3417; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3841 = _T_429 ? 1'h0 : _GEN_3481; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_435 = memReg_60_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_436 = |_T_435; // @[fifo.scala 109:63]
  wire [4:0] _memReg_60_branch_mask_T = memReg_60_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3846 = |_T_435 ? _memReg_60_branch_mask_T : _GEN_3418; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3847 = _T_436 ? 1'h0 : _GEN_3482; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_442 = memReg_61_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_443 = |_T_442; // @[fifo.scala 109:63]
  wire [4:0] _memReg_61_branch_mask_T = memReg_61_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3852 = |_T_442 ? _memReg_61_branch_mask_T : _GEN_3419; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3853 = _T_443 ? 1'h0 : _GEN_3483; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_449 = memReg_62_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_450 = |_T_449; // @[fifo.scala 109:63]
  wire [4:0] _memReg_62_branch_mask_T = memReg_62_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _GEN_3858 = |_T_449 ? _memReg_62_branch_mask_T : _GEN_3420; // @[fifo.scala 109:68 110:35]
  wire  _GEN_3859 = _T_450 ? 1'h0 : _GEN_3484; // @[fifo.scala 113:68 114:36]
  wire [4:0] _T_456 = memReg_63_branch_mask & branchOps_branchMask; // @[fifo.scala 109:39]
  wire  _T_457 = |_T_456; // @[fifo.scala 109:63]
  wire [4:0] _memReg_63_branch_mask_T = memReg_63_branch_mask ^ branchOps_branchMask; // @[fifo.scala 110:60]
  wire [4:0] _T_462 = _GEN_2013 & branchOps_branchMask; // @[utils.scala 101:27]
  wire  _GEN_4000 = |_T_462 ? 1'h0 : _GEN_1949; // @[utils.scala 101:56 103:28 107:28]
  wire  _GEN_4002 = branchOps_passed ? _GEN_1949 : _GEN_4000; // @[utils.scala 90:30 98:26]
  assign read_data_valid = _T_2 & _GEN_1629; // @[fifo.scala 122:32]
  assign read_data_branch_valid = branchOps_valid ? _GEN_4002 : _GEN_1949; // @[utils.scala 112:24 89:27]
  assign isEmpty = emptyReg; // @[fifo.scala 89:11]
  assign isFull = fullReg; // @[fifo.scala 148:10]
  always @(posedge clock) begin
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_0_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_0_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_0_valid <= _GEN_798;
      end
    end else begin
      memReg_0_valid <= _GEN_798;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h0 == writePtr) begin // @[fifo.scala 82:22]
        memReg_0_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (branchOps_passed) begin // @[fifo.scala 108:32]
        memReg_0_branch_valid <= _GEN_3422;
      end else if (_T_16) begin // @[fifo.scala 113:68]
        memReg_0_branch_valid <= 1'h0; // @[fifo.scala 114:36]
      end else begin
        memReg_0_branch_valid <= _GEN_3422;
      end
    end else begin
      memReg_0_branch_valid <= _GEN_3422;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_0_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (branchOps_passed) begin // @[fifo.scala 108:32]
        if (|_T_15) begin // @[fifo.scala 109:68]
          memReg_0_branch_mask <= _memReg_0_branch_mask_T; // @[fifo.scala 110:35]
        end else begin
          memReg_0_branch_mask <= _GEN_3358;
        end
      end else begin
        memReg_0_branch_mask <= _GEN_3358;
      end
    end else begin
      memReg_0_branch_mask <= _GEN_3358;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_1_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_1_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_1_valid <= _GEN_799;
      end
    end else begin
      memReg_1_valid <= _GEN_799;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h1 == writePtr) begin // @[fifo.scala 82:22]
        memReg_1_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h1 | 6'h1 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_1_branch_valid <= _GEN_3423;
        end else begin
          memReg_1_branch_valid <= _GEN_3493;
        end
      end else begin
        memReg_1_branch_valid <= _GEN_3423;
      end
    end else begin
      memReg_1_branch_valid <= _GEN_3423;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_1_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h1 | 6'h1 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_1_branch_mask <= _GEN_3492;
        end else begin
          memReg_1_branch_mask <= _GEN_3359;
        end
      end else begin
        memReg_1_branch_mask <= _GEN_3359;
      end
    end else begin
      memReg_1_branch_mask <= _GEN_3359;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_2_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_2_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_2_valid <= _GEN_800;
      end
    end else begin
      memReg_2_valid <= _GEN_800;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h2 == writePtr) begin // @[fifo.scala 82:22]
        memReg_2_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h2 | 6'h2 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_2_branch_valid <= _GEN_3424;
        end else begin
          memReg_2_branch_valid <= _GEN_3499;
        end
      end else begin
        memReg_2_branch_valid <= _GEN_3424;
      end
    end else begin
      memReg_2_branch_valid <= _GEN_3424;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_2_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h2 | 6'h2 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_2_branch_mask <= _GEN_3498;
        end else begin
          memReg_2_branch_mask <= _GEN_3360;
        end
      end else begin
        memReg_2_branch_mask <= _GEN_3360;
      end
    end else begin
      memReg_2_branch_mask <= _GEN_3360;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_3_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_3_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_3_valid <= _GEN_801;
      end
    end else begin
      memReg_3_valid <= _GEN_801;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h3 == writePtr) begin // @[fifo.scala 82:22]
        memReg_3_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h3 | 6'h3 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_3_branch_valid <= _GEN_3425;
        end else begin
          memReg_3_branch_valid <= _GEN_3505;
        end
      end else begin
        memReg_3_branch_valid <= _GEN_3425;
      end
    end else begin
      memReg_3_branch_valid <= _GEN_3425;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_3_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h3 | 6'h3 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_3_branch_mask <= _GEN_3504;
        end else begin
          memReg_3_branch_mask <= _GEN_3361;
        end
      end else begin
        memReg_3_branch_mask <= _GEN_3361;
      end
    end else begin
      memReg_3_branch_mask <= _GEN_3361;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_4_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_4_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_4_valid <= _GEN_802;
      end
    end else begin
      memReg_4_valid <= _GEN_802;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h4 == writePtr) begin // @[fifo.scala 82:22]
        memReg_4_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h4 | 6'h4 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_4_branch_valid <= _GEN_3426;
        end else begin
          memReg_4_branch_valid <= _GEN_3511;
        end
      end else begin
        memReg_4_branch_valid <= _GEN_3426;
      end
    end else begin
      memReg_4_branch_valid <= _GEN_3426;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_4_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h4 | 6'h4 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_4_branch_mask <= _GEN_3510;
        end else begin
          memReg_4_branch_mask <= _GEN_3362;
        end
      end else begin
        memReg_4_branch_mask <= _GEN_3362;
      end
    end else begin
      memReg_4_branch_mask <= _GEN_3362;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_5_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_5_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_5_valid <= _GEN_803;
      end
    end else begin
      memReg_5_valid <= _GEN_803;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h5 == writePtr) begin // @[fifo.scala 82:22]
        memReg_5_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h5 | 6'h5 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_5_branch_valid <= _GEN_3427;
        end else begin
          memReg_5_branch_valid <= _GEN_3517;
        end
      end else begin
        memReg_5_branch_valid <= _GEN_3427;
      end
    end else begin
      memReg_5_branch_valid <= _GEN_3427;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_5_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h5 | 6'h5 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_5_branch_mask <= _GEN_3516;
        end else begin
          memReg_5_branch_mask <= _GEN_3363;
        end
      end else begin
        memReg_5_branch_mask <= _GEN_3363;
      end
    end else begin
      memReg_5_branch_mask <= _GEN_3363;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_6_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_6_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_6_valid <= _GEN_804;
      end
    end else begin
      memReg_6_valid <= _GEN_804;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h6 == writePtr) begin // @[fifo.scala 82:22]
        memReg_6_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h6 | 6'h6 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_6_branch_valid <= _GEN_3428;
        end else begin
          memReg_6_branch_valid <= _GEN_3523;
        end
      end else begin
        memReg_6_branch_valid <= _GEN_3428;
      end
    end else begin
      memReg_6_branch_valid <= _GEN_3428;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_6_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h6 | 6'h6 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_6_branch_mask <= _GEN_3522;
        end else begin
          memReg_6_branch_mask <= _GEN_3364;
        end
      end else begin
        memReg_6_branch_mask <= _GEN_3364;
      end
    end else begin
      memReg_6_branch_mask <= _GEN_3364;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_7_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_7_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_7_valid <= _GEN_805;
      end
    end else begin
      memReg_7_valid <= _GEN_805;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h7 == writePtr) begin // @[fifo.scala 82:22]
        memReg_7_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h7 | 6'h7 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_7_branch_valid <= _GEN_3429;
        end else begin
          memReg_7_branch_valid <= _GEN_3529;
        end
      end else begin
        memReg_7_branch_valid <= _GEN_3429;
      end
    end else begin
      memReg_7_branch_valid <= _GEN_3429;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_7_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h7 | 6'h7 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_7_branch_mask <= _GEN_3528;
        end else begin
          memReg_7_branch_mask <= _GEN_3365;
        end
      end else begin
        memReg_7_branch_mask <= _GEN_3365;
      end
    end else begin
      memReg_7_branch_mask <= _GEN_3365;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_8_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_8_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_8_valid <= _GEN_806;
      end
    end else begin
      memReg_8_valid <= _GEN_806;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h8 == writePtr) begin // @[fifo.scala 82:22]
        memReg_8_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h8 | 6'h8 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_8_branch_valid <= _GEN_3430;
        end else begin
          memReg_8_branch_valid <= _GEN_3535;
        end
      end else begin
        memReg_8_branch_valid <= _GEN_3430;
      end
    end else begin
      memReg_8_branch_valid <= _GEN_3430;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_8_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h8 | 6'h8 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_8_branch_mask <= _GEN_3534;
        end else begin
          memReg_8_branch_mask <= _GEN_3366;
        end
      end else begin
        memReg_8_branch_mask <= _GEN_3366;
      end
    end else begin
      memReg_8_branch_mask <= _GEN_3366;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_9_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_9_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_9_valid <= _GEN_807;
      end
    end else begin
      memReg_9_valid <= _GEN_807;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h9 == writePtr) begin // @[fifo.scala 82:22]
        memReg_9_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h9 | 6'h9 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_9_branch_valid <= _GEN_3431;
        end else begin
          memReg_9_branch_valid <= _GEN_3541;
        end
      end else begin
        memReg_9_branch_valid <= _GEN_3431;
      end
    end else begin
      memReg_9_branch_valid <= _GEN_3431;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_9_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h9 | 6'h9 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_9_branch_mask <= _GEN_3540;
        end else begin
          memReg_9_branch_mask <= _GEN_3367;
        end
      end else begin
        memReg_9_branch_mask <= _GEN_3367;
      end
    end else begin
      memReg_9_branch_mask <= _GEN_3367;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_10_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_10_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_10_valid <= _GEN_808;
      end
    end else begin
      memReg_10_valid <= _GEN_808;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'ha == writePtr) begin // @[fifo.scala 82:22]
        memReg_10_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'ha | 6'ha <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_10_branch_valid <= _GEN_3432;
        end else begin
          memReg_10_branch_valid <= _GEN_3547;
        end
      end else begin
        memReg_10_branch_valid <= _GEN_3432;
      end
    end else begin
      memReg_10_branch_valid <= _GEN_3432;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_10_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'ha | 6'ha <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_10_branch_mask <= _GEN_3546;
        end else begin
          memReg_10_branch_mask <= _GEN_3368;
        end
      end else begin
        memReg_10_branch_mask <= _GEN_3368;
      end
    end else begin
      memReg_10_branch_mask <= _GEN_3368;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_11_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_11_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_11_valid <= _GEN_809;
      end
    end else begin
      memReg_11_valid <= _GEN_809;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'hb == writePtr) begin // @[fifo.scala 82:22]
        memReg_11_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'hb | 6'hb <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_11_branch_valid <= _GEN_3433;
        end else begin
          memReg_11_branch_valid <= _GEN_3553;
        end
      end else begin
        memReg_11_branch_valid <= _GEN_3433;
      end
    end else begin
      memReg_11_branch_valid <= _GEN_3433;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_11_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'hb | 6'hb <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_11_branch_mask <= _GEN_3552;
        end else begin
          memReg_11_branch_mask <= _GEN_3369;
        end
      end else begin
        memReg_11_branch_mask <= _GEN_3369;
      end
    end else begin
      memReg_11_branch_mask <= _GEN_3369;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_12_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_12_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_12_valid <= _GEN_810;
      end
    end else begin
      memReg_12_valid <= _GEN_810;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'hc == writePtr) begin // @[fifo.scala 82:22]
        memReg_12_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'hc | 6'hc <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_12_branch_valid <= _GEN_3434;
        end else begin
          memReg_12_branch_valid <= _GEN_3559;
        end
      end else begin
        memReg_12_branch_valid <= _GEN_3434;
      end
    end else begin
      memReg_12_branch_valid <= _GEN_3434;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_12_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'hc | 6'hc <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_12_branch_mask <= _GEN_3558;
        end else begin
          memReg_12_branch_mask <= _GEN_3370;
        end
      end else begin
        memReg_12_branch_mask <= _GEN_3370;
      end
    end else begin
      memReg_12_branch_mask <= _GEN_3370;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_13_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_13_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_13_valid <= _GEN_811;
      end
    end else begin
      memReg_13_valid <= _GEN_811;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'hd == writePtr) begin // @[fifo.scala 82:22]
        memReg_13_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'hd | 6'hd <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_13_branch_valid <= _GEN_3435;
        end else begin
          memReg_13_branch_valid <= _GEN_3565;
        end
      end else begin
        memReg_13_branch_valid <= _GEN_3435;
      end
    end else begin
      memReg_13_branch_valid <= _GEN_3435;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_13_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'hd | 6'hd <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_13_branch_mask <= _GEN_3564;
        end else begin
          memReg_13_branch_mask <= _GEN_3371;
        end
      end else begin
        memReg_13_branch_mask <= _GEN_3371;
      end
    end else begin
      memReg_13_branch_mask <= _GEN_3371;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_14_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_14_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_14_valid <= _GEN_812;
      end
    end else begin
      memReg_14_valid <= _GEN_812;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'he == writePtr) begin // @[fifo.scala 82:22]
        memReg_14_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'he | 6'he <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_14_branch_valid <= _GEN_3436;
        end else begin
          memReg_14_branch_valid <= _GEN_3571;
        end
      end else begin
        memReg_14_branch_valid <= _GEN_3436;
      end
    end else begin
      memReg_14_branch_valid <= _GEN_3436;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_14_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'he | 6'he <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_14_branch_mask <= _GEN_3570;
        end else begin
          memReg_14_branch_mask <= _GEN_3372;
        end
      end else begin
        memReg_14_branch_mask <= _GEN_3372;
      end
    end else begin
      memReg_14_branch_mask <= _GEN_3372;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_15_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_15_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_15_valid <= _GEN_813;
      end
    end else begin
      memReg_15_valid <= _GEN_813;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'hf == writePtr) begin // @[fifo.scala 82:22]
        memReg_15_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'hf | 6'hf <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_15_branch_valid <= _GEN_3437;
        end else begin
          memReg_15_branch_valid <= _GEN_3577;
        end
      end else begin
        memReg_15_branch_valid <= _GEN_3437;
      end
    end else begin
      memReg_15_branch_valid <= _GEN_3437;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_15_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'hf | 6'hf <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_15_branch_mask <= _GEN_3576;
        end else begin
          memReg_15_branch_mask <= _GEN_3373;
        end
      end else begin
        memReg_15_branch_mask <= _GEN_3373;
      end
    end else begin
      memReg_15_branch_mask <= _GEN_3373;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_16_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_16_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_16_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_16_valid <= _GEN_814;
      end
    end else begin
      memReg_16_valid <= _GEN_814;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_16_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h10 == writePtr) begin // @[fifo.scala 82:22]
        memReg_16_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_16_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h10 | 6'h10 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_16_branch_valid <= _GEN_3438;
        end else begin
          memReg_16_branch_valid <= _GEN_3583;
        end
      end else begin
        memReg_16_branch_valid <= _GEN_3438;
      end
    end else begin
      memReg_16_branch_valid <= _GEN_3438;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_16_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h10 | 6'h10 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_16_branch_mask <= _GEN_3582;
        end else begin
          memReg_16_branch_mask <= _GEN_3374;
        end
      end else begin
        memReg_16_branch_mask <= _GEN_3374;
      end
    end else begin
      memReg_16_branch_mask <= _GEN_3374;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_17_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_17_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_17_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_17_valid <= _GEN_815;
      end
    end else begin
      memReg_17_valid <= _GEN_815;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_17_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h11 == writePtr) begin // @[fifo.scala 82:22]
        memReg_17_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_17_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h11 | 6'h11 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_17_branch_valid <= _GEN_3439;
        end else begin
          memReg_17_branch_valid <= _GEN_3589;
        end
      end else begin
        memReg_17_branch_valid <= _GEN_3439;
      end
    end else begin
      memReg_17_branch_valid <= _GEN_3439;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_17_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h11 | 6'h11 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_17_branch_mask <= _GEN_3588;
        end else begin
          memReg_17_branch_mask <= _GEN_3375;
        end
      end else begin
        memReg_17_branch_mask <= _GEN_3375;
      end
    end else begin
      memReg_17_branch_mask <= _GEN_3375;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_18_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_18_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_18_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_18_valid <= _GEN_816;
      end
    end else begin
      memReg_18_valid <= _GEN_816;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_18_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h12 == writePtr) begin // @[fifo.scala 82:22]
        memReg_18_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_18_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h12 | 6'h12 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_18_branch_valid <= _GEN_3440;
        end else begin
          memReg_18_branch_valid <= _GEN_3595;
        end
      end else begin
        memReg_18_branch_valid <= _GEN_3440;
      end
    end else begin
      memReg_18_branch_valid <= _GEN_3440;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_18_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h12 | 6'h12 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_18_branch_mask <= _GEN_3594;
        end else begin
          memReg_18_branch_mask <= _GEN_3376;
        end
      end else begin
        memReg_18_branch_mask <= _GEN_3376;
      end
    end else begin
      memReg_18_branch_mask <= _GEN_3376;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_19_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_19_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_19_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_19_valid <= _GEN_817;
      end
    end else begin
      memReg_19_valid <= _GEN_817;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_19_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h13 == writePtr) begin // @[fifo.scala 82:22]
        memReg_19_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_19_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h13 | 6'h13 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_19_branch_valid <= _GEN_3441;
        end else begin
          memReg_19_branch_valid <= _GEN_3601;
        end
      end else begin
        memReg_19_branch_valid <= _GEN_3441;
      end
    end else begin
      memReg_19_branch_valid <= _GEN_3441;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_19_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h13 | 6'h13 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_19_branch_mask <= _GEN_3600;
        end else begin
          memReg_19_branch_mask <= _GEN_3377;
        end
      end else begin
        memReg_19_branch_mask <= _GEN_3377;
      end
    end else begin
      memReg_19_branch_mask <= _GEN_3377;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_20_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_20_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_20_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_20_valid <= _GEN_818;
      end
    end else begin
      memReg_20_valid <= _GEN_818;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_20_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h14 == writePtr) begin // @[fifo.scala 82:22]
        memReg_20_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_20_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h14 | 6'h14 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_20_branch_valid <= _GEN_3442;
        end else begin
          memReg_20_branch_valid <= _GEN_3607;
        end
      end else begin
        memReg_20_branch_valid <= _GEN_3442;
      end
    end else begin
      memReg_20_branch_valid <= _GEN_3442;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_20_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h14 | 6'h14 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_20_branch_mask <= _GEN_3606;
        end else begin
          memReg_20_branch_mask <= _GEN_3378;
        end
      end else begin
        memReg_20_branch_mask <= _GEN_3378;
      end
    end else begin
      memReg_20_branch_mask <= _GEN_3378;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_21_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_21_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_21_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_21_valid <= _GEN_819;
      end
    end else begin
      memReg_21_valid <= _GEN_819;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_21_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h15 == writePtr) begin // @[fifo.scala 82:22]
        memReg_21_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_21_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h15 | 6'h15 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_21_branch_valid <= _GEN_3443;
        end else begin
          memReg_21_branch_valid <= _GEN_3613;
        end
      end else begin
        memReg_21_branch_valid <= _GEN_3443;
      end
    end else begin
      memReg_21_branch_valid <= _GEN_3443;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_21_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h15 | 6'h15 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_21_branch_mask <= _GEN_3612;
        end else begin
          memReg_21_branch_mask <= _GEN_3379;
        end
      end else begin
        memReg_21_branch_mask <= _GEN_3379;
      end
    end else begin
      memReg_21_branch_mask <= _GEN_3379;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_22_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_22_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_22_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_22_valid <= _GEN_820;
      end
    end else begin
      memReg_22_valid <= _GEN_820;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_22_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h16 == writePtr) begin // @[fifo.scala 82:22]
        memReg_22_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_22_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h16 | 6'h16 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_22_branch_valid <= _GEN_3444;
        end else begin
          memReg_22_branch_valid <= _GEN_3619;
        end
      end else begin
        memReg_22_branch_valid <= _GEN_3444;
      end
    end else begin
      memReg_22_branch_valid <= _GEN_3444;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_22_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h16 | 6'h16 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_22_branch_mask <= _GEN_3618;
        end else begin
          memReg_22_branch_mask <= _GEN_3380;
        end
      end else begin
        memReg_22_branch_mask <= _GEN_3380;
      end
    end else begin
      memReg_22_branch_mask <= _GEN_3380;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_23_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_23_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_23_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_23_valid <= _GEN_821;
      end
    end else begin
      memReg_23_valid <= _GEN_821;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_23_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h17 == writePtr) begin // @[fifo.scala 82:22]
        memReg_23_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_23_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h17 | 6'h17 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_23_branch_valid <= _GEN_3445;
        end else begin
          memReg_23_branch_valid <= _GEN_3625;
        end
      end else begin
        memReg_23_branch_valid <= _GEN_3445;
      end
    end else begin
      memReg_23_branch_valid <= _GEN_3445;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_23_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h17 | 6'h17 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_23_branch_mask <= _GEN_3624;
        end else begin
          memReg_23_branch_mask <= _GEN_3381;
        end
      end else begin
        memReg_23_branch_mask <= _GEN_3381;
      end
    end else begin
      memReg_23_branch_mask <= _GEN_3381;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_24_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_24_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_24_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_24_valid <= _GEN_822;
      end
    end else begin
      memReg_24_valid <= _GEN_822;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_24_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h18 == writePtr) begin // @[fifo.scala 82:22]
        memReg_24_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_24_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h18 | 6'h18 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_24_branch_valid <= _GEN_3446;
        end else begin
          memReg_24_branch_valid <= _GEN_3631;
        end
      end else begin
        memReg_24_branch_valid <= _GEN_3446;
      end
    end else begin
      memReg_24_branch_valid <= _GEN_3446;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_24_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h18 | 6'h18 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_24_branch_mask <= _GEN_3630;
        end else begin
          memReg_24_branch_mask <= _GEN_3382;
        end
      end else begin
        memReg_24_branch_mask <= _GEN_3382;
      end
    end else begin
      memReg_24_branch_mask <= _GEN_3382;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_25_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_25_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_25_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_25_valid <= _GEN_823;
      end
    end else begin
      memReg_25_valid <= _GEN_823;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_25_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h19 == writePtr) begin // @[fifo.scala 82:22]
        memReg_25_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_25_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h19 | 6'h19 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_25_branch_valid <= _GEN_3447;
        end else begin
          memReg_25_branch_valid <= _GEN_3637;
        end
      end else begin
        memReg_25_branch_valid <= _GEN_3447;
      end
    end else begin
      memReg_25_branch_valid <= _GEN_3447;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_25_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h19 | 6'h19 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_25_branch_mask <= _GEN_3636;
        end else begin
          memReg_25_branch_mask <= _GEN_3383;
        end
      end else begin
        memReg_25_branch_mask <= _GEN_3383;
      end
    end else begin
      memReg_25_branch_mask <= _GEN_3383;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_26_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_26_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_26_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_26_valid <= _GEN_824;
      end
    end else begin
      memReg_26_valid <= _GEN_824;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_26_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h1a == writePtr) begin // @[fifo.scala 82:22]
        memReg_26_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_26_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h1a | 6'h1a <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_26_branch_valid <= _GEN_3448;
        end else begin
          memReg_26_branch_valid <= _GEN_3643;
        end
      end else begin
        memReg_26_branch_valid <= _GEN_3448;
      end
    end else begin
      memReg_26_branch_valid <= _GEN_3448;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_26_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h1a | 6'h1a <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_26_branch_mask <= _GEN_3642;
        end else begin
          memReg_26_branch_mask <= _GEN_3384;
        end
      end else begin
        memReg_26_branch_mask <= _GEN_3384;
      end
    end else begin
      memReg_26_branch_mask <= _GEN_3384;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_27_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_27_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_27_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_27_valid <= _GEN_825;
      end
    end else begin
      memReg_27_valid <= _GEN_825;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_27_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h1b == writePtr) begin // @[fifo.scala 82:22]
        memReg_27_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_27_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h1b | 6'h1b <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_27_branch_valid <= _GEN_3449;
        end else begin
          memReg_27_branch_valid <= _GEN_3649;
        end
      end else begin
        memReg_27_branch_valid <= _GEN_3449;
      end
    end else begin
      memReg_27_branch_valid <= _GEN_3449;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_27_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h1b | 6'h1b <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_27_branch_mask <= _GEN_3648;
        end else begin
          memReg_27_branch_mask <= _GEN_3385;
        end
      end else begin
        memReg_27_branch_mask <= _GEN_3385;
      end
    end else begin
      memReg_27_branch_mask <= _GEN_3385;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_28_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_28_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_28_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_28_valid <= _GEN_826;
      end
    end else begin
      memReg_28_valid <= _GEN_826;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_28_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h1c == writePtr) begin // @[fifo.scala 82:22]
        memReg_28_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_28_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h1c | 6'h1c <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_28_branch_valid <= _GEN_3450;
        end else begin
          memReg_28_branch_valid <= _GEN_3655;
        end
      end else begin
        memReg_28_branch_valid <= _GEN_3450;
      end
    end else begin
      memReg_28_branch_valid <= _GEN_3450;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_28_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h1c | 6'h1c <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_28_branch_mask <= _GEN_3654;
        end else begin
          memReg_28_branch_mask <= _GEN_3386;
        end
      end else begin
        memReg_28_branch_mask <= _GEN_3386;
      end
    end else begin
      memReg_28_branch_mask <= _GEN_3386;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_29_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_29_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_29_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_29_valid <= _GEN_827;
      end
    end else begin
      memReg_29_valid <= _GEN_827;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_29_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h1d == writePtr) begin // @[fifo.scala 82:22]
        memReg_29_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_29_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h1d | 6'h1d <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_29_branch_valid <= _GEN_3451;
        end else begin
          memReg_29_branch_valid <= _GEN_3661;
        end
      end else begin
        memReg_29_branch_valid <= _GEN_3451;
      end
    end else begin
      memReg_29_branch_valid <= _GEN_3451;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_29_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h1d | 6'h1d <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_29_branch_mask <= _GEN_3660;
        end else begin
          memReg_29_branch_mask <= _GEN_3387;
        end
      end else begin
        memReg_29_branch_mask <= _GEN_3387;
      end
    end else begin
      memReg_29_branch_mask <= _GEN_3387;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_30_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_30_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_30_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_30_valid <= _GEN_828;
      end
    end else begin
      memReg_30_valid <= _GEN_828;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_30_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h1e == writePtr) begin // @[fifo.scala 82:22]
        memReg_30_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_30_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h1e | 6'h1e <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_30_branch_valid <= _GEN_3452;
        end else begin
          memReg_30_branch_valid <= _GEN_3667;
        end
      end else begin
        memReg_30_branch_valid <= _GEN_3452;
      end
    end else begin
      memReg_30_branch_valid <= _GEN_3452;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_30_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h1e | 6'h1e <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_30_branch_mask <= _GEN_3666;
        end else begin
          memReg_30_branch_mask <= _GEN_3388;
        end
      end else begin
        memReg_30_branch_mask <= _GEN_3388;
      end
    end else begin
      memReg_30_branch_mask <= _GEN_3388;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_31_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_31_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_31_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_31_valid <= _GEN_829;
      end
    end else begin
      memReg_31_valid <= _GEN_829;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_31_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h1f == writePtr) begin // @[fifo.scala 82:22]
        memReg_31_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_31_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h1f | 6'h1f <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_31_branch_valid <= _GEN_3453;
        end else begin
          memReg_31_branch_valid <= _GEN_3673;
        end
      end else begin
        memReg_31_branch_valid <= _GEN_3453;
      end
    end else begin
      memReg_31_branch_valid <= _GEN_3453;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_31_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h1f | 6'h1f <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_31_branch_mask <= _GEN_3672;
        end else begin
          memReg_31_branch_mask <= _GEN_3389;
        end
      end else begin
        memReg_31_branch_mask <= _GEN_3389;
      end
    end else begin
      memReg_31_branch_mask <= _GEN_3389;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_32_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_32_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_32_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_32_valid <= _GEN_830;
      end
    end else begin
      memReg_32_valid <= _GEN_830;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_32_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h20 == writePtr) begin // @[fifo.scala 82:22]
        memReg_32_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_32_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h20 | 6'h20 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_32_branch_valid <= _GEN_3454;
        end else begin
          memReg_32_branch_valid <= _GEN_3679;
        end
      end else begin
        memReg_32_branch_valid <= _GEN_3454;
      end
    end else begin
      memReg_32_branch_valid <= _GEN_3454;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_32_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h20 | 6'h20 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_32_branch_mask <= _GEN_3678;
        end else begin
          memReg_32_branch_mask <= _GEN_3390;
        end
      end else begin
        memReg_32_branch_mask <= _GEN_3390;
      end
    end else begin
      memReg_32_branch_mask <= _GEN_3390;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_33_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_33_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_33_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_33_valid <= _GEN_831;
      end
    end else begin
      memReg_33_valid <= _GEN_831;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_33_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h21 == writePtr) begin // @[fifo.scala 82:22]
        memReg_33_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_33_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h21 | 6'h21 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_33_branch_valid <= _GEN_3455;
        end else begin
          memReg_33_branch_valid <= _GEN_3685;
        end
      end else begin
        memReg_33_branch_valid <= _GEN_3455;
      end
    end else begin
      memReg_33_branch_valid <= _GEN_3455;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_33_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h21 | 6'h21 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_33_branch_mask <= _GEN_3684;
        end else begin
          memReg_33_branch_mask <= _GEN_3391;
        end
      end else begin
        memReg_33_branch_mask <= _GEN_3391;
      end
    end else begin
      memReg_33_branch_mask <= _GEN_3391;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_34_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_34_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_34_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_34_valid <= _GEN_832;
      end
    end else begin
      memReg_34_valid <= _GEN_832;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_34_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h22 == writePtr) begin // @[fifo.scala 82:22]
        memReg_34_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_34_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h22 | 6'h22 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_34_branch_valid <= _GEN_3456;
        end else begin
          memReg_34_branch_valid <= _GEN_3691;
        end
      end else begin
        memReg_34_branch_valid <= _GEN_3456;
      end
    end else begin
      memReg_34_branch_valid <= _GEN_3456;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_34_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h22 | 6'h22 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_34_branch_mask <= _GEN_3690;
        end else begin
          memReg_34_branch_mask <= _GEN_3392;
        end
      end else begin
        memReg_34_branch_mask <= _GEN_3392;
      end
    end else begin
      memReg_34_branch_mask <= _GEN_3392;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_35_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_35_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_35_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_35_valid <= _GEN_833;
      end
    end else begin
      memReg_35_valid <= _GEN_833;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_35_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h23 == writePtr) begin // @[fifo.scala 82:22]
        memReg_35_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_35_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h23 | 6'h23 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_35_branch_valid <= _GEN_3457;
        end else begin
          memReg_35_branch_valid <= _GEN_3697;
        end
      end else begin
        memReg_35_branch_valid <= _GEN_3457;
      end
    end else begin
      memReg_35_branch_valid <= _GEN_3457;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_35_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h23 | 6'h23 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_35_branch_mask <= _GEN_3696;
        end else begin
          memReg_35_branch_mask <= _GEN_3393;
        end
      end else begin
        memReg_35_branch_mask <= _GEN_3393;
      end
    end else begin
      memReg_35_branch_mask <= _GEN_3393;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_36_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_36_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_36_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_36_valid <= _GEN_834;
      end
    end else begin
      memReg_36_valid <= _GEN_834;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_36_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h24 == writePtr) begin // @[fifo.scala 82:22]
        memReg_36_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_36_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h24 | 6'h24 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_36_branch_valid <= _GEN_3458;
        end else begin
          memReg_36_branch_valid <= _GEN_3703;
        end
      end else begin
        memReg_36_branch_valid <= _GEN_3458;
      end
    end else begin
      memReg_36_branch_valid <= _GEN_3458;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_36_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h24 | 6'h24 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_36_branch_mask <= _GEN_3702;
        end else begin
          memReg_36_branch_mask <= _GEN_3394;
        end
      end else begin
        memReg_36_branch_mask <= _GEN_3394;
      end
    end else begin
      memReg_36_branch_mask <= _GEN_3394;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_37_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_37_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_37_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_37_valid <= _GEN_835;
      end
    end else begin
      memReg_37_valid <= _GEN_835;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_37_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h25 == writePtr) begin // @[fifo.scala 82:22]
        memReg_37_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_37_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h25 | 6'h25 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_37_branch_valid <= _GEN_3459;
        end else begin
          memReg_37_branch_valid <= _GEN_3709;
        end
      end else begin
        memReg_37_branch_valid <= _GEN_3459;
      end
    end else begin
      memReg_37_branch_valid <= _GEN_3459;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_37_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h25 | 6'h25 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_37_branch_mask <= _GEN_3708;
        end else begin
          memReg_37_branch_mask <= _GEN_3395;
        end
      end else begin
        memReg_37_branch_mask <= _GEN_3395;
      end
    end else begin
      memReg_37_branch_mask <= _GEN_3395;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_38_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_38_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_38_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_38_valid <= _GEN_836;
      end
    end else begin
      memReg_38_valid <= _GEN_836;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_38_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h26 == writePtr) begin // @[fifo.scala 82:22]
        memReg_38_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_38_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h26 | 6'h26 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_38_branch_valid <= _GEN_3460;
        end else begin
          memReg_38_branch_valid <= _GEN_3715;
        end
      end else begin
        memReg_38_branch_valid <= _GEN_3460;
      end
    end else begin
      memReg_38_branch_valid <= _GEN_3460;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_38_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h26 | 6'h26 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_38_branch_mask <= _GEN_3714;
        end else begin
          memReg_38_branch_mask <= _GEN_3396;
        end
      end else begin
        memReg_38_branch_mask <= _GEN_3396;
      end
    end else begin
      memReg_38_branch_mask <= _GEN_3396;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_39_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_39_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_39_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_39_valid <= _GEN_837;
      end
    end else begin
      memReg_39_valid <= _GEN_837;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_39_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h27 == writePtr) begin // @[fifo.scala 82:22]
        memReg_39_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_39_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h27 | 6'h27 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_39_branch_valid <= _GEN_3461;
        end else begin
          memReg_39_branch_valid <= _GEN_3721;
        end
      end else begin
        memReg_39_branch_valid <= _GEN_3461;
      end
    end else begin
      memReg_39_branch_valid <= _GEN_3461;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_39_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h27 | 6'h27 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_39_branch_mask <= _GEN_3720;
        end else begin
          memReg_39_branch_mask <= _GEN_3397;
        end
      end else begin
        memReg_39_branch_mask <= _GEN_3397;
      end
    end else begin
      memReg_39_branch_mask <= _GEN_3397;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_40_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_40_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_40_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_40_valid <= _GEN_838;
      end
    end else begin
      memReg_40_valid <= _GEN_838;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_40_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h28 == writePtr) begin // @[fifo.scala 82:22]
        memReg_40_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_40_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h28 | 6'h28 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_40_branch_valid <= _GEN_3462;
        end else begin
          memReg_40_branch_valid <= _GEN_3727;
        end
      end else begin
        memReg_40_branch_valid <= _GEN_3462;
      end
    end else begin
      memReg_40_branch_valid <= _GEN_3462;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_40_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h28 | 6'h28 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_40_branch_mask <= _GEN_3726;
        end else begin
          memReg_40_branch_mask <= _GEN_3398;
        end
      end else begin
        memReg_40_branch_mask <= _GEN_3398;
      end
    end else begin
      memReg_40_branch_mask <= _GEN_3398;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_41_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_41_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_41_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_41_valid <= _GEN_839;
      end
    end else begin
      memReg_41_valid <= _GEN_839;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_41_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h29 == writePtr) begin // @[fifo.scala 82:22]
        memReg_41_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_41_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h29 | 6'h29 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_41_branch_valid <= _GEN_3463;
        end else begin
          memReg_41_branch_valid <= _GEN_3733;
        end
      end else begin
        memReg_41_branch_valid <= _GEN_3463;
      end
    end else begin
      memReg_41_branch_valid <= _GEN_3463;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_41_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h29 | 6'h29 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_41_branch_mask <= _GEN_3732;
        end else begin
          memReg_41_branch_mask <= _GEN_3399;
        end
      end else begin
        memReg_41_branch_mask <= _GEN_3399;
      end
    end else begin
      memReg_41_branch_mask <= _GEN_3399;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_42_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_42_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_42_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_42_valid <= _GEN_840;
      end
    end else begin
      memReg_42_valid <= _GEN_840;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_42_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h2a == writePtr) begin // @[fifo.scala 82:22]
        memReg_42_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_42_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h2a | 6'h2a <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_42_branch_valid <= _GEN_3464;
        end else begin
          memReg_42_branch_valid <= _GEN_3739;
        end
      end else begin
        memReg_42_branch_valid <= _GEN_3464;
      end
    end else begin
      memReg_42_branch_valid <= _GEN_3464;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_42_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h2a | 6'h2a <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_42_branch_mask <= _GEN_3738;
        end else begin
          memReg_42_branch_mask <= _GEN_3400;
        end
      end else begin
        memReg_42_branch_mask <= _GEN_3400;
      end
    end else begin
      memReg_42_branch_mask <= _GEN_3400;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_43_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_43_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_43_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_43_valid <= _GEN_841;
      end
    end else begin
      memReg_43_valid <= _GEN_841;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_43_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h2b == writePtr) begin // @[fifo.scala 82:22]
        memReg_43_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_43_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h2b | 6'h2b <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_43_branch_valid <= _GEN_3465;
        end else begin
          memReg_43_branch_valid <= _GEN_3745;
        end
      end else begin
        memReg_43_branch_valid <= _GEN_3465;
      end
    end else begin
      memReg_43_branch_valid <= _GEN_3465;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_43_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h2b | 6'h2b <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_43_branch_mask <= _GEN_3744;
        end else begin
          memReg_43_branch_mask <= _GEN_3401;
        end
      end else begin
        memReg_43_branch_mask <= _GEN_3401;
      end
    end else begin
      memReg_43_branch_mask <= _GEN_3401;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_44_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_44_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_44_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_44_valid <= _GEN_842;
      end
    end else begin
      memReg_44_valid <= _GEN_842;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_44_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h2c == writePtr) begin // @[fifo.scala 82:22]
        memReg_44_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_44_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h2c | 6'h2c <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_44_branch_valid <= _GEN_3466;
        end else begin
          memReg_44_branch_valid <= _GEN_3751;
        end
      end else begin
        memReg_44_branch_valid <= _GEN_3466;
      end
    end else begin
      memReg_44_branch_valid <= _GEN_3466;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_44_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h2c | 6'h2c <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_44_branch_mask <= _GEN_3750;
        end else begin
          memReg_44_branch_mask <= _GEN_3402;
        end
      end else begin
        memReg_44_branch_mask <= _GEN_3402;
      end
    end else begin
      memReg_44_branch_mask <= _GEN_3402;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_45_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_45_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_45_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_45_valid <= _GEN_843;
      end
    end else begin
      memReg_45_valid <= _GEN_843;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_45_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h2d == writePtr) begin // @[fifo.scala 82:22]
        memReg_45_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_45_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h2d | 6'h2d <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_45_branch_valid <= _GEN_3467;
        end else begin
          memReg_45_branch_valid <= _GEN_3757;
        end
      end else begin
        memReg_45_branch_valid <= _GEN_3467;
      end
    end else begin
      memReg_45_branch_valid <= _GEN_3467;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_45_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h2d | 6'h2d <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_45_branch_mask <= _GEN_3756;
        end else begin
          memReg_45_branch_mask <= _GEN_3403;
        end
      end else begin
        memReg_45_branch_mask <= _GEN_3403;
      end
    end else begin
      memReg_45_branch_mask <= _GEN_3403;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_46_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_46_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_46_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_46_valid <= _GEN_844;
      end
    end else begin
      memReg_46_valid <= _GEN_844;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_46_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h2e == writePtr) begin // @[fifo.scala 82:22]
        memReg_46_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_46_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h2e | 6'h2e <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_46_branch_valid <= _GEN_3468;
        end else begin
          memReg_46_branch_valid <= _GEN_3763;
        end
      end else begin
        memReg_46_branch_valid <= _GEN_3468;
      end
    end else begin
      memReg_46_branch_valid <= _GEN_3468;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_46_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h2e | 6'h2e <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_46_branch_mask <= _GEN_3762;
        end else begin
          memReg_46_branch_mask <= _GEN_3404;
        end
      end else begin
        memReg_46_branch_mask <= _GEN_3404;
      end
    end else begin
      memReg_46_branch_mask <= _GEN_3404;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_47_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_47_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_47_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_47_valid <= _GEN_845;
      end
    end else begin
      memReg_47_valid <= _GEN_845;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_47_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h2f == writePtr) begin // @[fifo.scala 82:22]
        memReg_47_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_47_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h2f | 6'h2f <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_47_branch_valid <= _GEN_3469;
        end else begin
          memReg_47_branch_valid <= _GEN_3769;
        end
      end else begin
        memReg_47_branch_valid <= _GEN_3469;
      end
    end else begin
      memReg_47_branch_valid <= _GEN_3469;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_47_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h2f | 6'h2f <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_47_branch_mask <= _GEN_3768;
        end else begin
          memReg_47_branch_mask <= _GEN_3405;
        end
      end else begin
        memReg_47_branch_mask <= _GEN_3405;
      end
    end else begin
      memReg_47_branch_mask <= _GEN_3405;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_48_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_48_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_48_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_48_valid <= _GEN_846;
      end
    end else begin
      memReg_48_valid <= _GEN_846;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_48_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h30 == writePtr) begin // @[fifo.scala 82:22]
        memReg_48_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_48_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h30 | 6'h30 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_48_branch_valid <= _GEN_3470;
        end else begin
          memReg_48_branch_valid <= _GEN_3775;
        end
      end else begin
        memReg_48_branch_valid <= _GEN_3470;
      end
    end else begin
      memReg_48_branch_valid <= _GEN_3470;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_48_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h30 | 6'h30 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_48_branch_mask <= _GEN_3774;
        end else begin
          memReg_48_branch_mask <= _GEN_3406;
        end
      end else begin
        memReg_48_branch_mask <= _GEN_3406;
      end
    end else begin
      memReg_48_branch_mask <= _GEN_3406;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_49_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_49_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_49_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_49_valid <= _GEN_847;
      end
    end else begin
      memReg_49_valid <= _GEN_847;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_49_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h31 == writePtr) begin // @[fifo.scala 82:22]
        memReg_49_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_49_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h31 | 6'h31 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_49_branch_valid <= _GEN_3471;
        end else begin
          memReg_49_branch_valid <= _GEN_3781;
        end
      end else begin
        memReg_49_branch_valid <= _GEN_3471;
      end
    end else begin
      memReg_49_branch_valid <= _GEN_3471;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_49_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h31 | 6'h31 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_49_branch_mask <= _GEN_3780;
        end else begin
          memReg_49_branch_mask <= _GEN_3407;
        end
      end else begin
        memReg_49_branch_mask <= _GEN_3407;
      end
    end else begin
      memReg_49_branch_mask <= _GEN_3407;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_50_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_50_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_50_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_50_valid <= _GEN_848;
      end
    end else begin
      memReg_50_valid <= _GEN_848;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_50_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h32 == writePtr) begin // @[fifo.scala 82:22]
        memReg_50_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_50_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h32 | 6'h32 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_50_branch_valid <= _GEN_3472;
        end else begin
          memReg_50_branch_valid <= _GEN_3787;
        end
      end else begin
        memReg_50_branch_valid <= _GEN_3472;
      end
    end else begin
      memReg_50_branch_valid <= _GEN_3472;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_50_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h32 | 6'h32 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_50_branch_mask <= _GEN_3786;
        end else begin
          memReg_50_branch_mask <= _GEN_3408;
        end
      end else begin
        memReg_50_branch_mask <= _GEN_3408;
      end
    end else begin
      memReg_50_branch_mask <= _GEN_3408;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_51_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_51_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_51_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_51_valid <= _GEN_849;
      end
    end else begin
      memReg_51_valid <= _GEN_849;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_51_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h33 == writePtr) begin // @[fifo.scala 82:22]
        memReg_51_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_51_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h33 | 6'h33 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_51_branch_valid <= _GEN_3473;
        end else begin
          memReg_51_branch_valid <= _GEN_3793;
        end
      end else begin
        memReg_51_branch_valid <= _GEN_3473;
      end
    end else begin
      memReg_51_branch_valid <= _GEN_3473;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_51_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h33 | 6'h33 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_51_branch_mask <= _GEN_3792;
        end else begin
          memReg_51_branch_mask <= _GEN_3409;
        end
      end else begin
        memReg_51_branch_mask <= _GEN_3409;
      end
    end else begin
      memReg_51_branch_mask <= _GEN_3409;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_52_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_52_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_52_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_52_valid <= _GEN_850;
      end
    end else begin
      memReg_52_valid <= _GEN_850;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_52_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h34 == writePtr) begin // @[fifo.scala 82:22]
        memReg_52_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_52_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h34 | 6'h34 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_52_branch_valid <= _GEN_3474;
        end else begin
          memReg_52_branch_valid <= _GEN_3799;
        end
      end else begin
        memReg_52_branch_valid <= _GEN_3474;
      end
    end else begin
      memReg_52_branch_valid <= _GEN_3474;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_52_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h34 | 6'h34 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_52_branch_mask <= _GEN_3798;
        end else begin
          memReg_52_branch_mask <= _GEN_3410;
        end
      end else begin
        memReg_52_branch_mask <= _GEN_3410;
      end
    end else begin
      memReg_52_branch_mask <= _GEN_3410;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_53_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_53_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_53_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_53_valid <= _GEN_851;
      end
    end else begin
      memReg_53_valid <= _GEN_851;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_53_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h35 == writePtr) begin // @[fifo.scala 82:22]
        memReg_53_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_53_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h35 | 6'h35 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_53_branch_valid <= _GEN_3475;
        end else begin
          memReg_53_branch_valid <= _GEN_3805;
        end
      end else begin
        memReg_53_branch_valid <= _GEN_3475;
      end
    end else begin
      memReg_53_branch_valid <= _GEN_3475;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_53_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h35 | 6'h35 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_53_branch_mask <= _GEN_3804;
        end else begin
          memReg_53_branch_mask <= _GEN_3411;
        end
      end else begin
        memReg_53_branch_mask <= _GEN_3411;
      end
    end else begin
      memReg_53_branch_mask <= _GEN_3411;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_54_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_54_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_54_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_54_valid <= _GEN_852;
      end
    end else begin
      memReg_54_valid <= _GEN_852;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_54_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h36 == writePtr) begin // @[fifo.scala 82:22]
        memReg_54_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_54_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h36 | 6'h36 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_54_branch_valid <= _GEN_3476;
        end else begin
          memReg_54_branch_valid <= _GEN_3811;
        end
      end else begin
        memReg_54_branch_valid <= _GEN_3476;
      end
    end else begin
      memReg_54_branch_valid <= _GEN_3476;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_54_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h36 | 6'h36 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_54_branch_mask <= _GEN_3810;
        end else begin
          memReg_54_branch_mask <= _GEN_3412;
        end
      end else begin
        memReg_54_branch_mask <= _GEN_3412;
      end
    end else begin
      memReg_54_branch_mask <= _GEN_3412;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_55_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_55_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_55_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_55_valid <= _GEN_853;
      end
    end else begin
      memReg_55_valid <= _GEN_853;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_55_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h37 == writePtr) begin // @[fifo.scala 82:22]
        memReg_55_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_55_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h37 | 6'h37 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_55_branch_valid <= _GEN_3477;
        end else begin
          memReg_55_branch_valid <= _GEN_3817;
        end
      end else begin
        memReg_55_branch_valid <= _GEN_3477;
      end
    end else begin
      memReg_55_branch_valid <= _GEN_3477;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_55_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h37 | 6'h37 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_55_branch_mask <= _GEN_3816;
        end else begin
          memReg_55_branch_mask <= _GEN_3413;
        end
      end else begin
        memReg_55_branch_mask <= _GEN_3413;
      end
    end else begin
      memReg_55_branch_mask <= _GEN_3413;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_56_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_56_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_56_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_56_valid <= _GEN_854;
      end
    end else begin
      memReg_56_valid <= _GEN_854;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_56_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h38 == writePtr) begin // @[fifo.scala 82:22]
        memReg_56_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_56_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h38 | 6'h38 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_56_branch_valid <= _GEN_3478;
        end else begin
          memReg_56_branch_valid <= _GEN_3823;
        end
      end else begin
        memReg_56_branch_valid <= _GEN_3478;
      end
    end else begin
      memReg_56_branch_valid <= _GEN_3478;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_56_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h38 | 6'h38 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_56_branch_mask <= _GEN_3822;
        end else begin
          memReg_56_branch_mask <= _GEN_3414;
        end
      end else begin
        memReg_56_branch_mask <= _GEN_3414;
      end
    end else begin
      memReg_56_branch_mask <= _GEN_3414;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_57_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_57_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_57_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_57_valid <= _GEN_855;
      end
    end else begin
      memReg_57_valid <= _GEN_855;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_57_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h39 == writePtr) begin // @[fifo.scala 82:22]
        memReg_57_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_57_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h39 | 6'h39 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_57_branch_valid <= _GEN_3479;
        end else begin
          memReg_57_branch_valid <= _GEN_3829;
        end
      end else begin
        memReg_57_branch_valid <= _GEN_3479;
      end
    end else begin
      memReg_57_branch_valid <= _GEN_3479;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_57_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h39 | 6'h39 <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_57_branch_mask <= _GEN_3828;
        end else begin
          memReg_57_branch_mask <= _GEN_3415;
        end
      end else begin
        memReg_57_branch_mask <= _GEN_3415;
      end
    end else begin
      memReg_57_branch_mask <= _GEN_3415;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_58_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_58_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_58_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_58_valid <= _GEN_856;
      end
    end else begin
      memReg_58_valid <= _GEN_856;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_58_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h3a == writePtr) begin // @[fifo.scala 82:22]
        memReg_58_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_58_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h3a | 6'h3a <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_58_branch_valid <= _GEN_3480;
        end else begin
          memReg_58_branch_valid <= _GEN_3835;
        end
      end else begin
        memReg_58_branch_valid <= _GEN_3480;
      end
    end else begin
      memReg_58_branch_valid <= _GEN_3480;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_58_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h3a | 6'h3a <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_58_branch_mask <= _GEN_3834;
        end else begin
          memReg_58_branch_mask <= _GEN_3416;
        end
      end else begin
        memReg_58_branch_mask <= _GEN_3416;
      end
    end else begin
      memReg_58_branch_mask <= _GEN_3416;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_59_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_59_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_59_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_59_valid <= _GEN_857;
      end
    end else begin
      memReg_59_valid <= _GEN_857;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_59_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h3b == writePtr) begin // @[fifo.scala 82:22]
        memReg_59_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_59_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h3b | 6'h3b <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_59_branch_valid <= _GEN_3481;
        end else begin
          memReg_59_branch_valid <= _GEN_3841;
        end
      end else begin
        memReg_59_branch_valid <= _GEN_3481;
      end
    end else begin
      memReg_59_branch_valid <= _GEN_3481;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_59_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h3b | 6'h3b <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_59_branch_mask <= _GEN_3840;
        end else begin
          memReg_59_branch_mask <= _GEN_3417;
        end
      end else begin
        memReg_59_branch_mask <= _GEN_3417;
      end
    end else begin
      memReg_59_branch_mask <= _GEN_3417;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_60_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_60_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_60_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_60_valid <= _GEN_858;
      end
    end else begin
      memReg_60_valid <= _GEN_858;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_60_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h3c == writePtr) begin // @[fifo.scala 82:22]
        memReg_60_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_60_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h3c | 6'h3c <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_60_branch_valid <= _GEN_3482;
        end else begin
          memReg_60_branch_valid <= _GEN_3847;
        end
      end else begin
        memReg_60_branch_valid <= _GEN_3482;
      end
    end else begin
      memReg_60_branch_valid <= _GEN_3482;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_60_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h3c | 6'h3c <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_60_branch_mask <= _GEN_3846;
        end else begin
          memReg_60_branch_mask <= _GEN_3418;
        end
      end else begin
        memReg_60_branch_mask <= _GEN_3418;
      end
    end else begin
      memReg_60_branch_mask <= _GEN_3418;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_61_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_61_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_61_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_61_valid <= _GEN_859;
      end
    end else begin
      memReg_61_valid <= _GEN_859;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_61_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h3d == writePtr) begin // @[fifo.scala 82:22]
        memReg_61_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_61_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h3d | 6'h3d <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_61_branch_valid <= _GEN_3483;
        end else begin
          memReg_61_branch_valid <= _GEN_3853;
        end
      end else begin
        memReg_61_branch_valid <= _GEN_3483;
      end
    end else begin
      memReg_61_branch_valid <= _GEN_3483;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_61_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h3d | 6'h3d <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_61_branch_mask <= _GEN_3852;
        end else begin
          memReg_61_branch_mask <= _GEN_3419;
        end
      end else begin
        memReg_61_branch_mask <= _GEN_3419;
      end
    end else begin
      memReg_61_branch_mask <= _GEN_3419;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_62_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_62_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_62_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_62_valid <= _GEN_860;
      end
    end else begin
      memReg_62_valid <= _GEN_860;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_62_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h3e == writePtr) begin // @[fifo.scala 82:22]
        memReg_62_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_62_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h3e | 6'h3e <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_62_branch_valid <= _GEN_3484;
        end else begin
          memReg_62_branch_valid <= _GEN_3859;
        end
      end else begin
        memReg_62_branch_valid <= _GEN_3484;
      end
    end else begin
      memReg_62_branch_valid <= _GEN_3484;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_62_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (startPointer <= 6'h3e | 6'h3e <= endPointer) begin // @[fifo.scala 107:54]
        if (branchOps_passed) begin // @[fifo.scala 108:32]
          memReg_62_branch_mask <= _GEN_3858;
        end else begin
          memReg_62_branch_mask <= _GEN_3420;
        end
      end else begin
        memReg_62_branch_mask <= _GEN_3420;
      end
    end else begin
      memReg_62_branch_mask <= _GEN_3420;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_63_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (invalidateEnable) begin // @[fifo.scala 141:26]
      if (memReg_63_address == invalidateAddr) begin // @[fifo.scala 143:50]
        memReg_63_valid <= 1'h0; // @[fifo.scala 144:25]
      end else begin
        memReg_63_valid <= _GEN_861;
      end
    end else begin
      memReg_63_valid <= _GEN_861;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_63_address <= 32'h0; // @[fifo.scala 27:33]
    end else if (incrWrite) begin // @[fifo.scala 81:17]
      if (6'h3f == writePtr) begin // @[fifo.scala 82:22]
        memReg_63_address <= write_data_address; // @[fifo.scala 82:22]
      end
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_63_branch_valid <= 1'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (branchOps_passed) begin // @[fifo.scala 108:32]
        memReg_63_branch_valid <= _GEN_3485;
      end else if (_T_457) begin // @[fifo.scala 113:68]
        memReg_63_branch_valid <= 1'h0; // @[fifo.scala 114:36]
      end else begin
        memReg_63_branch_valid <= _GEN_3485;
      end
    end else begin
      memReg_63_branch_valid <= _GEN_3485;
    end
    if (reset) begin // @[fifo.scala 27:33]
      memReg_63_branch_mask <= 5'h0; // @[fifo.scala 27:33]
    end else if (branchOps_valid) begin // @[fifo.scala 105:25]
      if (branchOps_passed) begin // @[fifo.scala 108:32]
        if (|_T_456) begin // @[fifo.scala 109:68]
          memReg_63_branch_mask <= _memReg_63_branch_mask_T; // @[fifo.scala 110:35]
        end else begin
          memReg_63_branch_mask <= _GEN_3421;
        end
      end else begin
        memReg_63_branch_mask <= _GEN_3421;
      end
    end else begin
      memReg_63_branch_mask <= _GEN_3421;
    end
    if (reset) begin // @[fifo.scala 33:25]
      readPtr <= 6'h0; // @[fifo.scala 33:25]
    end else if (incrRead) begin // @[fifo.scala 35:15]
      if (readPtr == 6'h3f) begin // @[fifo.scala 34:22]
        readPtr <= 6'h0;
      end else begin
        readPtr <= _nextVal_T_2;
      end
    end
    emptyReg <= reset | _GEN_27; // @[fifo.scala 43:{25,25}]
    if (reset) begin // @[fifo.scala 33:25]
      writePtr <= 6'h0; // @[fifo.scala 33:25]
    end else if (incrWrite) begin // @[fifo.scala 35:15]
      if (writePtr == 6'h3f) begin // @[fifo.scala 34:22]
        writePtr <= 6'h0;
      end else begin
        writePtr <= _nextVal_T_5;
      end
    end
    if (reset) begin // @[fifo.scala 44:34]
      fullReg <= 1'h0; // @[fifo.scala 44:34]
    end else if (!(2'h0 == op)) begin // @[fifo.scala 49:14]
      if (2'h1 == op) begin // @[fifo.scala 49:14]
        if (~emptyReg) begin // @[fifo.scala 52:23]
          fullReg <= 1'h0; // @[fifo.scala 53:17]
        end
      end else if (2'h2 == op) begin // @[fifo.scala 49:14]
        fullReg <= _GEN_7;
      end else begin
        fullReg <= _GEN_16;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  memReg_0_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  memReg_0_address = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  memReg_0_branch_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  memReg_0_branch_mask = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  memReg_1_valid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  memReg_1_address = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  memReg_1_branch_valid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  memReg_1_branch_mask = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  memReg_2_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  memReg_2_address = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  memReg_2_branch_valid = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  memReg_2_branch_mask = _RAND_11[4:0];
  _RAND_12 = {1{`RANDOM}};
  memReg_3_valid = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  memReg_3_address = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  memReg_3_branch_valid = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  memReg_3_branch_mask = _RAND_15[4:0];
  _RAND_16 = {1{`RANDOM}};
  memReg_4_valid = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  memReg_4_address = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  memReg_4_branch_valid = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  memReg_4_branch_mask = _RAND_19[4:0];
  _RAND_20 = {1{`RANDOM}};
  memReg_5_valid = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  memReg_5_address = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  memReg_5_branch_valid = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  memReg_5_branch_mask = _RAND_23[4:0];
  _RAND_24 = {1{`RANDOM}};
  memReg_6_valid = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  memReg_6_address = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  memReg_6_branch_valid = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  memReg_6_branch_mask = _RAND_27[4:0];
  _RAND_28 = {1{`RANDOM}};
  memReg_7_valid = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  memReg_7_address = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  memReg_7_branch_valid = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  memReg_7_branch_mask = _RAND_31[4:0];
  _RAND_32 = {1{`RANDOM}};
  memReg_8_valid = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  memReg_8_address = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  memReg_8_branch_valid = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  memReg_8_branch_mask = _RAND_35[4:0];
  _RAND_36 = {1{`RANDOM}};
  memReg_9_valid = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  memReg_9_address = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  memReg_9_branch_valid = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  memReg_9_branch_mask = _RAND_39[4:0];
  _RAND_40 = {1{`RANDOM}};
  memReg_10_valid = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  memReg_10_address = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  memReg_10_branch_valid = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  memReg_10_branch_mask = _RAND_43[4:0];
  _RAND_44 = {1{`RANDOM}};
  memReg_11_valid = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  memReg_11_address = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  memReg_11_branch_valid = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  memReg_11_branch_mask = _RAND_47[4:0];
  _RAND_48 = {1{`RANDOM}};
  memReg_12_valid = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  memReg_12_address = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  memReg_12_branch_valid = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  memReg_12_branch_mask = _RAND_51[4:0];
  _RAND_52 = {1{`RANDOM}};
  memReg_13_valid = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  memReg_13_address = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  memReg_13_branch_valid = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  memReg_13_branch_mask = _RAND_55[4:0];
  _RAND_56 = {1{`RANDOM}};
  memReg_14_valid = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  memReg_14_address = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  memReg_14_branch_valid = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  memReg_14_branch_mask = _RAND_59[4:0];
  _RAND_60 = {1{`RANDOM}};
  memReg_15_valid = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  memReg_15_address = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  memReg_15_branch_valid = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  memReg_15_branch_mask = _RAND_63[4:0];
  _RAND_64 = {1{`RANDOM}};
  memReg_16_valid = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  memReg_16_address = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  memReg_16_branch_valid = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  memReg_16_branch_mask = _RAND_67[4:0];
  _RAND_68 = {1{`RANDOM}};
  memReg_17_valid = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  memReg_17_address = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  memReg_17_branch_valid = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  memReg_17_branch_mask = _RAND_71[4:0];
  _RAND_72 = {1{`RANDOM}};
  memReg_18_valid = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  memReg_18_address = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  memReg_18_branch_valid = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  memReg_18_branch_mask = _RAND_75[4:0];
  _RAND_76 = {1{`RANDOM}};
  memReg_19_valid = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  memReg_19_address = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  memReg_19_branch_valid = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  memReg_19_branch_mask = _RAND_79[4:0];
  _RAND_80 = {1{`RANDOM}};
  memReg_20_valid = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  memReg_20_address = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  memReg_20_branch_valid = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  memReg_20_branch_mask = _RAND_83[4:0];
  _RAND_84 = {1{`RANDOM}};
  memReg_21_valid = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  memReg_21_address = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  memReg_21_branch_valid = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  memReg_21_branch_mask = _RAND_87[4:0];
  _RAND_88 = {1{`RANDOM}};
  memReg_22_valid = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  memReg_22_address = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  memReg_22_branch_valid = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  memReg_22_branch_mask = _RAND_91[4:0];
  _RAND_92 = {1{`RANDOM}};
  memReg_23_valid = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  memReg_23_address = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  memReg_23_branch_valid = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  memReg_23_branch_mask = _RAND_95[4:0];
  _RAND_96 = {1{`RANDOM}};
  memReg_24_valid = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  memReg_24_address = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  memReg_24_branch_valid = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  memReg_24_branch_mask = _RAND_99[4:0];
  _RAND_100 = {1{`RANDOM}};
  memReg_25_valid = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  memReg_25_address = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  memReg_25_branch_valid = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  memReg_25_branch_mask = _RAND_103[4:0];
  _RAND_104 = {1{`RANDOM}};
  memReg_26_valid = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  memReg_26_address = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  memReg_26_branch_valid = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  memReg_26_branch_mask = _RAND_107[4:0];
  _RAND_108 = {1{`RANDOM}};
  memReg_27_valid = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  memReg_27_address = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  memReg_27_branch_valid = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  memReg_27_branch_mask = _RAND_111[4:0];
  _RAND_112 = {1{`RANDOM}};
  memReg_28_valid = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  memReg_28_address = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  memReg_28_branch_valid = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  memReg_28_branch_mask = _RAND_115[4:0];
  _RAND_116 = {1{`RANDOM}};
  memReg_29_valid = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  memReg_29_address = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  memReg_29_branch_valid = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  memReg_29_branch_mask = _RAND_119[4:0];
  _RAND_120 = {1{`RANDOM}};
  memReg_30_valid = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  memReg_30_address = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  memReg_30_branch_valid = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  memReg_30_branch_mask = _RAND_123[4:0];
  _RAND_124 = {1{`RANDOM}};
  memReg_31_valid = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  memReg_31_address = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  memReg_31_branch_valid = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  memReg_31_branch_mask = _RAND_127[4:0];
  _RAND_128 = {1{`RANDOM}};
  memReg_32_valid = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  memReg_32_address = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  memReg_32_branch_valid = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  memReg_32_branch_mask = _RAND_131[4:0];
  _RAND_132 = {1{`RANDOM}};
  memReg_33_valid = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  memReg_33_address = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  memReg_33_branch_valid = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  memReg_33_branch_mask = _RAND_135[4:0];
  _RAND_136 = {1{`RANDOM}};
  memReg_34_valid = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  memReg_34_address = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  memReg_34_branch_valid = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  memReg_34_branch_mask = _RAND_139[4:0];
  _RAND_140 = {1{`RANDOM}};
  memReg_35_valid = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  memReg_35_address = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  memReg_35_branch_valid = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  memReg_35_branch_mask = _RAND_143[4:0];
  _RAND_144 = {1{`RANDOM}};
  memReg_36_valid = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  memReg_36_address = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  memReg_36_branch_valid = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  memReg_36_branch_mask = _RAND_147[4:0];
  _RAND_148 = {1{`RANDOM}};
  memReg_37_valid = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  memReg_37_address = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  memReg_37_branch_valid = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  memReg_37_branch_mask = _RAND_151[4:0];
  _RAND_152 = {1{`RANDOM}};
  memReg_38_valid = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  memReg_38_address = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  memReg_38_branch_valid = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  memReg_38_branch_mask = _RAND_155[4:0];
  _RAND_156 = {1{`RANDOM}};
  memReg_39_valid = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  memReg_39_address = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  memReg_39_branch_valid = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  memReg_39_branch_mask = _RAND_159[4:0];
  _RAND_160 = {1{`RANDOM}};
  memReg_40_valid = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  memReg_40_address = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  memReg_40_branch_valid = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  memReg_40_branch_mask = _RAND_163[4:0];
  _RAND_164 = {1{`RANDOM}};
  memReg_41_valid = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  memReg_41_address = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  memReg_41_branch_valid = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  memReg_41_branch_mask = _RAND_167[4:0];
  _RAND_168 = {1{`RANDOM}};
  memReg_42_valid = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  memReg_42_address = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  memReg_42_branch_valid = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  memReg_42_branch_mask = _RAND_171[4:0];
  _RAND_172 = {1{`RANDOM}};
  memReg_43_valid = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  memReg_43_address = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  memReg_43_branch_valid = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  memReg_43_branch_mask = _RAND_175[4:0];
  _RAND_176 = {1{`RANDOM}};
  memReg_44_valid = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  memReg_44_address = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  memReg_44_branch_valid = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  memReg_44_branch_mask = _RAND_179[4:0];
  _RAND_180 = {1{`RANDOM}};
  memReg_45_valid = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  memReg_45_address = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  memReg_45_branch_valid = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  memReg_45_branch_mask = _RAND_183[4:0];
  _RAND_184 = {1{`RANDOM}};
  memReg_46_valid = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  memReg_46_address = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  memReg_46_branch_valid = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  memReg_46_branch_mask = _RAND_187[4:0];
  _RAND_188 = {1{`RANDOM}};
  memReg_47_valid = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  memReg_47_address = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  memReg_47_branch_valid = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  memReg_47_branch_mask = _RAND_191[4:0];
  _RAND_192 = {1{`RANDOM}};
  memReg_48_valid = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  memReg_48_address = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  memReg_48_branch_valid = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  memReg_48_branch_mask = _RAND_195[4:0];
  _RAND_196 = {1{`RANDOM}};
  memReg_49_valid = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  memReg_49_address = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  memReg_49_branch_valid = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  memReg_49_branch_mask = _RAND_199[4:0];
  _RAND_200 = {1{`RANDOM}};
  memReg_50_valid = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  memReg_50_address = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  memReg_50_branch_valid = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  memReg_50_branch_mask = _RAND_203[4:0];
  _RAND_204 = {1{`RANDOM}};
  memReg_51_valid = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  memReg_51_address = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  memReg_51_branch_valid = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  memReg_51_branch_mask = _RAND_207[4:0];
  _RAND_208 = {1{`RANDOM}};
  memReg_52_valid = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  memReg_52_address = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  memReg_52_branch_valid = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  memReg_52_branch_mask = _RAND_211[4:0];
  _RAND_212 = {1{`RANDOM}};
  memReg_53_valid = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  memReg_53_address = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  memReg_53_branch_valid = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  memReg_53_branch_mask = _RAND_215[4:0];
  _RAND_216 = {1{`RANDOM}};
  memReg_54_valid = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  memReg_54_address = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  memReg_54_branch_valid = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  memReg_54_branch_mask = _RAND_219[4:0];
  _RAND_220 = {1{`RANDOM}};
  memReg_55_valid = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  memReg_55_address = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  memReg_55_branch_valid = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  memReg_55_branch_mask = _RAND_223[4:0];
  _RAND_224 = {1{`RANDOM}};
  memReg_56_valid = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  memReg_56_address = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  memReg_56_branch_valid = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  memReg_56_branch_mask = _RAND_227[4:0];
  _RAND_228 = {1{`RANDOM}};
  memReg_57_valid = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  memReg_57_address = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  memReg_57_branch_valid = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  memReg_57_branch_mask = _RAND_231[4:0];
  _RAND_232 = {1{`RANDOM}};
  memReg_58_valid = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  memReg_58_address = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  memReg_58_branch_valid = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  memReg_58_branch_mask = _RAND_235[4:0];
  _RAND_236 = {1{`RANDOM}};
  memReg_59_valid = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  memReg_59_address = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  memReg_59_branch_valid = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  memReg_59_branch_mask = _RAND_239[4:0];
  _RAND_240 = {1{`RANDOM}};
  memReg_60_valid = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  memReg_60_address = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  memReg_60_branch_valid = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  memReg_60_branch_mask = _RAND_243[4:0];
  _RAND_244 = {1{`RANDOM}};
  memReg_61_valid = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  memReg_61_address = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  memReg_61_branch_valid = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  memReg_61_branch_mask = _RAND_247[4:0];
  _RAND_248 = {1{`RANDOM}};
  memReg_62_valid = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  memReg_62_address = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  memReg_62_branch_valid = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  memReg_62_branch_mask = _RAND_251[4:0];
  _RAND_252 = {1{`RANDOM}};
  memReg_63_valid = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  memReg_63_address = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  memReg_63_branch_valid = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  memReg_63_branch_mask = _RAND_255[4:0];
  _RAND_256 = {1{`RANDOM}};
  readPtr = _RAND_256[5:0];
  _RAND_257 = {1{`RANDOM}};
  emptyReg = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  writePtr = _RAND_258[5:0];
  _RAND_259 = {1{`RANDOM}};
  fullReg = _RAND_259[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module core_Anon_1(
  input         clock,
  input         reset,
  input         request_valid,
  input  [31:0] request_address,
  input  [31:0] request_instruction,
  input  [4:0]  request_branchMask,
  input  [3:0]  request_robAddr,
  input  [5:0]  request_prfDest,
  output [31:0] dPort_AWADDR,
  output        dPort_AWVALID,
  input         dPort_AWREADY,
  output [63:0] dPort_WDATA,
  output        dPort_WLAST,
  output        dPort_WVALID,
  input         dPort_WREADY,
  input  [1:0]  dPort_BRESP,
  input         dPort_BVALID,
  output        dPort_BREADY,
  output [31:0] dPort_ARADDR,
  output        dPort_ARVALID,
  input         dPort_ARREADY,
  input  [63:0] dPort_RDATA,
  input         dPort_RLAST,
  input         dPort_RVALID,
  output        dPort_RREADY,
  output [2:0]  dPort_AWSNOOP,
  output [3:0]  dPort_ARSNOOP,
  input  [3:0]  dPort_RRESP,
  input         dPort_ACVALID,
  output        dPort_ACREADY,
  input  [31:0] dPort_ACADDR,
  input  [3:0]  dPort_ACSNOOP,
  output        dPort_CRVALID,
  input         dPort_CRREADY,
  output [4:0]  dPort_CRRESP,
  output        dPort_CDVALID,
  input         dPort_CDREADY,
  output [63:0] dPort_CDDATA,
  output        dPort_CDLAST,
  output [31:0] peripheral_AWADDR,
  output [7:0]  peripheral_AWLEN,
  output [2:0]  peripheral_AWSIZE,
  output [1:0]  peripheral_AWBURST,
  output [2:0]  peripheral_AWPROT,
  output        peripheral_AWVALID,
  input         peripheral_AWREADY,
  output [31:0] peripheral_WDATA,
  output [3:0]  peripheral_WSTRB,
  output        peripheral_WLAST,
  output        peripheral_WVALID,
  input         peripheral_WREADY,
  input  [1:0]  peripheral_BID,
  input  [1:0]  peripheral_BRESP,
  input         peripheral_BVALID,
  output        peripheral_BREADY,
  output [31:0] peripheral_ARADDR,
  output [7:0]  peripheral_ARLEN,
  output [2:0]  peripheral_ARSIZE,
  output [1:0]  peripheral_ARBURST,
  output [2:0]  peripheral_ARPROT,
  output        peripheral_ARVALID,
  input         peripheral_ARREADY,
  input  [1:0]  peripheral_RID,
  input  [31:0] peripheral_RDATA,
  input  [1:0]  peripheral_RRESP,
  input         peripheral_RLAST,
  input         peripheral_RVALID,
  output        peripheral_RREADY,
  output        responseOut_valid,
  output [5:0]  responseOut_prfDest,
  output [3:0]  responseOut_robAddr,
  output [63:0] responseOut_result,
  output [31:0] responseOut_instruction,
  output        canAllocate,
  input         writeDataIn_valid,
  input  [63:0] writeDataIn_data,
  input         initiateFence,
  output        fenceInstructions_ready,
  input         fenceInstructions_fired,
  output        writeCommit_ready,
  input         writeCommit_fired,
  output        writeInstructionCommit_ready,
  input         writeInstructionCommit_fired,
  input         branchOps_valid,
  input  [4:0]  branchOps_branchMask,
  input         branchOps_passed,
  input         loadCommit_ready,
  output        loadCommit_valid,
  output        loadCommit_state
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  requestScheduler_clock; // @[cacheModule.scala 48:32]
  wire  requestScheduler_reset; // @[cacheModule.scala 48:32]
  wire  requestScheduler_requestIn_valid; // @[cacheModule.scala 48:32]
  wire [31:0] requestScheduler_requestIn_address; // @[cacheModule.scala 48:32]
  wire [31:0] requestScheduler_requestIn_core_instruction; // @[cacheModule.scala 48:32]
  wire [3:0] requestScheduler_requestIn_core_robAddr; // @[cacheModule.scala 48:32]
  wire [5:0] requestScheduler_requestIn_core_prfDest; // @[cacheModule.scala 48:32]
  wire [4:0] requestScheduler_requestIn_branch_mask; // @[cacheModule.scala 48:32]
  wire  requestScheduler_canAllocate; // @[cacheModule.scala 48:32]
  wire  requestScheduler_requestOut_valid; // @[cacheModule.scala 48:32]
  wire [31:0] requestScheduler_requestOut_address; // @[cacheModule.scala 48:32]
  wire [31:0] requestScheduler_requestOut_core_instruction; // @[cacheModule.scala 48:32]
  wire [3:0] requestScheduler_requestOut_core_robAddr; // @[cacheModule.scala 48:32]
  wire [5:0] requestScheduler_requestOut_core_prfDest; // @[cacheModule.scala 48:32]
  wire  requestScheduler_requestOut_branch_valid; // @[cacheModule.scala 48:32]
  wire [4:0] requestScheduler_requestOut_branch_mask; // @[cacheModule.scala 48:32]
  wire  requestScheduler_requestOut_writeData_valid; // @[cacheModule.scala 48:32]
  wire [63:0] requestScheduler_requestOut_writeData_data; // @[cacheModule.scala 48:32]
  wire  requestScheduler_controlSignal_isSpeculative; // @[cacheModule.scala 48:32]
  wire  requestScheduler_controlSignal_inorderReady; // @[cacheModule.scala 48:32]
  wire  requestScheduler_controlSignal_speculativeReady; // @[cacheModule.scala 48:32]
  wire  requestScheduler_fenceReady; // @[cacheModule.scala 48:32]
  wire  requestScheduler_branchOps_valid; // @[cacheModule.scala 48:32]
  wire [4:0] requestScheduler_branchOps_branchMask; // @[cacheModule.scala 48:32]
  wire  requestScheduler_branchOps_passed; // @[cacheModule.scala 48:32]
  wire  arbiter_clock; // @[cacheModule.scala 49:23]
  wire  arbiter_reset; // @[cacheModule.scala 49:23]
  wire  arbiter_request_request_valid; // @[cacheModule.scala 49:23]
  wire [31:0] arbiter_request_request_address; // @[cacheModule.scala 49:23]
  wire [31:0] arbiter_request_request_core_instruction; // @[cacheModule.scala 49:23]
  wire [3:0] arbiter_request_request_core_robAddr; // @[cacheModule.scala 49:23]
  wire [5:0] arbiter_request_request_core_prfDest; // @[cacheModule.scala 49:23]
  wire  arbiter_request_request_branch_valid; // @[cacheModule.scala 49:23]
  wire [4:0] arbiter_request_request_branch_mask; // @[cacheModule.scala 49:23]
  wire  arbiter_request_request_writeData_valid; // @[cacheModule.scala 49:23]
  wire [63:0] arbiter_request_request_writeData_data; // @[cacheModule.scala 49:23]
  wire  arbiter_request_isSpeculative; // @[cacheModule.scala 49:23]
  wire  arbiter_request_inorderReady; // @[cacheModule.scala 49:23]
  wire  arbiter_request_speculativeReady; // @[cacheModule.scala 49:23]
  wire  arbiter_toPeripheral_ready; // @[cacheModule.scala 49:23]
  wire  arbiter_toPeripheral_request_valid; // @[cacheModule.scala 49:23]
  wire [31:0] arbiter_toPeripheral_request_address; // @[cacheModule.scala 49:23]
  wire [31:0] arbiter_toPeripheral_request_core_instruction; // @[cacheModule.scala 49:23]
  wire [3:0] arbiter_toPeripheral_request_core_robAddr; // @[cacheModule.scala 49:23]
  wire [5:0] arbiter_toPeripheral_request_core_prfDest; // @[cacheModule.scala 49:23]
  wire  arbiter_toPeripheral_request_branch_valid; // @[cacheModule.scala 49:23]
  wire [4:0] arbiter_toPeripheral_request_branch_mask; // @[cacheModule.scala 49:23]
  wire  arbiter_toPeripheral_request_writeData_valid; // @[cacheModule.scala 49:23]
  wire [63:0] arbiter_toPeripheral_request_writeData_data; // @[cacheModule.scala 49:23]
  wire  arbiter_toCacheLookup_ready; // @[cacheModule.scala 49:23]
  wire  arbiter_toCacheLookup_holdInOrder; // @[cacheModule.scala 49:23]
  wire [1:0] arbiter_toCacheLookup_requestType; // @[cacheModule.scala 49:23]
  wire  arbiter_toCacheLookup_request_valid; // @[cacheModule.scala 49:23]
  wire [31:0] arbiter_toCacheLookup_request_address; // @[cacheModule.scala 49:23]
  wire [31:0] arbiter_toCacheLookup_request_core_instruction; // @[cacheModule.scala 49:23]
  wire [3:0] arbiter_toCacheLookup_request_core_robAddr; // @[cacheModule.scala 49:23]
  wire [5:0] arbiter_toCacheLookup_request_core_prfDest; // @[cacheModule.scala 49:23]
  wire  arbiter_toCacheLookup_request_branch_valid; // @[cacheModule.scala 49:23]
  wire [4:0] arbiter_toCacheLookup_request_branch_mask; // @[cacheModule.scala 49:23]
  wire  arbiter_toCacheLookup_request_writeData_valid; // @[cacheModule.scala 49:23]
  wire [63:0] arbiter_toCacheLookup_request_writeData_data; // @[cacheModule.scala 49:23]
  wire [511:0] arbiter_toCacheLookup_request_cacheLine_cacheLine; // @[cacheModule.scala 49:23]
  wire [1:0] arbiter_toCacheLookup_request_cacheLine_response; // @[cacheModule.scala 49:23]
  wire  arbiter_replayRequest_ready; // @[cacheModule.scala 49:23]
  wire  arbiter_replayRequest_request_valid; // @[cacheModule.scala 49:23]
  wire [31:0] arbiter_replayRequest_request_address; // @[cacheModule.scala 49:23]
  wire [31:0] arbiter_replayRequest_request_core_instruction; // @[cacheModule.scala 49:23]
  wire [3:0] arbiter_replayRequest_request_core_robAddr; // @[cacheModule.scala 49:23]
  wire [5:0] arbiter_replayRequest_request_core_prfDest; // @[cacheModule.scala 49:23]
  wire  arbiter_replayRequest_request_branch_valid; // @[cacheModule.scala 49:23]
  wire [4:0] arbiter_replayRequest_request_branch_mask; // @[cacheModule.scala 49:23]
  wire  arbiter_replayRequest_request_writeData_valid; // @[cacheModule.scala 49:23]
  wire [63:0] arbiter_replayRequest_request_writeData_data; // @[cacheModule.scala 49:23]
  wire [511:0] arbiter_replayRequest_request_cacheLine_cacheLine; // @[cacheModule.scala 49:23]
  wire [1:0] arbiter_replayRequest_request_cacheLine_response; // @[cacheModule.scala 49:23]
  wire  arbiter_coherencyRequest_ready; // @[cacheModule.scala 49:23]
  wire  arbiter_coherencyRequest_request_valid; // @[cacheModule.scala 49:23]
  wire [31:0] arbiter_coherencyRequest_request_address; // @[cacheModule.scala 49:23]
  wire [1:0] arbiter_coherencyRequest_request_response; // @[cacheModule.scala 49:23]
  wire  arbiter_writeDataIn_valid; // @[cacheModule.scala 49:23]
  wire [63:0] arbiter_writeDataIn_data; // @[cacheModule.scala 49:23]
  wire  arbiter_writeCommit_ready; // @[cacheModule.scala 49:23]
  wire  arbiter_writeCommit_fired; // @[cacheModule.scala 49:23]
  wire  arbiter_branchOps_valid; // @[cacheModule.scala 49:23]
  wire [4:0] arbiter_branchOps_branchMask; // @[cacheModule.scala 49:23]
  wire  arbiter_branchOps_passed; // @[cacheModule.scala 49:23]
  wire  arbiter_responseOut_valid; // @[cacheModule.scala 49:23]
  wire [31:0] arbiter_responseOut_instruction; // @[cacheModule.scala 49:23]
  wire  arbiter_fenceReady; // @[cacheModule.scala 49:23]
  wire  arbiter_writeInstuctionCommitFired; // @[cacheModule.scala 49:23]
  wire  cacheLookup_clock; // @[cacheModule.scala 50:27]
  wire  cacheLookup_reset; // @[cacheModule.scala 50:27]
  wire  cacheLookup_request_ready; // @[cacheModule.scala 50:27]
  wire  cacheLookup_request_holdInOrder; // @[cacheModule.scala 50:27]
  wire [1:0] cacheLookup_request_requestType; // @[cacheModule.scala 50:27]
  wire  cacheLookup_request_request_valid; // @[cacheModule.scala 50:27]
  wire [31:0] cacheLookup_request_request_address; // @[cacheModule.scala 50:27]
  wire [31:0] cacheLookup_request_request_core_instruction; // @[cacheModule.scala 50:27]
  wire [3:0] cacheLookup_request_request_core_robAddr; // @[cacheModule.scala 50:27]
  wire [5:0] cacheLookup_request_request_core_prfDest; // @[cacheModule.scala 50:27]
  wire  cacheLookup_request_request_branch_valid; // @[cacheModule.scala 50:27]
  wire [4:0] cacheLookup_request_request_branch_mask; // @[cacheModule.scala 50:27]
  wire  cacheLookup_request_request_writeData_valid; // @[cacheModule.scala 50:27]
  wire [63:0] cacheLookup_request_request_writeData_data; // @[cacheModule.scala 50:27]
  wire [511:0] cacheLookup_request_request_cacheLine_cacheLine; // @[cacheModule.scala 50:27]
  wire [1:0] cacheLookup_request_request_cacheLine_response; // @[cacheModule.scala 50:27]
  wire  cacheLookup_toReplay_ready; // @[cacheModule.scala 50:27]
  wire  cacheLookup_toReplay_request_valid; // @[cacheModule.scala 50:27]
  wire [31:0] cacheLookup_toReplay_request_address; // @[cacheModule.scala 50:27]
  wire [31:0] cacheLookup_toReplay_request_core_instruction; // @[cacheModule.scala 50:27]
  wire [3:0] cacheLookup_toReplay_request_core_robAddr; // @[cacheModule.scala 50:27]
  wire [5:0] cacheLookup_toReplay_request_core_prfDest; // @[cacheModule.scala 50:27]
  wire  cacheLookup_toReplay_request_branch_valid; // @[cacheModule.scala 50:27]
  wire [4:0] cacheLookup_toReplay_request_branch_mask; // @[cacheModule.scala 50:27]
  wire  cacheLookup_toReplay_request_writeData_valid; // @[cacheModule.scala 50:27]
  wire [63:0] cacheLookup_toReplay_request_writeData_data; // @[cacheModule.scala 50:27]
  wire [1:0] cacheLookup_toReplay_request_cacheLine_response; // @[cacheModule.scala 50:27]
  wire  cacheLookup_toWriteBack_ready; // @[cacheModule.scala 50:27]
  wire  cacheLookup_toWriteBack_request_valid; // @[cacheModule.scala 50:27]
  wire [31:0] cacheLookup_toWriteBack_request_address; // @[cacheModule.scala 50:27]
  wire [511:0] cacheLookup_toWriteBack_request_data; // @[cacheModule.scala 50:27]
  wire  cacheLookup_toCoherency_ready; // @[cacheModule.scala 50:27]
  wire  cacheLookup_toCoherency_request_valid; // @[cacheModule.scala 50:27]
  wire [1:0] cacheLookup_toCoherency_request_response; // @[cacheModule.scala 50:27]
  wire [511:0] cacheLookup_toCoherency_request_cacheLine; // @[cacheModule.scala 50:27]
  wire  cacheLookup_toCoherency_request_dataValid; // @[cacheModule.scala 50:27]
  wire  cacheLookup_toResponse_request_valid; // @[cacheModule.scala 50:27]
  wire [31:0] cacheLookup_toResponse_request_address; // @[cacheModule.scala 50:27]
  wire [31:0] cacheLookup_toResponse_request_core_instruction; // @[cacheModule.scala 50:27]
  wire [3:0] cacheLookup_toResponse_request_core_robAddr; // @[cacheModule.scala 50:27]
  wire [5:0] cacheLookup_toResponse_request_core_prfDest; // @[cacheModule.scala 50:27]
  wire  cacheLookup_toResponse_request_branch_valid; // @[cacheModule.scala 50:27]
  wire [4:0] cacheLookup_toResponse_request_branch_mask; // @[cacheModule.scala 50:27]
  wire [63:0] cacheLookup_toResponse_request_writeData_data; // @[cacheModule.scala 50:27]
  wire  cacheLookup_writeInstructionCommit_ready; // @[cacheModule.scala 50:27]
  wire  cacheLookup_writeInstructionCommit_fired; // @[cacheModule.scala 50:27]
  wire  cacheLookup_branchOps_valid; // @[cacheModule.scala 50:27]
  wire [4:0] cacheLookup_branchOps_branchMask; // @[cacheModule.scala 50:27]
  wire  cacheLookup_branchOps_passed; // @[cacheModule.scala 50:27]
  wire  replayUnit_clock; // @[cacheModule.scala 51:26]
  wire  replayUnit_reset; // @[cacheModule.scala 51:26]
  wire  replayUnit_requestIn_ready; // @[cacheModule.scala 51:26]
  wire  replayUnit_requestIn_request_valid; // @[cacheModule.scala 51:26]
  wire [31:0] replayUnit_requestIn_request_address; // @[cacheModule.scala 51:26]
  wire [31:0] replayUnit_requestIn_request_core_instruction; // @[cacheModule.scala 51:26]
  wire [3:0] replayUnit_requestIn_request_core_robAddr; // @[cacheModule.scala 51:26]
  wire [5:0] replayUnit_requestIn_request_core_prfDest; // @[cacheModule.scala 51:26]
  wire  replayUnit_requestIn_request_branch_valid; // @[cacheModule.scala 51:26]
  wire [4:0] replayUnit_requestIn_request_branch_mask; // @[cacheModule.scala 51:26]
  wire  replayUnit_requestIn_request_writeData_valid; // @[cacheModule.scala 51:26]
  wire [63:0] replayUnit_requestIn_request_writeData_data; // @[cacheModule.scala 51:26]
  wire [1:0] replayUnit_requestIn_request_cacheLine_response; // @[cacheModule.scala 51:26]
  wire  replayUnit_requestOut_ready; // @[cacheModule.scala 51:26]
  wire  replayUnit_requestOut_request_valid; // @[cacheModule.scala 51:26]
  wire [31:0] replayUnit_requestOut_request_address; // @[cacheModule.scala 51:26]
  wire [31:0] replayUnit_requestOut_request_core_instruction; // @[cacheModule.scala 51:26]
  wire [3:0] replayUnit_requestOut_request_core_robAddr; // @[cacheModule.scala 51:26]
  wire [5:0] replayUnit_requestOut_request_core_prfDest; // @[cacheModule.scala 51:26]
  wire  replayUnit_requestOut_request_branch_valid; // @[cacheModule.scala 51:26]
  wire [4:0] replayUnit_requestOut_request_branch_mask; // @[cacheModule.scala 51:26]
  wire  replayUnit_requestOut_request_writeData_valid; // @[cacheModule.scala 51:26]
  wire [63:0] replayUnit_requestOut_request_writeData_data; // @[cacheModule.scala 51:26]
  wire [1:0] replayUnit_requestOut_request_cacheLine_response; // @[cacheModule.scala 51:26]
  wire  replayUnit_responseIn_ready; // @[cacheModule.scala 51:26]
  wire  replayUnit_responseIn_request_valid; // @[cacheModule.scala 51:26]
  wire [31:0] replayUnit_responseIn_request_address; // @[cacheModule.scala 51:26]
  wire [31:0] replayUnit_responseIn_request_core_instruction; // @[cacheModule.scala 51:26]
  wire [3:0] replayUnit_responseIn_request_core_robAddr; // @[cacheModule.scala 51:26]
  wire [5:0] replayUnit_responseIn_request_core_prfDest; // @[cacheModule.scala 51:26]
  wire  replayUnit_responseIn_request_branch_valid; // @[cacheModule.scala 51:26]
  wire [4:0] replayUnit_responseIn_request_branch_mask; // @[cacheModule.scala 51:26]
  wire  replayUnit_responseIn_request_writeData_valid; // @[cacheModule.scala 51:26]
  wire [63:0] replayUnit_responseIn_request_writeData_data; // @[cacheModule.scala 51:26]
  wire [511:0] replayUnit_responseIn_request_cacheLine_cacheLine; // @[cacheModule.scala 51:26]
  wire [1:0] replayUnit_responseIn_request_cacheLine_response; // @[cacheModule.scala 51:26]
  wire  replayUnit_responseOut_ready; // @[cacheModule.scala 51:26]
  wire  replayUnit_responseOut_request_valid; // @[cacheModule.scala 51:26]
  wire [31:0] replayUnit_responseOut_request_address; // @[cacheModule.scala 51:26]
  wire [31:0] replayUnit_responseOut_request_core_instruction; // @[cacheModule.scala 51:26]
  wire [3:0] replayUnit_responseOut_request_core_robAddr; // @[cacheModule.scala 51:26]
  wire [5:0] replayUnit_responseOut_request_core_prfDest; // @[cacheModule.scala 51:26]
  wire  replayUnit_responseOut_request_branch_valid; // @[cacheModule.scala 51:26]
  wire [4:0] replayUnit_responseOut_request_branch_mask; // @[cacheModule.scala 51:26]
  wire  replayUnit_responseOut_request_writeData_valid; // @[cacheModule.scala 51:26]
  wire [63:0] replayUnit_responseOut_request_writeData_data; // @[cacheModule.scala 51:26]
  wire [511:0] replayUnit_responseOut_request_cacheLine_cacheLine; // @[cacheModule.scala 51:26]
  wire [1:0] replayUnit_responseOut_request_cacheLine_response; // @[cacheModule.scala 51:26]
  wire  replayUnit_writeBackIn_ready; // @[cacheModule.scala 51:26]
  wire  replayUnit_writeBackIn_request_valid; // @[cacheModule.scala 51:26]
  wire [31:0] replayUnit_writeBackIn_request_address; // @[cacheModule.scala 51:26]
  wire [511:0] replayUnit_writeBackIn_request_data; // @[cacheModule.scala 51:26]
  wire  replayUnit_writeBackOut_ready; // @[cacheModule.scala 51:26]
  wire  replayUnit_writeBackOut_request_valid; // @[cacheModule.scala 51:26]
  wire [31:0] replayUnit_writeBackOut_request_address; // @[cacheModule.scala 51:26]
  wire [511:0] replayUnit_writeBackOut_request_data; // @[cacheModule.scala 51:26]
  wire  replayUnit_branchOps_valid; // @[cacheModule.scala 51:26]
  wire [4:0] replayUnit_branchOps_branchMask; // @[cacheModule.scala 51:26]
  wire  replayUnit_branchOps_passed; // @[cacheModule.scala 51:26]
  wire  replayUnit_fenceReady; // @[cacheModule.scala 51:26]
  wire  peripheralUnit_clock; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_reset; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_request_ready; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_request_request_valid; // @[cacheModule.scala 52:30]
  wire [31:0] peripheralUnit_request_request_address; // @[cacheModule.scala 52:30]
  wire [31:0] peripheralUnit_request_request_core_instruction; // @[cacheModule.scala 52:30]
  wire [3:0] peripheralUnit_request_request_core_robAddr; // @[cacheModule.scala 52:30]
  wire [5:0] peripheralUnit_request_request_core_prfDest; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_request_request_branch_valid; // @[cacheModule.scala 52:30]
  wire [4:0] peripheralUnit_request_request_branch_mask; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_request_request_writeData_valid; // @[cacheModule.scala 52:30]
  wire [63:0] peripheralUnit_request_request_writeData_data; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_responseOut_ready; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_responseOut_request_valid; // @[cacheModule.scala 52:30]
  wire [31:0] peripheralUnit_responseOut_request_address; // @[cacheModule.scala 52:30]
  wire [31:0] peripheralUnit_responseOut_request_core_instruction; // @[cacheModule.scala 52:30]
  wire [3:0] peripheralUnit_responseOut_request_core_robAddr; // @[cacheModule.scala 52:30]
  wire [5:0] peripheralUnit_responseOut_request_core_prfDest; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_responseOut_request_branch_valid; // @[cacheModule.scala 52:30]
  wire [4:0] peripheralUnit_responseOut_request_branch_mask; // @[cacheModule.scala 52:30]
  wire [63:0] peripheralUnit_responseOut_request_writeData_data; // @[cacheModule.scala 52:30]
  wire [31:0] peripheralUnit_bus_AWADDR; // @[cacheModule.scala 52:30]
  wire [7:0] peripheralUnit_bus_AWLEN; // @[cacheModule.scala 52:30]
  wire [2:0] peripheralUnit_bus_AWSIZE; // @[cacheModule.scala 52:30]
  wire [1:0] peripheralUnit_bus_AWBURST; // @[cacheModule.scala 52:30]
  wire [2:0] peripheralUnit_bus_AWPROT; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_bus_AWVALID; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_bus_AWREADY; // @[cacheModule.scala 52:30]
  wire [31:0] peripheralUnit_bus_WDATA; // @[cacheModule.scala 52:30]
  wire [3:0] peripheralUnit_bus_WSTRB; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_bus_WLAST; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_bus_WVALID; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_bus_WREADY; // @[cacheModule.scala 52:30]
  wire [1:0] peripheralUnit_bus_BID; // @[cacheModule.scala 52:30]
  wire [1:0] peripheralUnit_bus_BRESP; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_bus_BVALID; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_bus_BREADY; // @[cacheModule.scala 52:30]
  wire [31:0] peripheralUnit_bus_ARADDR; // @[cacheModule.scala 52:30]
  wire [7:0] peripheralUnit_bus_ARLEN; // @[cacheModule.scala 52:30]
  wire [2:0] peripheralUnit_bus_ARSIZE; // @[cacheModule.scala 52:30]
  wire [1:0] peripheralUnit_bus_ARBURST; // @[cacheModule.scala 52:30]
  wire [2:0] peripheralUnit_bus_ARPROT; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_bus_ARVALID; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_bus_ARREADY; // @[cacheModule.scala 52:30]
  wire [1:0] peripheralUnit_bus_RID; // @[cacheModule.scala 52:30]
  wire [31:0] peripheralUnit_bus_RDATA; // @[cacheModule.scala 52:30]
  wire [1:0] peripheralUnit_bus_RRESP; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_bus_RLAST; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_bus_RVALID; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_bus_RREADY; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_writeInstructionCommit_ready; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_writeInstructionCommit_fired; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_branchOps_valid; // @[cacheModule.scala 52:30]
  wire [4:0] peripheralUnit_branchOps_branchMask; // @[cacheModule.scala 52:30]
  wire  peripheralUnit_branchOps_passed; // @[cacheModule.scala 52:30]
  wire  aceUnit_clock; // @[cacheModule.scala 59:23]
  wire  aceUnit_reset; // @[cacheModule.scala 59:23]
  wire  aceUnit_readRequest_ready; // @[cacheModule.scala 59:23]
  wire  aceUnit_readRequest_request_valid; // @[cacheModule.scala 59:23]
  wire [31:0] aceUnit_readRequest_request_address; // @[cacheModule.scala 59:23]
  wire [31:0] aceUnit_readRequest_request_core_instruction; // @[cacheModule.scala 59:23]
  wire [3:0] aceUnit_readRequest_request_core_robAddr; // @[cacheModule.scala 59:23]
  wire [5:0] aceUnit_readRequest_request_core_prfDest; // @[cacheModule.scala 59:23]
  wire  aceUnit_readRequest_request_branch_valid; // @[cacheModule.scala 59:23]
  wire [4:0] aceUnit_readRequest_request_branch_mask; // @[cacheModule.scala 59:23]
  wire  aceUnit_readRequest_request_writeData_valid; // @[cacheModule.scala 59:23]
  wire [63:0] aceUnit_readRequest_request_writeData_data; // @[cacheModule.scala 59:23]
  wire [1:0] aceUnit_readRequest_request_cacheLine_response; // @[cacheModule.scala 59:23]
  wire  aceUnit_readResponse_ready; // @[cacheModule.scala 59:23]
  wire  aceUnit_readResponse_request_valid; // @[cacheModule.scala 59:23]
  wire [31:0] aceUnit_readResponse_request_address; // @[cacheModule.scala 59:23]
  wire [31:0] aceUnit_readResponse_request_core_instruction; // @[cacheModule.scala 59:23]
  wire [3:0] aceUnit_readResponse_request_core_robAddr; // @[cacheModule.scala 59:23]
  wire [5:0] aceUnit_readResponse_request_core_prfDest; // @[cacheModule.scala 59:23]
  wire  aceUnit_readResponse_request_branch_valid; // @[cacheModule.scala 59:23]
  wire [4:0] aceUnit_readResponse_request_branch_mask; // @[cacheModule.scala 59:23]
  wire  aceUnit_readResponse_request_writeData_valid; // @[cacheModule.scala 59:23]
  wire [63:0] aceUnit_readResponse_request_writeData_data; // @[cacheModule.scala 59:23]
  wire [511:0] aceUnit_readResponse_request_cacheLine_cacheLine; // @[cacheModule.scala 59:23]
  wire [1:0] aceUnit_readResponse_request_cacheLine_response; // @[cacheModule.scala 59:23]
  wire  aceUnit_writeRequest_ready; // @[cacheModule.scala 59:23]
  wire  aceUnit_writeRequest_request_valid; // @[cacheModule.scala 59:23]
  wire [31:0] aceUnit_writeRequest_request_address; // @[cacheModule.scala 59:23]
  wire [511:0] aceUnit_writeRequest_request_data; // @[cacheModule.scala 59:23]
  wire  aceUnit_coherencyRequest_ready; // @[cacheModule.scala 59:23]
  wire  aceUnit_coherencyRequest_request_valid; // @[cacheModule.scala 59:23]
  wire [31:0] aceUnit_coherencyRequest_request_address; // @[cacheModule.scala 59:23]
  wire [1:0] aceUnit_coherencyRequest_request_response; // @[cacheModule.scala 59:23]
  wire  aceUnit_coherencyResponse_ready; // @[cacheModule.scala 59:23]
  wire  aceUnit_coherencyResponse_request_valid; // @[cacheModule.scala 59:23]
  wire [1:0] aceUnit_coherencyResponse_request_response; // @[cacheModule.scala 59:23]
  wire [511:0] aceUnit_coherencyResponse_request_cacheLine; // @[cacheModule.scala 59:23]
  wire  aceUnit_coherencyResponse_request_dataValid; // @[cacheModule.scala 59:23]
  wire  aceUnit_fenceReady; // @[cacheModule.scala 59:23]
  wire  aceUnit_branchOps_valid; // @[cacheModule.scala 59:23]
  wire [4:0] aceUnit_branchOps_branchMask; // @[cacheModule.scala 59:23]
  wire  aceUnit_branchOps_passed; // @[cacheModule.scala 59:23]
  wire [31:0] aceUnit_bus_AWADDR; // @[cacheModule.scala 59:23]
  wire  aceUnit_bus_AWVALID; // @[cacheModule.scala 59:23]
  wire  aceUnit_bus_AWREADY; // @[cacheModule.scala 59:23]
  wire [63:0] aceUnit_bus_WDATA; // @[cacheModule.scala 59:23]
  wire  aceUnit_bus_WLAST; // @[cacheModule.scala 59:23]
  wire  aceUnit_bus_WVALID; // @[cacheModule.scala 59:23]
  wire  aceUnit_bus_WREADY; // @[cacheModule.scala 59:23]
  wire [1:0] aceUnit_bus_BRESP; // @[cacheModule.scala 59:23]
  wire  aceUnit_bus_BVALID; // @[cacheModule.scala 59:23]
  wire  aceUnit_bus_BREADY; // @[cacheModule.scala 59:23]
  wire [31:0] aceUnit_bus_ARADDR; // @[cacheModule.scala 59:23]
  wire  aceUnit_bus_ARVALID; // @[cacheModule.scala 59:23]
  wire  aceUnit_bus_ARREADY; // @[cacheModule.scala 59:23]
  wire [63:0] aceUnit_bus_RDATA; // @[cacheModule.scala 59:23]
  wire  aceUnit_bus_RLAST; // @[cacheModule.scala 59:23]
  wire  aceUnit_bus_RVALID; // @[cacheModule.scala 59:23]
  wire  aceUnit_bus_RREADY; // @[cacheModule.scala 59:23]
  wire [2:0] aceUnit_bus_AWSNOOP; // @[cacheModule.scala 59:23]
  wire [3:0] aceUnit_bus_ARSNOOP; // @[cacheModule.scala 59:23]
  wire [3:0] aceUnit_bus_RRESP; // @[cacheModule.scala 59:23]
  wire  aceUnit_bus_ACVALID; // @[cacheModule.scala 59:23]
  wire  aceUnit_bus_ACREADY; // @[cacheModule.scala 59:23]
  wire [31:0] aceUnit_bus_ACADDR; // @[cacheModule.scala 59:23]
  wire [3:0] aceUnit_bus_ACSNOOP; // @[cacheModule.scala 59:23]
  wire  aceUnit_bus_CRVALID; // @[cacheModule.scala 59:23]
  wire  aceUnit_bus_CRREADY; // @[cacheModule.scala 59:23]
  wire [4:0] aceUnit_bus_CRRESP; // @[cacheModule.scala 59:23]
  wire  aceUnit_bus_CDVALID; // @[cacheModule.scala 59:23]
  wire  aceUnit_bus_CDREADY; // @[cacheModule.scala 59:23]
  wire [63:0] aceUnit_bus_CDDATA; // @[cacheModule.scala 59:23]
  wire  aceUnit_bus_CDLAST; // @[cacheModule.scala 59:23]
  wire  commitFifo_clock; // @[cacheModule.scala 66:26]
  wire  commitFifo_reset; // @[cacheModule.scala 66:26]
  wire  commitFifo_write_data_valid; // @[cacheModule.scala 66:26]
  wire [31:0] commitFifo_write_data_address; // @[cacheModule.scala 66:26]
  wire  commitFifo_write_data_branch_valid; // @[cacheModule.scala 66:26]
  wire [4:0] commitFifo_write_data_branch_mask; // @[cacheModule.scala 66:26]
  wire  commitFifo_read_ready; // @[cacheModule.scala 66:26]
  wire  commitFifo_read_data_valid; // @[cacheModule.scala 66:26]
  wire  commitFifo_read_data_branch_valid; // @[cacheModule.scala 66:26]
  wire  commitFifo_isEmpty; // @[cacheModule.scala 66:26]
  wire  commitFifo_branchOps_valid; // @[cacheModule.scala 66:26]
  wire [4:0] commitFifo_branchOps_branchMask; // @[cacheModule.scala 66:26]
  wire  commitFifo_branchOps_passed; // @[cacheModule.scala 66:26]
  wire  commitFifo_isFull; // @[cacheModule.scala 66:26]
  wire [31:0] commitFifo_invalidateAddr; // @[cacheModule.scala 66:26]
  wire  commitFifo_invalidateEnable; // @[cacheModule.scala 66:26]
  wire  _responseOut_valid_T = cacheLookup_toResponse_request_valid & cacheLookup_toResponse_request_branch_valid; // @[cacheModule.scala 139:103]
  wire [4:0] _GEN_8 = peripheralUnit_responseOut_request_valid ? peripheralUnit_responseOut_request_branch_mask : 5'h0; // @[cacheModule.scala 161:56 162:27 utils.scala 49:41]
  wire  _GEN_9 = peripheralUnit_responseOut_request_valid & peripheralUnit_responseOut_request_branch_valid; // @[cacheModule.scala 161:56 162:27 utils.scala 48:41]
  wire [31:0] _GEN_13 = peripheralUnit_responseOut_request_valid ? peripheralUnit_responseOut_request_address : 32'h0; // @[cacheModule.scala 161:56 162:27 utils.scala 49:41]
  wire  _GEN_14 = peripheralUnit_responseOut_request_valid; // @[cacheModule.scala 161:56 162:27 utils.scala 48:41]
  wire  _GEN_29 = commitFifo_isEmpty ? 1'h0 : commitFifo_read_data_valid; // @[cacheModule.scala 174:22 176:29 177:24]
  wire  _GEN_30 = commitFifo_isEmpty | ~commitFifo_isEmpty & commitFifo_read_data_branch_valid; // @[cacheModule.scala 175:22 176:29 178:24]
  reg  fenceInititatedReg; // @[cacheModule.scala 183:35]
  reg  canInititatedFenceReg; // @[cacheModule.scala 184:38]
  wire  _subModulesReady_T = requestScheduler_fenceReady & arbiter_fenceReady; // @[cacheModule.scala 186:33]
  wire  _subModulesReady_T_1 = _subModulesReady_T & replayUnit_fenceReady; // @[cacheModule.scala 187:24]
  wire  _subModulesReady_T_2 = _subModulesReady_T_1 & aceUnit_fenceReady; // @[cacheModule.scala 188:27]
  reg  subModulesReady_REG; // @[cacheModule.scala 190:20]
  reg  subModulesReady_REG_1; // @[cacheModule.scala 190:12]
  wire  subModulesReady = _subModulesReady_T_2 & subModulesReady_REG_1; // @[cacheModule.scala 189:24]
  requestScheduler requestScheduler ( // @[cacheModule.scala 48:32]
    .clock(requestScheduler_clock),
    .reset(requestScheduler_reset),
    .requestIn_valid(requestScheduler_requestIn_valid),
    .requestIn_address(requestScheduler_requestIn_address),
    .requestIn_core_instruction(requestScheduler_requestIn_core_instruction),
    .requestIn_core_robAddr(requestScheduler_requestIn_core_robAddr),
    .requestIn_core_prfDest(requestScheduler_requestIn_core_prfDest),
    .requestIn_branch_mask(requestScheduler_requestIn_branch_mask),
    .canAllocate(requestScheduler_canAllocate),
    .requestOut_valid(requestScheduler_requestOut_valid),
    .requestOut_address(requestScheduler_requestOut_address),
    .requestOut_core_instruction(requestScheduler_requestOut_core_instruction),
    .requestOut_core_robAddr(requestScheduler_requestOut_core_robAddr),
    .requestOut_core_prfDest(requestScheduler_requestOut_core_prfDest),
    .requestOut_branch_valid(requestScheduler_requestOut_branch_valid),
    .requestOut_branch_mask(requestScheduler_requestOut_branch_mask),
    .requestOut_writeData_valid(requestScheduler_requestOut_writeData_valid),
    .requestOut_writeData_data(requestScheduler_requestOut_writeData_data),
    .controlSignal_isSpeculative(requestScheduler_controlSignal_isSpeculative),
    .controlSignal_inorderReady(requestScheduler_controlSignal_inorderReady),
    .controlSignal_speculativeReady(requestScheduler_controlSignal_speculativeReady),
    .fenceReady(requestScheduler_fenceReady),
    .branchOps_valid(requestScheduler_branchOps_valid),
    .branchOps_branchMask(requestScheduler_branchOps_branchMask),
    .branchOps_passed(requestScheduler_branchOps_passed)
  );
  arbiter arbiter ( // @[cacheModule.scala 49:23]
    .clock(arbiter_clock),
    .reset(arbiter_reset),
    .request_request_valid(arbiter_request_request_valid),
    .request_request_address(arbiter_request_request_address),
    .request_request_core_instruction(arbiter_request_request_core_instruction),
    .request_request_core_robAddr(arbiter_request_request_core_robAddr),
    .request_request_core_prfDest(arbiter_request_request_core_prfDest),
    .request_request_branch_valid(arbiter_request_request_branch_valid),
    .request_request_branch_mask(arbiter_request_request_branch_mask),
    .request_request_writeData_valid(arbiter_request_request_writeData_valid),
    .request_request_writeData_data(arbiter_request_request_writeData_data),
    .request_isSpeculative(arbiter_request_isSpeculative),
    .request_inorderReady(arbiter_request_inorderReady),
    .request_speculativeReady(arbiter_request_speculativeReady),
    .toPeripheral_ready(arbiter_toPeripheral_ready),
    .toPeripheral_request_valid(arbiter_toPeripheral_request_valid),
    .toPeripheral_request_address(arbiter_toPeripheral_request_address),
    .toPeripheral_request_core_instruction(arbiter_toPeripheral_request_core_instruction),
    .toPeripheral_request_core_robAddr(arbiter_toPeripheral_request_core_robAddr),
    .toPeripheral_request_core_prfDest(arbiter_toPeripheral_request_core_prfDest),
    .toPeripheral_request_branch_valid(arbiter_toPeripheral_request_branch_valid),
    .toPeripheral_request_branch_mask(arbiter_toPeripheral_request_branch_mask),
    .toPeripheral_request_writeData_valid(arbiter_toPeripheral_request_writeData_valid),
    .toPeripheral_request_writeData_data(arbiter_toPeripheral_request_writeData_data),
    .toCacheLookup_ready(arbiter_toCacheLookup_ready),
    .toCacheLookup_holdInOrder(arbiter_toCacheLookup_holdInOrder),
    .toCacheLookup_requestType(arbiter_toCacheLookup_requestType),
    .toCacheLookup_request_valid(arbiter_toCacheLookup_request_valid),
    .toCacheLookup_request_address(arbiter_toCacheLookup_request_address),
    .toCacheLookup_request_core_instruction(arbiter_toCacheLookup_request_core_instruction),
    .toCacheLookup_request_core_robAddr(arbiter_toCacheLookup_request_core_robAddr),
    .toCacheLookup_request_core_prfDest(arbiter_toCacheLookup_request_core_prfDest),
    .toCacheLookup_request_branch_valid(arbiter_toCacheLookup_request_branch_valid),
    .toCacheLookup_request_branch_mask(arbiter_toCacheLookup_request_branch_mask),
    .toCacheLookup_request_writeData_valid(arbiter_toCacheLookup_request_writeData_valid),
    .toCacheLookup_request_writeData_data(arbiter_toCacheLookup_request_writeData_data),
    .toCacheLookup_request_cacheLine_cacheLine(arbiter_toCacheLookup_request_cacheLine_cacheLine),
    .toCacheLookup_request_cacheLine_response(arbiter_toCacheLookup_request_cacheLine_response),
    .replayRequest_ready(arbiter_replayRequest_ready),
    .replayRequest_request_valid(arbiter_replayRequest_request_valid),
    .replayRequest_request_address(arbiter_replayRequest_request_address),
    .replayRequest_request_core_instruction(arbiter_replayRequest_request_core_instruction),
    .replayRequest_request_core_robAddr(arbiter_replayRequest_request_core_robAddr),
    .replayRequest_request_core_prfDest(arbiter_replayRequest_request_core_prfDest),
    .replayRequest_request_branch_valid(arbiter_replayRequest_request_branch_valid),
    .replayRequest_request_branch_mask(arbiter_replayRequest_request_branch_mask),
    .replayRequest_request_writeData_valid(arbiter_replayRequest_request_writeData_valid),
    .replayRequest_request_writeData_data(arbiter_replayRequest_request_writeData_data),
    .replayRequest_request_cacheLine_cacheLine(arbiter_replayRequest_request_cacheLine_cacheLine),
    .replayRequest_request_cacheLine_response(arbiter_replayRequest_request_cacheLine_response),
    .coherencyRequest_ready(arbiter_coherencyRequest_ready),
    .coherencyRequest_request_valid(arbiter_coherencyRequest_request_valid),
    .coherencyRequest_request_address(arbiter_coherencyRequest_request_address),
    .coherencyRequest_request_response(arbiter_coherencyRequest_request_response),
    .writeDataIn_valid(arbiter_writeDataIn_valid),
    .writeDataIn_data(arbiter_writeDataIn_data),
    .writeCommit_ready(arbiter_writeCommit_ready),
    .writeCommit_fired(arbiter_writeCommit_fired),
    .branchOps_valid(arbiter_branchOps_valid),
    .branchOps_branchMask(arbiter_branchOps_branchMask),
    .branchOps_passed(arbiter_branchOps_passed),
    .responseOut_valid(arbiter_responseOut_valid),
    .responseOut_instruction(arbiter_responseOut_instruction),
    .fenceReady(arbiter_fenceReady),
    .writeInstuctionCommitFired(arbiter_writeInstuctionCommitFired)
  );
  cacheLookupUnit cacheLookup ( // @[cacheModule.scala 50:27]
    .clock(cacheLookup_clock),
    .reset(cacheLookup_reset),
    .request_ready(cacheLookup_request_ready),
    .request_holdInOrder(cacheLookup_request_holdInOrder),
    .request_requestType(cacheLookup_request_requestType),
    .request_request_valid(cacheLookup_request_request_valid),
    .request_request_address(cacheLookup_request_request_address),
    .request_request_core_instruction(cacheLookup_request_request_core_instruction),
    .request_request_core_robAddr(cacheLookup_request_request_core_robAddr),
    .request_request_core_prfDest(cacheLookup_request_request_core_prfDest),
    .request_request_branch_valid(cacheLookup_request_request_branch_valid),
    .request_request_branch_mask(cacheLookup_request_request_branch_mask),
    .request_request_writeData_valid(cacheLookup_request_request_writeData_valid),
    .request_request_writeData_data(cacheLookup_request_request_writeData_data),
    .request_request_cacheLine_cacheLine(cacheLookup_request_request_cacheLine_cacheLine),
    .request_request_cacheLine_response(cacheLookup_request_request_cacheLine_response),
    .toReplay_ready(cacheLookup_toReplay_ready),
    .toReplay_request_valid(cacheLookup_toReplay_request_valid),
    .toReplay_request_address(cacheLookup_toReplay_request_address),
    .toReplay_request_core_instruction(cacheLookup_toReplay_request_core_instruction),
    .toReplay_request_core_robAddr(cacheLookup_toReplay_request_core_robAddr),
    .toReplay_request_core_prfDest(cacheLookup_toReplay_request_core_prfDest),
    .toReplay_request_branch_valid(cacheLookup_toReplay_request_branch_valid),
    .toReplay_request_branch_mask(cacheLookup_toReplay_request_branch_mask),
    .toReplay_request_writeData_valid(cacheLookup_toReplay_request_writeData_valid),
    .toReplay_request_writeData_data(cacheLookup_toReplay_request_writeData_data),
    .toReplay_request_cacheLine_response(cacheLookup_toReplay_request_cacheLine_response),
    .toWriteBack_ready(cacheLookup_toWriteBack_ready),
    .toWriteBack_request_valid(cacheLookup_toWriteBack_request_valid),
    .toWriteBack_request_address(cacheLookup_toWriteBack_request_address),
    .toWriteBack_request_data(cacheLookup_toWriteBack_request_data),
    .toCoherency_ready(cacheLookup_toCoherency_ready),
    .toCoherency_request_valid(cacheLookup_toCoherency_request_valid),
    .toCoherency_request_response(cacheLookup_toCoherency_request_response),
    .toCoherency_request_cacheLine(cacheLookup_toCoherency_request_cacheLine),
    .toCoherency_request_dataValid(cacheLookup_toCoherency_request_dataValid),
    .toResponse_request_valid(cacheLookup_toResponse_request_valid),
    .toResponse_request_address(cacheLookup_toResponse_request_address),
    .toResponse_request_core_instruction(cacheLookup_toResponse_request_core_instruction),
    .toResponse_request_core_robAddr(cacheLookup_toResponse_request_core_robAddr),
    .toResponse_request_core_prfDest(cacheLookup_toResponse_request_core_prfDest),
    .toResponse_request_branch_valid(cacheLookup_toResponse_request_branch_valid),
    .toResponse_request_branch_mask(cacheLookup_toResponse_request_branch_mask),
    .toResponse_request_writeData_data(cacheLookup_toResponse_request_writeData_data),
    .writeInstructionCommit_ready(cacheLookup_writeInstructionCommit_ready),
    .writeInstructionCommit_fired(cacheLookup_writeInstructionCommit_fired),
    .branchOps_valid(cacheLookup_branchOps_valid),
    .branchOps_branchMask(cacheLookup_branchOps_branchMask),
    .branchOps_passed(cacheLookup_branchOps_passed)
  );
  replayUnit replayUnit ( // @[cacheModule.scala 51:26]
    .clock(replayUnit_clock),
    .reset(replayUnit_reset),
    .requestIn_ready(replayUnit_requestIn_ready),
    .requestIn_request_valid(replayUnit_requestIn_request_valid),
    .requestIn_request_address(replayUnit_requestIn_request_address),
    .requestIn_request_core_instruction(replayUnit_requestIn_request_core_instruction),
    .requestIn_request_core_robAddr(replayUnit_requestIn_request_core_robAddr),
    .requestIn_request_core_prfDest(replayUnit_requestIn_request_core_prfDest),
    .requestIn_request_branch_valid(replayUnit_requestIn_request_branch_valid),
    .requestIn_request_branch_mask(replayUnit_requestIn_request_branch_mask),
    .requestIn_request_writeData_valid(replayUnit_requestIn_request_writeData_valid),
    .requestIn_request_writeData_data(replayUnit_requestIn_request_writeData_data),
    .requestIn_request_cacheLine_response(replayUnit_requestIn_request_cacheLine_response),
    .requestOut_ready(replayUnit_requestOut_ready),
    .requestOut_request_valid(replayUnit_requestOut_request_valid),
    .requestOut_request_address(replayUnit_requestOut_request_address),
    .requestOut_request_core_instruction(replayUnit_requestOut_request_core_instruction),
    .requestOut_request_core_robAddr(replayUnit_requestOut_request_core_robAddr),
    .requestOut_request_core_prfDest(replayUnit_requestOut_request_core_prfDest),
    .requestOut_request_branch_valid(replayUnit_requestOut_request_branch_valid),
    .requestOut_request_branch_mask(replayUnit_requestOut_request_branch_mask),
    .requestOut_request_writeData_valid(replayUnit_requestOut_request_writeData_valid),
    .requestOut_request_writeData_data(replayUnit_requestOut_request_writeData_data),
    .requestOut_request_cacheLine_response(replayUnit_requestOut_request_cacheLine_response),
    .responseIn_ready(replayUnit_responseIn_ready),
    .responseIn_request_valid(replayUnit_responseIn_request_valid),
    .responseIn_request_address(replayUnit_responseIn_request_address),
    .responseIn_request_core_instruction(replayUnit_responseIn_request_core_instruction),
    .responseIn_request_core_robAddr(replayUnit_responseIn_request_core_robAddr),
    .responseIn_request_core_prfDest(replayUnit_responseIn_request_core_prfDest),
    .responseIn_request_branch_valid(replayUnit_responseIn_request_branch_valid),
    .responseIn_request_branch_mask(replayUnit_responseIn_request_branch_mask),
    .responseIn_request_writeData_valid(replayUnit_responseIn_request_writeData_valid),
    .responseIn_request_writeData_data(replayUnit_responseIn_request_writeData_data),
    .responseIn_request_cacheLine_cacheLine(replayUnit_responseIn_request_cacheLine_cacheLine),
    .responseIn_request_cacheLine_response(replayUnit_responseIn_request_cacheLine_response),
    .responseOut_ready(replayUnit_responseOut_ready),
    .responseOut_request_valid(replayUnit_responseOut_request_valid),
    .responseOut_request_address(replayUnit_responseOut_request_address),
    .responseOut_request_core_instruction(replayUnit_responseOut_request_core_instruction),
    .responseOut_request_core_robAddr(replayUnit_responseOut_request_core_robAddr),
    .responseOut_request_core_prfDest(replayUnit_responseOut_request_core_prfDest),
    .responseOut_request_branch_valid(replayUnit_responseOut_request_branch_valid),
    .responseOut_request_branch_mask(replayUnit_responseOut_request_branch_mask),
    .responseOut_request_writeData_valid(replayUnit_responseOut_request_writeData_valid),
    .responseOut_request_writeData_data(replayUnit_responseOut_request_writeData_data),
    .responseOut_request_cacheLine_cacheLine(replayUnit_responseOut_request_cacheLine_cacheLine),
    .responseOut_request_cacheLine_response(replayUnit_responseOut_request_cacheLine_response),
    .writeBackIn_ready(replayUnit_writeBackIn_ready),
    .writeBackIn_request_valid(replayUnit_writeBackIn_request_valid),
    .writeBackIn_request_address(replayUnit_writeBackIn_request_address),
    .writeBackIn_request_data(replayUnit_writeBackIn_request_data),
    .writeBackOut_ready(replayUnit_writeBackOut_ready),
    .writeBackOut_request_valid(replayUnit_writeBackOut_request_valid),
    .writeBackOut_request_address(replayUnit_writeBackOut_request_address),
    .writeBackOut_request_data(replayUnit_writeBackOut_request_data),
    .branchOps_valid(replayUnit_branchOps_valid),
    .branchOps_branchMask(replayUnit_branchOps_branchMask),
    .branchOps_passed(replayUnit_branchOps_passed),
    .fenceReady(replayUnit_fenceReady)
  );
  peripheralUnit peripheralUnit ( // @[cacheModule.scala 52:30]
    .clock(peripheralUnit_clock),
    .reset(peripheralUnit_reset),
    .request_ready(peripheralUnit_request_ready),
    .request_request_valid(peripheralUnit_request_request_valid),
    .request_request_address(peripheralUnit_request_request_address),
    .request_request_core_instruction(peripheralUnit_request_request_core_instruction),
    .request_request_core_robAddr(peripheralUnit_request_request_core_robAddr),
    .request_request_core_prfDest(peripheralUnit_request_request_core_prfDest),
    .request_request_branch_valid(peripheralUnit_request_request_branch_valid),
    .request_request_branch_mask(peripheralUnit_request_request_branch_mask),
    .request_request_writeData_valid(peripheralUnit_request_request_writeData_valid),
    .request_request_writeData_data(peripheralUnit_request_request_writeData_data),
    .responseOut_ready(peripheralUnit_responseOut_ready),
    .responseOut_request_valid(peripheralUnit_responseOut_request_valid),
    .responseOut_request_address(peripheralUnit_responseOut_request_address),
    .responseOut_request_core_instruction(peripheralUnit_responseOut_request_core_instruction),
    .responseOut_request_core_robAddr(peripheralUnit_responseOut_request_core_robAddr),
    .responseOut_request_core_prfDest(peripheralUnit_responseOut_request_core_prfDest),
    .responseOut_request_branch_valid(peripheralUnit_responseOut_request_branch_valid),
    .responseOut_request_branch_mask(peripheralUnit_responseOut_request_branch_mask),
    .responseOut_request_writeData_data(peripheralUnit_responseOut_request_writeData_data),
    .bus_AWADDR(peripheralUnit_bus_AWADDR),
    .bus_AWLEN(peripheralUnit_bus_AWLEN),
    .bus_AWSIZE(peripheralUnit_bus_AWSIZE),
    .bus_AWBURST(peripheralUnit_bus_AWBURST),
    .bus_AWPROT(peripheralUnit_bus_AWPROT),
    .bus_AWVALID(peripheralUnit_bus_AWVALID),
    .bus_AWREADY(peripheralUnit_bus_AWREADY),
    .bus_WDATA(peripheralUnit_bus_WDATA),
    .bus_WSTRB(peripheralUnit_bus_WSTRB),
    .bus_WLAST(peripheralUnit_bus_WLAST),
    .bus_WVALID(peripheralUnit_bus_WVALID),
    .bus_WREADY(peripheralUnit_bus_WREADY),
    .bus_BID(peripheralUnit_bus_BID),
    .bus_BRESP(peripheralUnit_bus_BRESP),
    .bus_BVALID(peripheralUnit_bus_BVALID),
    .bus_BREADY(peripheralUnit_bus_BREADY),
    .bus_ARADDR(peripheralUnit_bus_ARADDR),
    .bus_ARLEN(peripheralUnit_bus_ARLEN),
    .bus_ARSIZE(peripheralUnit_bus_ARSIZE),
    .bus_ARBURST(peripheralUnit_bus_ARBURST),
    .bus_ARPROT(peripheralUnit_bus_ARPROT),
    .bus_ARVALID(peripheralUnit_bus_ARVALID),
    .bus_ARREADY(peripheralUnit_bus_ARREADY),
    .bus_RID(peripheralUnit_bus_RID),
    .bus_RDATA(peripheralUnit_bus_RDATA),
    .bus_RRESP(peripheralUnit_bus_RRESP),
    .bus_RLAST(peripheralUnit_bus_RLAST),
    .bus_RVALID(peripheralUnit_bus_RVALID),
    .bus_RREADY(peripheralUnit_bus_RREADY),
    .writeInstructionCommit_ready(peripheralUnit_writeInstructionCommit_ready),
    .writeInstructionCommit_fired(peripheralUnit_writeInstructionCommit_fired),
    .branchOps_valid(peripheralUnit_branchOps_valid),
    .branchOps_branchMask(peripheralUnit_branchOps_branchMask),
    .branchOps_passed(peripheralUnit_branchOps_passed)
  );
  ACEUnit aceUnit ( // @[cacheModule.scala 59:23]
    .clock(aceUnit_clock),
    .reset(aceUnit_reset),
    .readRequest_ready(aceUnit_readRequest_ready),
    .readRequest_request_valid(aceUnit_readRequest_request_valid),
    .readRequest_request_address(aceUnit_readRequest_request_address),
    .readRequest_request_core_instruction(aceUnit_readRequest_request_core_instruction),
    .readRequest_request_core_robAddr(aceUnit_readRequest_request_core_robAddr),
    .readRequest_request_core_prfDest(aceUnit_readRequest_request_core_prfDest),
    .readRequest_request_branch_valid(aceUnit_readRequest_request_branch_valid),
    .readRequest_request_branch_mask(aceUnit_readRequest_request_branch_mask),
    .readRequest_request_writeData_valid(aceUnit_readRequest_request_writeData_valid),
    .readRequest_request_writeData_data(aceUnit_readRequest_request_writeData_data),
    .readRequest_request_cacheLine_response(aceUnit_readRequest_request_cacheLine_response),
    .readResponse_ready(aceUnit_readResponse_ready),
    .readResponse_request_valid(aceUnit_readResponse_request_valid),
    .readResponse_request_address(aceUnit_readResponse_request_address),
    .readResponse_request_core_instruction(aceUnit_readResponse_request_core_instruction),
    .readResponse_request_core_robAddr(aceUnit_readResponse_request_core_robAddr),
    .readResponse_request_core_prfDest(aceUnit_readResponse_request_core_prfDest),
    .readResponse_request_branch_valid(aceUnit_readResponse_request_branch_valid),
    .readResponse_request_branch_mask(aceUnit_readResponse_request_branch_mask),
    .readResponse_request_writeData_valid(aceUnit_readResponse_request_writeData_valid),
    .readResponse_request_writeData_data(aceUnit_readResponse_request_writeData_data),
    .readResponse_request_cacheLine_cacheLine(aceUnit_readResponse_request_cacheLine_cacheLine),
    .readResponse_request_cacheLine_response(aceUnit_readResponse_request_cacheLine_response),
    .writeRequest_ready(aceUnit_writeRequest_ready),
    .writeRequest_request_valid(aceUnit_writeRequest_request_valid),
    .writeRequest_request_address(aceUnit_writeRequest_request_address),
    .writeRequest_request_data(aceUnit_writeRequest_request_data),
    .coherencyRequest_ready(aceUnit_coherencyRequest_ready),
    .coherencyRequest_request_valid(aceUnit_coherencyRequest_request_valid),
    .coherencyRequest_request_address(aceUnit_coherencyRequest_request_address),
    .coherencyRequest_request_response(aceUnit_coherencyRequest_request_response),
    .coherencyResponse_ready(aceUnit_coherencyResponse_ready),
    .coherencyResponse_request_valid(aceUnit_coherencyResponse_request_valid),
    .coherencyResponse_request_response(aceUnit_coherencyResponse_request_response),
    .coherencyResponse_request_cacheLine(aceUnit_coherencyResponse_request_cacheLine),
    .coherencyResponse_request_dataValid(aceUnit_coherencyResponse_request_dataValid),
    .fenceReady(aceUnit_fenceReady),
    .branchOps_valid(aceUnit_branchOps_valid),
    .branchOps_branchMask(aceUnit_branchOps_branchMask),
    .branchOps_passed(aceUnit_branchOps_passed),
    .bus_AWADDR(aceUnit_bus_AWADDR),
    .bus_AWVALID(aceUnit_bus_AWVALID),
    .bus_AWREADY(aceUnit_bus_AWREADY),
    .bus_WDATA(aceUnit_bus_WDATA),
    .bus_WLAST(aceUnit_bus_WLAST),
    .bus_WVALID(aceUnit_bus_WVALID),
    .bus_WREADY(aceUnit_bus_WREADY),
    .bus_BRESP(aceUnit_bus_BRESP),
    .bus_BVALID(aceUnit_bus_BVALID),
    .bus_BREADY(aceUnit_bus_BREADY),
    .bus_ARADDR(aceUnit_bus_ARADDR),
    .bus_ARVALID(aceUnit_bus_ARVALID),
    .bus_ARREADY(aceUnit_bus_ARREADY),
    .bus_RDATA(aceUnit_bus_RDATA),
    .bus_RLAST(aceUnit_bus_RLAST),
    .bus_RVALID(aceUnit_bus_RVALID),
    .bus_RREADY(aceUnit_bus_RREADY),
    .bus_AWSNOOP(aceUnit_bus_AWSNOOP),
    .bus_ARSNOOP(aceUnit_bus_ARSNOOP),
    .bus_RRESP(aceUnit_bus_RRESP),
    .bus_ACVALID(aceUnit_bus_ACVALID),
    .bus_ACREADY(aceUnit_bus_ACREADY),
    .bus_ACADDR(aceUnit_bus_ACADDR),
    .bus_ACSNOOP(aceUnit_bus_ACSNOOP),
    .bus_CRVALID(aceUnit_bus_CRVALID),
    .bus_CRREADY(aceUnit_bus_CRREADY),
    .bus_CRRESP(aceUnit_bus_CRRESP),
    .bus_CDVALID(aceUnit_bus_CDVALID),
    .bus_CDREADY(aceUnit_bus_CDREADY),
    .bus_CDDATA(aceUnit_bus_CDDATA),
    .bus_CDLAST(aceUnit_bus_CDLAST)
  );
  fifoRecordInvalidateI commitFifo ( // @[cacheModule.scala 66:26]
    .clock(commitFifo_clock),
    .reset(commitFifo_reset),
    .write_data_valid(commitFifo_write_data_valid),
    .write_data_address(commitFifo_write_data_address),
    .write_data_branch_valid(commitFifo_write_data_branch_valid),
    .write_data_branch_mask(commitFifo_write_data_branch_mask),
    .read_ready(commitFifo_read_ready),
    .read_data_valid(commitFifo_read_data_valid),
    .read_data_branch_valid(commitFifo_read_data_branch_valid),
    .isEmpty(commitFifo_isEmpty),
    .branchOps_valid(commitFifo_branchOps_valid),
    .branchOps_branchMask(commitFifo_branchOps_branchMask),
    .branchOps_passed(commitFifo_branchOps_passed),
    .isFull(commitFifo_isFull),
    .invalidateAddr(commitFifo_invalidateAddr),
    .invalidateEnable(commitFifo_invalidateEnable)
  );
  assign dPort_AWADDR = aceUnit_bus_AWADDR; // @[cacheModule.scala 125:15]
  assign dPort_AWVALID = aceUnit_bus_AWVALID; // @[cacheModule.scala 125:15]
  assign dPort_WDATA = aceUnit_bus_WDATA; // @[cacheModule.scala 125:15]
  assign dPort_WLAST = aceUnit_bus_WLAST; // @[cacheModule.scala 125:15]
  assign dPort_WVALID = aceUnit_bus_WVALID; // @[cacheModule.scala 125:15]
  assign dPort_BREADY = aceUnit_bus_BREADY; // @[cacheModule.scala 125:15]
  assign dPort_ARADDR = aceUnit_bus_ARADDR; // @[cacheModule.scala 125:15]
  assign dPort_ARVALID = aceUnit_bus_ARVALID; // @[cacheModule.scala 125:15]
  assign dPort_RREADY = aceUnit_bus_RREADY; // @[cacheModule.scala 125:15]
  assign dPort_AWSNOOP = aceUnit_bus_AWSNOOP; // @[cacheModule.scala 125:15]
  assign dPort_ARSNOOP = aceUnit_bus_ARSNOOP; // @[cacheModule.scala 125:15]
  assign dPort_ACREADY = aceUnit_bus_ACREADY; // @[cacheModule.scala 125:15]
  assign dPort_CRVALID = aceUnit_bus_CRVALID; // @[cacheModule.scala 125:15]
  assign dPort_CRRESP = aceUnit_bus_CRRESP; // @[cacheModule.scala 125:15]
  assign dPort_CDVALID = aceUnit_bus_CDVALID; // @[cacheModule.scala 125:15]
  assign dPort_CDDATA = aceUnit_bus_CDDATA; // @[cacheModule.scala 125:15]
  assign dPort_CDLAST = aceUnit_bus_CDLAST; // @[cacheModule.scala 125:15]
  assign peripheral_AWADDR = peripheralUnit_bus_AWADDR; // @[cacheModule.scala 133:22]
  assign peripheral_AWLEN = peripheralUnit_bus_AWLEN; // @[cacheModule.scala 133:22]
  assign peripheral_AWSIZE = peripheralUnit_bus_AWSIZE; // @[cacheModule.scala 133:22]
  assign peripheral_AWBURST = peripheralUnit_bus_AWBURST; // @[cacheModule.scala 133:22]
  assign peripheral_AWPROT = peripheralUnit_bus_AWPROT; // @[cacheModule.scala 133:22]
  assign peripheral_AWVALID = peripheralUnit_bus_AWVALID; // @[cacheModule.scala 133:22]
  assign peripheral_WDATA = peripheralUnit_bus_WDATA; // @[cacheModule.scala 133:22]
  assign peripheral_WSTRB = peripheralUnit_bus_WSTRB; // @[cacheModule.scala 133:22]
  assign peripheral_WLAST = peripheralUnit_bus_WLAST; // @[cacheModule.scala 133:22]
  assign peripheral_WVALID = peripheralUnit_bus_WVALID; // @[cacheModule.scala 133:22]
  assign peripheral_BREADY = peripheralUnit_bus_BREADY; // @[cacheModule.scala 133:22]
  assign peripheral_ARADDR = peripheralUnit_bus_ARADDR; // @[cacheModule.scala 133:22]
  assign peripheral_ARLEN = peripheralUnit_bus_ARLEN; // @[cacheModule.scala 133:22]
  assign peripheral_ARSIZE = peripheralUnit_bus_ARSIZE; // @[cacheModule.scala 133:22]
  assign peripheral_ARBURST = peripheralUnit_bus_ARBURST; // @[cacheModule.scala 133:22]
  assign peripheral_ARPROT = peripheralUnit_bus_ARPROT; // @[cacheModule.scala 133:22]
  assign peripheral_ARVALID = peripheralUnit_bus_ARVALID; // @[cacheModule.scala 133:22]
  assign peripheral_RREADY = peripheralUnit_bus_RREADY; // @[cacheModule.scala 133:22]
  assign responseOut_valid = cacheLookup_toResponse_request_valid ? cacheLookup_toResponse_request_valid &
    cacheLookup_toResponse_request_branch_valid : peripheralUnit_responseOut_request_valid; // @[cacheModule.scala 139:27]
  assign responseOut_prfDest = cacheLookup_toResponse_request_valid ? cacheLookup_toResponse_request_core_prfDest :
    peripheralUnit_responseOut_request_core_prfDest; // @[cacheModule.scala 141:29]
  assign responseOut_robAddr = cacheLookup_toResponse_request_valid ? cacheLookup_toResponse_request_core_robAddr :
    peripheralUnit_responseOut_request_core_robAddr; // @[cacheModule.scala 142:29]
  assign responseOut_result = cacheLookup_toResponse_request_valid ? cacheLookup_toResponse_request_writeData_data :
    peripheralUnit_responseOut_request_writeData_data; // @[cacheModule.scala 143:28]
  assign responseOut_instruction = cacheLookup_toResponse_request_valid ?
    cacheLookup_toResponse_request_core_instruction : peripheralUnit_responseOut_request_core_instruction; // @[cacheModule.scala 144:33]
  assign canAllocate = fenceInititatedReg ? 1'h0 : requestScheduler_canAllocate & ~commitFifo_isFull; // @[cacheModule.scala 197:27 199:17 73:15]
  assign fenceInstructions_ready = fenceInititatedReg; // @[cacheModule.scala 197:27 198:29 40:27]
  assign writeCommit_ready = arbiter_writeCommit_ready; // @[cacheModule.scala 93:23]
  assign writeInstructionCommit_ready = cacheLookup_writeInstructionCommit_ready ?
    cacheLookup_writeInstructionCommit_ready : peripheralUnit_writeInstructionCommit_ready; // @[cacheModule.scala 146:49 147:40 149:43]
  assign loadCommit_valid = loadCommit_ready & _GEN_30; // @[cacheModule.scala 172:25 43:20]
  assign loadCommit_state = loadCommit_ready & _GEN_29; // @[cacheModule.scala 172:25 44:20]
  assign requestScheduler_clock = clock;
  assign requestScheduler_reset = reset;
  assign requestScheduler_requestIn_valid = request_valid; // @[cacheModule.scala 75:36]
  assign requestScheduler_requestIn_address = request_address; // @[cacheModule.scala 76:38]
  assign requestScheduler_requestIn_core_instruction = request_instruction; // @[cacheModule.scala 77:47]
  assign requestScheduler_requestIn_core_robAddr = request_robAddr; // @[cacheModule.scala 78:43]
  assign requestScheduler_requestIn_core_prfDest = request_prfDest; // @[cacheModule.scala 79:43]
  assign requestScheduler_requestIn_branch_mask = request_branchMask; // @[cacheModule.scala 80:42]
  assign requestScheduler_controlSignal_inorderReady = arbiter_request_inorderReady; // @[cacheModule.scala 98:47]
  assign requestScheduler_controlSignal_speculativeReady = arbiter_request_speculativeReady; // @[cacheModule.scala 99:51]
  assign requestScheduler_branchOps_valid = branchOps_valid; // @[cacheModule.scala 72:30]
  assign requestScheduler_branchOps_branchMask = branchOps_branchMask; // @[cacheModule.scala 72:30]
  assign requestScheduler_branchOps_passed = branchOps_passed; // @[cacheModule.scala 72:30]
  assign arbiter_clock = clock;
  assign arbiter_reset = reset;
  assign arbiter_request_request_valid = requestScheduler_requestOut_valid; // @[cacheModule.scala 101:27]
  assign arbiter_request_request_address = requestScheduler_requestOut_address; // @[cacheModule.scala 101:27]
  assign arbiter_request_request_core_instruction = requestScheduler_requestOut_core_instruction; // @[cacheModule.scala 101:27]
  assign arbiter_request_request_core_robAddr = requestScheduler_requestOut_core_robAddr; // @[cacheModule.scala 101:27]
  assign arbiter_request_request_core_prfDest = requestScheduler_requestOut_core_prfDest; // @[cacheModule.scala 101:27]
  assign arbiter_request_request_branch_valid = requestScheduler_requestOut_branch_valid; // @[cacheModule.scala 101:27]
  assign arbiter_request_request_branch_mask = requestScheduler_requestOut_branch_mask; // @[cacheModule.scala 101:27]
  assign arbiter_request_request_writeData_valid = requestScheduler_requestOut_writeData_valid; // @[cacheModule.scala 101:27]
  assign arbiter_request_request_writeData_data = requestScheduler_requestOut_writeData_data; // @[cacheModule.scala 101:27]
  assign arbiter_request_isSpeculative = requestScheduler_controlSignal_isSpeculative; // @[cacheModule.scala 100:33]
  assign arbiter_toPeripheral_ready = peripheralUnit_request_ready; // @[cacheModule.scala 135:26]
  assign arbiter_toCacheLookup_ready = cacheLookup_request_ready; // @[cacheModule.scala 109:23]
  assign arbiter_toCacheLookup_holdInOrder = cacheLookup_request_holdInOrder; // @[cacheModule.scala 109:23]
  assign arbiter_replayRequest_request_valid = replayUnit_responseOut_request_valid; // @[cacheModule.scala 102:25]
  assign arbiter_replayRequest_request_address = replayUnit_responseOut_request_address; // @[cacheModule.scala 102:25]
  assign arbiter_replayRequest_request_core_instruction = replayUnit_responseOut_request_core_instruction; // @[cacheModule.scala 102:25]
  assign arbiter_replayRequest_request_core_robAddr = replayUnit_responseOut_request_core_robAddr; // @[cacheModule.scala 102:25]
  assign arbiter_replayRequest_request_core_prfDest = replayUnit_responseOut_request_core_prfDest; // @[cacheModule.scala 102:25]
  assign arbiter_replayRequest_request_branch_valid = replayUnit_responseOut_request_branch_valid; // @[cacheModule.scala 102:25]
  assign arbiter_replayRequest_request_branch_mask = replayUnit_responseOut_request_branch_mask; // @[cacheModule.scala 102:25]
  assign arbiter_replayRequest_request_writeData_valid = replayUnit_responseOut_request_writeData_valid; // @[cacheModule.scala 102:25]
  assign arbiter_replayRequest_request_writeData_data = replayUnit_responseOut_request_writeData_data; // @[cacheModule.scala 102:25]
  assign arbiter_replayRequest_request_cacheLine_cacheLine = replayUnit_responseOut_request_cacheLine_cacheLine; // @[cacheModule.scala 102:25]
  assign arbiter_replayRequest_request_cacheLine_response = replayUnit_responseOut_request_cacheLine_response; // @[cacheModule.scala 102:25]
  assign arbiter_coherencyRequest_request_valid = aceUnit_coherencyRequest_request_valid; // @[cacheModule.scala 103:28]
  assign arbiter_coherencyRequest_request_address = aceUnit_coherencyRequest_request_address; // @[cacheModule.scala 103:28]
  assign arbiter_coherencyRequest_request_response = aceUnit_coherencyRequest_request_response; // @[cacheModule.scala 103:28]
  assign arbiter_writeDataIn_valid = writeDataIn_valid; // @[cacheModule.scala 92:23]
  assign arbiter_writeDataIn_data = writeDataIn_data; // @[cacheModule.scala 92:23]
  assign arbiter_writeCommit_fired = writeCommit_fired; // @[cacheModule.scala 93:23]
  assign arbiter_branchOps_valid = branchOps_valid; // @[cacheModule.scala 95:21]
  assign arbiter_branchOps_branchMask = branchOps_branchMask; // @[cacheModule.scala 95:21]
  assign arbiter_branchOps_passed = branchOps_passed; // @[cacheModule.scala 95:21]
  assign arbiter_responseOut_valid = responseOut_valid; // @[cacheModule.scala 94:23]
  assign arbiter_responseOut_instruction = responseOut_instruction; // @[cacheModule.scala 94:23]
  assign arbiter_writeInstuctionCommitFired = writeInstructionCommit_fired; // @[cacheModule.scala 104:38]
  assign cacheLookup_clock = clock;
  assign cacheLookup_reset = reset;
  assign cacheLookup_request_requestType = arbiter_toCacheLookup_requestType; // @[cacheModule.scala 109:23]
  assign cacheLookup_request_request_valid = arbiter_toCacheLookup_request_valid; // @[cacheModule.scala 109:23]
  assign cacheLookup_request_request_address = arbiter_toCacheLookup_request_address; // @[cacheModule.scala 109:23]
  assign cacheLookup_request_request_core_instruction = arbiter_toCacheLookup_request_core_instruction; // @[cacheModule.scala 109:23]
  assign cacheLookup_request_request_core_robAddr = arbiter_toCacheLookup_request_core_robAddr; // @[cacheModule.scala 109:23]
  assign cacheLookup_request_request_core_prfDest = arbiter_toCacheLookup_request_core_prfDest; // @[cacheModule.scala 109:23]
  assign cacheLookup_request_request_branch_valid = arbiter_toCacheLookup_request_branch_valid; // @[cacheModule.scala 109:23]
  assign cacheLookup_request_request_branch_mask = arbiter_toCacheLookup_request_branch_mask; // @[cacheModule.scala 109:23]
  assign cacheLookup_request_request_writeData_valid = arbiter_toCacheLookup_request_writeData_valid; // @[cacheModule.scala 109:23]
  assign cacheLookup_request_request_writeData_data = arbiter_toCacheLookup_request_writeData_data; // @[cacheModule.scala 109:23]
  assign cacheLookup_request_request_cacheLine_cacheLine = arbiter_toCacheLookup_request_cacheLine_cacheLine; // @[cacheModule.scala 109:23]
  assign cacheLookup_request_request_cacheLine_response = arbiter_toCacheLookup_request_cacheLine_response; // @[cacheModule.scala 109:23]
  assign cacheLookup_toReplay_ready = replayUnit_requestIn_ready; // @[cacheModule.scala 118:24]
  assign cacheLookup_toWriteBack_ready = replayUnit_writeBackIn_ready; // @[cacheModule.scala 120:26]
  assign cacheLookup_toCoherency_ready = aceUnit_coherencyResponse_ready; // @[cacheModule.scala 128:29]
  assign cacheLookup_writeInstructionCommit_fired = cacheLookup_writeInstructionCommit_ready &
    writeInstructionCommit_fired; // @[cacheModule.scala 146:49 147:40 110:44]
  assign cacheLookup_branchOps_valid = branchOps_valid; // @[cacheModule.scala 107:25]
  assign cacheLookup_branchOps_branchMask = branchOps_branchMask; // @[cacheModule.scala 107:25]
  assign cacheLookup_branchOps_passed = branchOps_passed; // @[cacheModule.scala 107:25]
  assign replayUnit_clock = clock;
  assign replayUnit_reset = reset;
  assign replayUnit_requestIn_request_valid = cacheLookup_toReplay_request_valid; // @[cacheModule.scala 118:24]
  assign replayUnit_requestIn_request_address = cacheLookup_toReplay_request_address; // @[cacheModule.scala 118:24]
  assign replayUnit_requestIn_request_core_instruction = cacheLookup_toReplay_request_core_instruction; // @[cacheModule.scala 118:24]
  assign replayUnit_requestIn_request_core_robAddr = cacheLookup_toReplay_request_core_robAddr; // @[cacheModule.scala 118:24]
  assign replayUnit_requestIn_request_core_prfDest = cacheLookup_toReplay_request_core_prfDest; // @[cacheModule.scala 118:24]
  assign replayUnit_requestIn_request_branch_valid = cacheLookup_toReplay_request_branch_valid; // @[cacheModule.scala 118:24]
  assign replayUnit_requestIn_request_branch_mask = cacheLookup_toReplay_request_branch_mask; // @[cacheModule.scala 118:24]
  assign replayUnit_requestIn_request_writeData_valid = cacheLookup_toReplay_request_writeData_valid; // @[cacheModule.scala 118:24]
  assign replayUnit_requestIn_request_writeData_data = cacheLookup_toReplay_request_writeData_data; // @[cacheModule.scala 118:24]
  assign replayUnit_requestIn_request_cacheLine_response = cacheLookup_toReplay_request_cacheLine_response; // @[cacheModule.scala 118:24]
  assign replayUnit_requestOut_ready = aceUnit_readRequest_ready; // @[cacheModule.scala 127:23]
  assign replayUnit_responseIn_request_valid = aceUnit_readResponse_request_valid; // @[cacheModule.scala 119:25]
  assign replayUnit_responseIn_request_address = aceUnit_readResponse_request_address; // @[cacheModule.scala 119:25]
  assign replayUnit_responseIn_request_core_instruction = aceUnit_readResponse_request_core_instruction; // @[cacheModule.scala 119:25]
  assign replayUnit_responseIn_request_core_robAddr = aceUnit_readResponse_request_core_robAddr; // @[cacheModule.scala 119:25]
  assign replayUnit_responseIn_request_core_prfDest = aceUnit_readResponse_request_core_prfDest; // @[cacheModule.scala 119:25]
  assign replayUnit_responseIn_request_branch_valid = aceUnit_readResponse_request_branch_valid; // @[cacheModule.scala 119:25]
  assign replayUnit_responseIn_request_branch_mask = aceUnit_readResponse_request_branch_mask; // @[cacheModule.scala 119:25]
  assign replayUnit_responseIn_request_writeData_valid = aceUnit_readResponse_request_writeData_valid; // @[cacheModule.scala 119:25]
  assign replayUnit_responseIn_request_writeData_data = aceUnit_readResponse_request_writeData_data; // @[cacheModule.scala 119:25]
  assign replayUnit_responseIn_request_cacheLine_cacheLine = aceUnit_readResponse_request_cacheLine_cacheLine; // @[cacheModule.scala 119:25]
  assign replayUnit_responseIn_request_cacheLine_response = aceUnit_readResponse_request_cacheLine_response; // @[cacheModule.scala 119:25]
  assign replayUnit_responseOut_ready = arbiter_replayRequest_ready; // @[cacheModule.scala 102:25]
  assign replayUnit_writeBackIn_request_valid = cacheLookup_toWriteBack_request_valid; // @[cacheModule.scala 120:26]
  assign replayUnit_writeBackIn_request_address = cacheLookup_toWriteBack_request_address; // @[cacheModule.scala 120:26]
  assign replayUnit_writeBackIn_request_data = cacheLookup_toWriteBack_request_data; // @[cacheModule.scala 120:26]
  assign replayUnit_writeBackOut_ready = aceUnit_writeRequest_ready; // @[cacheModule.scala 129:24]
  assign replayUnit_branchOps_valid = branchOps_valid; // @[cacheModule.scala 116:24]
  assign replayUnit_branchOps_branchMask = branchOps_branchMask; // @[cacheModule.scala 116:24]
  assign replayUnit_branchOps_passed = branchOps_passed; // @[cacheModule.scala 116:24]
  assign peripheralUnit_clock = clock;
  assign peripheralUnit_reset = reset;
  assign peripheralUnit_request_request_valid = arbiter_toPeripheral_request_valid; // @[cacheModule.scala 135:26]
  assign peripheralUnit_request_request_address = arbiter_toPeripheral_request_address; // @[cacheModule.scala 135:26]
  assign peripheralUnit_request_request_core_instruction = arbiter_toPeripheral_request_core_instruction; // @[cacheModule.scala 135:26]
  assign peripheralUnit_request_request_core_robAddr = arbiter_toPeripheral_request_core_robAddr; // @[cacheModule.scala 135:26]
  assign peripheralUnit_request_request_core_prfDest = arbiter_toPeripheral_request_core_prfDest; // @[cacheModule.scala 135:26]
  assign peripheralUnit_request_request_branch_valid = arbiter_toPeripheral_request_branch_valid; // @[cacheModule.scala 135:26]
  assign peripheralUnit_request_request_branch_mask = arbiter_toPeripheral_request_branch_mask; // @[cacheModule.scala 135:26]
  assign peripheralUnit_request_request_writeData_valid = arbiter_toPeripheral_request_writeData_valid; // @[cacheModule.scala 135:26]
  assign peripheralUnit_request_request_writeData_data = arbiter_toPeripheral_request_writeData_data; // @[cacheModule.scala 135:26]
  assign peripheralUnit_responseOut_ready = ~cacheLookup_toResponse_request_valid; // @[cacheModule.scala 136:39]
  assign peripheralUnit_bus_AWREADY = peripheral_AWREADY; // @[cacheModule.scala 133:22]
  assign peripheralUnit_bus_WREADY = peripheral_WREADY; // @[cacheModule.scala 133:22]
  assign peripheralUnit_bus_BID = peripheral_BID; // @[cacheModule.scala 133:22]
  assign peripheralUnit_bus_BRESP = peripheral_BRESP; // @[cacheModule.scala 133:22]
  assign peripheralUnit_bus_BVALID = peripheral_BVALID; // @[cacheModule.scala 133:22]
  assign peripheralUnit_bus_ARREADY = peripheral_ARREADY; // @[cacheModule.scala 133:22]
  assign peripheralUnit_bus_RID = peripheral_RID; // @[cacheModule.scala 133:22]
  assign peripheralUnit_bus_RDATA = peripheral_RDATA; // @[cacheModule.scala 133:22]
  assign peripheralUnit_bus_RRESP = peripheral_RRESP; // @[cacheModule.scala 133:22]
  assign peripheralUnit_bus_RLAST = peripheral_RLAST; // @[cacheModule.scala 133:22]
  assign peripheralUnit_bus_RVALID = peripheral_RVALID; // @[cacheModule.scala 133:22]
  assign peripheralUnit_writeInstructionCommit_fired = cacheLookup_writeInstructionCommit_ready ? 1'h0 :
    writeInstructionCommit_fired; // @[cacheModule.scala 137:47 146:49 149:43]
  assign peripheralUnit_branchOps_valid = branchOps_valid; // @[cacheModule.scala 132:28]
  assign peripheralUnit_branchOps_branchMask = branchOps_branchMask; // @[cacheModule.scala 132:28]
  assign peripheralUnit_branchOps_passed = branchOps_passed; // @[cacheModule.scala 132:28]
  assign aceUnit_clock = clock;
  assign aceUnit_reset = reset;
  assign aceUnit_readRequest_request_valid = replayUnit_requestOut_request_valid; // @[cacheModule.scala 127:23]
  assign aceUnit_readRequest_request_address = replayUnit_requestOut_request_address; // @[cacheModule.scala 127:23]
  assign aceUnit_readRequest_request_core_instruction = replayUnit_requestOut_request_core_instruction; // @[cacheModule.scala 127:23]
  assign aceUnit_readRequest_request_core_robAddr = replayUnit_requestOut_request_core_robAddr; // @[cacheModule.scala 127:23]
  assign aceUnit_readRequest_request_core_prfDest = replayUnit_requestOut_request_core_prfDest; // @[cacheModule.scala 127:23]
  assign aceUnit_readRequest_request_branch_valid = replayUnit_requestOut_request_branch_valid; // @[cacheModule.scala 127:23]
  assign aceUnit_readRequest_request_branch_mask = replayUnit_requestOut_request_branch_mask; // @[cacheModule.scala 127:23]
  assign aceUnit_readRequest_request_writeData_valid = replayUnit_requestOut_request_writeData_valid; // @[cacheModule.scala 127:23]
  assign aceUnit_readRequest_request_writeData_data = replayUnit_requestOut_request_writeData_data; // @[cacheModule.scala 127:23]
  assign aceUnit_readRequest_request_cacheLine_response = replayUnit_requestOut_request_cacheLine_response; // @[cacheModule.scala 127:23]
  assign aceUnit_readResponse_ready = replayUnit_responseIn_ready; // @[cacheModule.scala 119:25]
  assign aceUnit_writeRequest_request_valid = replayUnit_writeBackOut_request_valid; // @[cacheModule.scala 129:24]
  assign aceUnit_writeRequest_request_address = replayUnit_writeBackOut_request_address; // @[cacheModule.scala 129:24]
  assign aceUnit_writeRequest_request_data = replayUnit_writeBackOut_request_data; // @[cacheModule.scala 129:24]
  assign aceUnit_coherencyRequest_ready = arbiter_coherencyRequest_ready; // @[cacheModule.scala 103:28]
  assign aceUnit_coherencyResponse_request_valid = cacheLookup_toCoherency_request_valid; // @[cacheModule.scala 128:29]
  assign aceUnit_coherencyResponse_request_response = cacheLookup_toCoherency_request_response; // @[cacheModule.scala 128:29]
  assign aceUnit_coherencyResponse_request_cacheLine = cacheLookup_toCoherency_request_cacheLine; // @[cacheModule.scala 128:29]
  assign aceUnit_coherencyResponse_request_dataValid = cacheLookup_toCoherency_request_dataValid; // @[cacheModule.scala 128:29]
  assign aceUnit_branchOps_valid = branchOps_valid; // @[cacheModule.scala 124:21]
  assign aceUnit_branchOps_branchMask = branchOps_branchMask; // @[cacheModule.scala 124:21]
  assign aceUnit_branchOps_passed = branchOps_passed; // @[cacheModule.scala 124:21]
  assign aceUnit_bus_AWREADY = dPort_AWREADY; // @[cacheModule.scala 125:15]
  assign aceUnit_bus_WREADY = dPort_WREADY; // @[cacheModule.scala 125:15]
  assign aceUnit_bus_BRESP = dPort_BRESP; // @[cacheModule.scala 125:15]
  assign aceUnit_bus_BVALID = dPort_BVALID; // @[cacheModule.scala 125:15]
  assign aceUnit_bus_ARREADY = dPort_ARREADY; // @[cacheModule.scala 125:15]
  assign aceUnit_bus_RDATA = dPort_RDATA; // @[cacheModule.scala 125:15]
  assign aceUnit_bus_RLAST = dPort_RLAST; // @[cacheModule.scala 125:15]
  assign aceUnit_bus_RVALID = dPort_RVALID; // @[cacheModule.scala 125:15]
  assign aceUnit_bus_RRESP = dPort_RRESP; // @[cacheModule.scala 125:15]
  assign aceUnit_bus_ACVALID = dPort_ACVALID; // @[cacheModule.scala 125:15]
  assign aceUnit_bus_ACADDR = dPort_ACADDR; // @[cacheModule.scala 125:15]
  assign aceUnit_bus_ACSNOOP = dPort_ACSNOOP; // @[cacheModule.scala 125:15]
  assign aceUnit_bus_CRREADY = dPort_CRREADY; // @[cacheModule.scala 125:15]
  assign aceUnit_bus_CDREADY = dPort_CDREADY; // @[cacheModule.scala 125:15]
  assign commitFifo_clock = clock;
  assign commitFifo_reset = reset;
  assign commitFifo_write_data_valid = _responseOut_valid_T & cacheLookup_toResponse_request_core_instruction[6:0] == 7'h3
     ? cacheLookup_toResponse_request_valid : _GEN_14; // @[cacheModule.scala 159:165 160:27]
  assign commitFifo_write_data_address = _responseOut_valid_T & cacheLookup_toResponse_request_core_instruction[6:0] == 7'h3
     ? cacheLookup_toResponse_request_address : _GEN_13; // @[cacheModule.scala 159:165 160:27]
  assign commitFifo_write_data_branch_valid = _responseOut_valid_T & cacheLookup_toResponse_request_core_instruction[6:0
    ] == 7'h3 ? cacheLookup_toResponse_request_branch_valid : _GEN_9; // @[cacheModule.scala 159:165 160:27]
  assign commitFifo_write_data_branch_mask = _responseOut_valid_T & cacheLookup_toResponse_request_core_instruction[6:0]
     == 7'h3 ? cacheLookup_toResponse_request_branch_mask : _GEN_8; // @[cacheModule.scala 159:165 160:27]
  assign commitFifo_read_ready = loadCommit_ready; // @[cacheModule.scala 154:25 172:25 173:27]
  assign commitFifo_branchOps_valid = branchOps_valid; // @[cacheModule.scala 165:24]
  assign commitFifo_branchOps_branchMask = branchOps_branchMask; // @[cacheModule.scala 165:24]
  assign commitFifo_branchOps_passed = branchOps_passed; // @[cacheModule.scala 165:24]
  assign commitFifo_invalidateAddr = aceUnit_coherencyRequest_request_valid & aceUnit_coherencyRequest_request_response[
    1] ? aceUnit_coherencyRequest_request_address : 32'h0; // @[cacheModule.scala 155:29 167:95 168:31]
  assign commitFifo_invalidateEnable = aceUnit_coherencyRequest_request_valid &
    aceUnit_coherencyRequest_request_response[1]; // @[cacheModule.scala 167:47]
  always @(posedge clock) begin
    if (reset) begin // @[cacheModule.scala 183:35]
      fenceInititatedReg <= 1'h0; // @[cacheModule.scala 183:35]
    end else if (fenceInititatedReg) begin // @[cacheModule.scala 197:27]
      if (fenceInstructions_fired) begin // @[cacheModule.scala 200:30]
        fenceInititatedReg <= 1'h0;
      end else begin
        fenceInititatedReg <= 1'h1;
      end
    end else begin
      fenceInititatedReg <= canInititatedFenceReg & subModulesReady; // @[cacheModule.scala 195:22]
    end
    if (reset) begin // @[cacheModule.scala 184:38]
      canInititatedFenceReg <= 1'h0; // @[cacheModule.scala 184:38]
    end else if (fenceInititatedReg) begin // @[cacheModule.scala 197:27]
      if (fenceInstructions_fired) begin // @[cacheModule.scala 200:30]
        canInititatedFenceReg <= 1'h0;
      end else begin
        canInititatedFenceReg <= 1'h1;
      end
    end else if (~canInititatedFenceReg) begin // @[cacheModule.scala 193:31]
      canInititatedFenceReg <= initiateFence;
    end
    subModulesReady_REG <= ~cacheLookup_request_holdInOrder; // @[cacheModule.scala 190:21]
    subModulesReady_REG_1 <= subModulesReady_REG; // @[cacheModule.scala 190:12]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fenceInititatedReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  canInititatedFenceReg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  subModulesReady_REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  subModulesReady_REG_1 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReadWriteSmem(
  input         clock,
  input         io_wenable,
  input         io_renable,
  input  [5:0]  io_raddr,
  input  [5:0]  io_waddr,
  input  [63:0] io_dataIn,
  output [63:0] io_dataOut
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mem [0:63]; // @[SRAM_block.scala 15:24]
  wire  mem_io_dataOut_MPORT_en; // @[SRAM_block.scala 15:24]
  wire [5:0] mem_io_dataOut_MPORT_addr; // @[SRAM_block.scala 15:24]
  wire [63:0] mem_io_dataOut_MPORT_data; // @[SRAM_block.scala 15:24]
  wire [63:0] mem_MPORT_data; // @[SRAM_block.scala 15:24]
  wire [5:0] mem_MPORT_addr; // @[SRAM_block.scala 15:24]
  wire  mem_MPORT_mask; // @[SRAM_block.scala 15:24]
  wire  mem_MPORT_en; // @[SRAM_block.scala 15:24]
  reg  mem_io_dataOut_MPORT_en_pipe_0;
  reg [5:0] mem_io_dataOut_MPORT_addr_pipe_0;
  assign mem_io_dataOut_MPORT_en = mem_io_dataOut_MPORT_en_pipe_0;
  assign mem_io_dataOut_MPORT_addr = mem_io_dataOut_MPORT_addr_pipe_0;
  assign mem_io_dataOut_MPORT_data = mem[mem_io_dataOut_MPORT_addr]; // @[SRAM_block.scala 15:24]
  assign mem_MPORT_data = io_dataIn;
  assign mem_MPORT_addr = io_waddr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_wenable;
  assign io_dataOut = mem_io_dataOut_MPORT_data; // @[SRAM_block.scala 21:14]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SRAM_block.scala 15:24]
    end
    mem_io_dataOut_MPORT_en_pipe_0 <= io_renable;
    if (io_renable) begin
      mem_io_dataOut_MPORT_addr_pipe_0 <= io_raddr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    mem[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_dataOut_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_dataOut_MPORT_addr_pipe_0 = _RAND_2[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LVT_set(
  input         clock,
  input         io_wenable,
  input         io_r1enable,
  input         io_r2enable,
  input         io_r3enable,
  input  [5:0]  io_r1addr,
  input  [5:0]  io_r2addr,
  input  [5:0]  io_r3addr,
  input  [5:0]  io_waddr,
  input  [63:0] io_wdata,
  output [63:0] io_r1data,
  output [63:0] io_r2data,
  output [63:0] io_r3data
);
  wire  b1_clock; // @[LVT_set.scala 20:18]
  wire  b1_io_wenable; // @[LVT_set.scala 20:18]
  wire  b1_io_renable; // @[LVT_set.scala 20:18]
  wire [5:0] b1_io_raddr; // @[LVT_set.scala 20:18]
  wire [5:0] b1_io_waddr; // @[LVT_set.scala 20:18]
  wire [63:0] b1_io_dataIn; // @[LVT_set.scala 20:18]
  wire [63:0] b1_io_dataOut; // @[LVT_set.scala 20:18]
  wire  b2_clock; // @[LVT_set.scala 21:18]
  wire  b2_io_wenable; // @[LVT_set.scala 21:18]
  wire  b2_io_renable; // @[LVT_set.scala 21:18]
  wire [5:0] b2_io_raddr; // @[LVT_set.scala 21:18]
  wire [5:0] b2_io_waddr; // @[LVT_set.scala 21:18]
  wire [63:0] b2_io_dataIn; // @[LVT_set.scala 21:18]
  wire [63:0] b2_io_dataOut; // @[LVT_set.scala 21:18]
  wire  b3_clock; // @[LVT_set.scala 22:18]
  wire  b3_io_wenable; // @[LVT_set.scala 22:18]
  wire  b3_io_renable; // @[LVT_set.scala 22:18]
  wire [5:0] b3_io_raddr; // @[LVT_set.scala 22:18]
  wire [5:0] b3_io_waddr; // @[LVT_set.scala 22:18]
  wire [63:0] b3_io_dataIn; // @[LVT_set.scala 22:18]
  wire [63:0] b3_io_dataOut; // @[LVT_set.scala 22:18]
  ReadWriteSmem b1 ( // @[LVT_set.scala 20:18]
    .clock(b1_clock),
    .io_wenable(b1_io_wenable),
    .io_renable(b1_io_renable),
    .io_raddr(b1_io_raddr),
    .io_waddr(b1_io_waddr),
    .io_dataIn(b1_io_dataIn),
    .io_dataOut(b1_io_dataOut)
  );
  ReadWriteSmem b2 ( // @[LVT_set.scala 21:18]
    .clock(b2_clock),
    .io_wenable(b2_io_wenable),
    .io_renable(b2_io_renable),
    .io_raddr(b2_io_raddr),
    .io_waddr(b2_io_waddr),
    .io_dataIn(b2_io_dataIn),
    .io_dataOut(b2_io_dataOut)
  );
  ReadWriteSmem b3 ( // @[LVT_set.scala 22:18]
    .clock(b3_clock),
    .io_wenable(b3_io_wenable),
    .io_renable(b3_io_renable),
    .io_raddr(b3_io_raddr),
    .io_waddr(b3_io_waddr),
    .io_dataIn(b3_io_dataIn),
    .io_dataOut(b3_io_dataOut)
  );
  assign io_r1data = b1_io_dataOut; // @[LVT_set.scala 35:13]
  assign io_r2data = b2_io_dataOut; // @[LVT_set.scala 36:13]
  assign io_r3data = b3_io_dataOut; // @[LVT_set.scala 37:13]
  assign b1_clock = clock;
  assign b1_io_wenable = io_wenable; // @[LVT_set.scala 24:17]
  assign b1_io_renable = io_r1enable; // @[LVT_set.scala 31:17]
  assign b1_io_raddr = io_r1addr; // @[LVT_set.scala 39:15]
  assign b1_io_waddr = io_waddr; // @[LVT_set.scala 43:15]
  assign b1_io_dataIn = io_wdata; // @[LVT_set.scala 27:16]
  assign b2_clock = clock;
  assign b2_io_wenable = io_wenable; // @[LVT_set.scala 25:17]
  assign b2_io_renable = io_r2enable; // @[LVT_set.scala 32:17]
  assign b2_io_raddr = io_r2addr; // @[LVT_set.scala 40:15]
  assign b2_io_waddr = io_waddr; // @[LVT_set.scala 44:15]
  assign b2_io_dataIn = io_wdata; // @[LVT_set.scala 28:16]
  assign b3_clock = clock;
  assign b3_io_wenable = io_wenable; // @[LVT_set.scala 26:17]
  assign b3_io_renable = io_r3enable; // @[LVT_set.scala 33:17]
  assign b3_io_raddr = io_r3addr; // @[LVT_set.scala 41:15]
  assign b3_io_waddr = io_waddr; // @[LVT_set.scala 45:15]
  assign b3_io_dataIn = io_wdata; // @[LVT_set.scala 29:16]
endmodule
module LVT_Mem(
  input         clock,
  input         reset,
  input  [5:0]  io_R1_addr,
  output [63:0] io_R1_data,
  input         io_R1_en,
  input  [5:0]  io_R2_addr,
  output [63:0] io_R2_data,
  input         io_R2_en,
  input  [5:0]  io_R3_addr,
  output [63:0] io_R3_data,
  input         io_R3_en,
  input  [5:0]  io_W1_addr,
  input  [63:0] io_W1_data,
  input         io_W1_en,
  input  [5:0]  io_W2_addr,
  input  [63:0] io_W2_data,
  input         io_W2_en,
  input  [5:0]  io_W3_addr,
  input  [63:0] io_W3_data,
  input         io_W3_en,
  input  [5:0]  io_W4_addr,
  input  [63:0] io_W4_data,
  input         io_W4_en
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] LVT [0:63]; // @[LVT_Mem.scala 32:16]
  wire  LVT_r1_sel_reg_MPORT_en; // @[LVT_Mem.scala 32:16]
  wire [5:0] LVT_r1_sel_reg_MPORT_addr; // @[LVT_Mem.scala 32:16]
  wire [1:0] LVT_r1_sel_reg_MPORT_data; // @[LVT_Mem.scala 32:16]
  wire  LVT_r2_sel_reg_MPORT_en; // @[LVT_Mem.scala 32:16]
  wire [5:0] LVT_r2_sel_reg_MPORT_addr; // @[LVT_Mem.scala 32:16]
  wire [1:0] LVT_r2_sel_reg_MPORT_data; // @[LVT_Mem.scala 32:16]
  wire  LVT_r3_sel_reg_MPORT_en; // @[LVT_Mem.scala 32:16]
  wire [5:0] LVT_r3_sel_reg_MPORT_addr; // @[LVT_Mem.scala 32:16]
  wire [1:0] LVT_r3_sel_reg_MPORT_data; // @[LVT_Mem.scala 32:16]
  wire [1:0] LVT_MPORT_data; // @[LVT_Mem.scala 32:16]
  wire [5:0] LVT_MPORT_addr; // @[LVT_Mem.scala 32:16]
  wire  LVT_MPORT_mask; // @[LVT_Mem.scala 32:16]
  wire  LVT_MPORT_en; // @[LVT_Mem.scala 32:16]
  wire [1:0] LVT_MPORT_1_data; // @[LVT_Mem.scala 32:16]
  wire [5:0] LVT_MPORT_1_addr; // @[LVT_Mem.scala 32:16]
  wire  LVT_MPORT_1_mask; // @[LVT_Mem.scala 32:16]
  wire  LVT_MPORT_1_en; // @[LVT_Mem.scala 32:16]
  wire [1:0] LVT_MPORT_2_data; // @[LVT_Mem.scala 32:16]
  wire [5:0] LVT_MPORT_2_addr; // @[LVT_Mem.scala 32:16]
  wire  LVT_MPORT_2_mask; // @[LVT_Mem.scala 32:16]
  wire  LVT_MPORT_2_en; // @[LVT_Mem.scala 32:16]
  wire [1:0] LVT_MPORT_3_data; // @[LVT_Mem.scala 32:16]
  wire [5:0] LVT_MPORT_3_addr; // @[LVT_Mem.scala 32:16]
  wire  LVT_MPORT_3_mask; // @[LVT_Mem.scala 32:16]
  wire  LVT_MPORT_3_en; // @[LVT_Mem.scala 32:16]
  wire  s1_clock; // @[LVT_Mem.scala 35:18]
  wire  s1_io_wenable; // @[LVT_Mem.scala 35:18]
  wire  s1_io_r1enable; // @[LVT_Mem.scala 35:18]
  wire  s1_io_r2enable; // @[LVT_Mem.scala 35:18]
  wire  s1_io_r3enable; // @[LVT_Mem.scala 35:18]
  wire [5:0] s1_io_r1addr; // @[LVT_Mem.scala 35:18]
  wire [5:0] s1_io_r2addr; // @[LVT_Mem.scala 35:18]
  wire [5:0] s1_io_r3addr; // @[LVT_Mem.scala 35:18]
  wire [5:0] s1_io_waddr; // @[LVT_Mem.scala 35:18]
  wire [63:0] s1_io_wdata; // @[LVT_Mem.scala 35:18]
  wire [63:0] s1_io_r1data; // @[LVT_Mem.scala 35:18]
  wire [63:0] s1_io_r2data; // @[LVT_Mem.scala 35:18]
  wire [63:0] s1_io_r3data; // @[LVT_Mem.scala 35:18]
  wire  s2_clock; // @[LVT_Mem.scala 36:18]
  wire  s2_io_wenable; // @[LVT_Mem.scala 36:18]
  wire  s2_io_r1enable; // @[LVT_Mem.scala 36:18]
  wire  s2_io_r2enable; // @[LVT_Mem.scala 36:18]
  wire  s2_io_r3enable; // @[LVT_Mem.scala 36:18]
  wire [5:0] s2_io_r1addr; // @[LVT_Mem.scala 36:18]
  wire [5:0] s2_io_r2addr; // @[LVT_Mem.scala 36:18]
  wire [5:0] s2_io_r3addr; // @[LVT_Mem.scala 36:18]
  wire [5:0] s2_io_waddr; // @[LVT_Mem.scala 36:18]
  wire [63:0] s2_io_wdata; // @[LVT_Mem.scala 36:18]
  wire [63:0] s2_io_r1data; // @[LVT_Mem.scala 36:18]
  wire [63:0] s2_io_r2data; // @[LVT_Mem.scala 36:18]
  wire [63:0] s2_io_r3data; // @[LVT_Mem.scala 36:18]
  wire  s3_clock; // @[LVT_Mem.scala 37:18]
  wire  s3_io_wenable; // @[LVT_Mem.scala 37:18]
  wire  s3_io_r1enable; // @[LVT_Mem.scala 37:18]
  wire  s3_io_r2enable; // @[LVT_Mem.scala 37:18]
  wire  s3_io_r3enable; // @[LVT_Mem.scala 37:18]
  wire [5:0] s3_io_r1addr; // @[LVT_Mem.scala 37:18]
  wire [5:0] s3_io_r2addr; // @[LVT_Mem.scala 37:18]
  wire [5:0] s3_io_r3addr; // @[LVT_Mem.scala 37:18]
  wire [5:0] s3_io_waddr; // @[LVT_Mem.scala 37:18]
  wire [63:0] s3_io_wdata; // @[LVT_Mem.scala 37:18]
  wire [63:0] s3_io_r1data; // @[LVT_Mem.scala 37:18]
  wire [63:0] s3_io_r2data; // @[LVT_Mem.scala 37:18]
  wire [63:0] s3_io_r3data; // @[LVT_Mem.scala 37:18]
  wire  s4_clock; // @[LVT_Mem.scala 38:18]
  wire  s4_io_wenable; // @[LVT_Mem.scala 38:18]
  wire  s4_io_r1enable; // @[LVT_Mem.scala 38:18]
  wire  s4_io_r2enable; // @[LVT_Mem.scala 38:18]
  wire  s4_io_r3enable; // @[LVT_Mem.scala 38:18]
  wire [5:0] s4_io_r1addr; // @[LVT_Mem.scala 38:18]
  wire [5:0] s4_io_r2addr; // @[LVT_Mem.scala 38:18]
  wire [5:0] s4_io_r3addr; // @[LVT_Mem.scala 38:18]
  wire [5:0] s4_io_waddr; // @[LVT_Mem.scala 38:18]
  wire [63:0] s4_io_wdata; // @[LVT_Mem.scala 38:18]
  wire [63:0] s4_io_r1data; // @[LVT_Mem.scala 38:18]
  wire [63:0] s4_io_r2data; // @[LVT_Mem.scala 38:18]
  wire [63:0] s4_io_r3data; // @[LVT_Mem.scala 38:18]
  reg [1:0] r1_sel_reg; // @[LVT_Mem.scala 69:27]
  reg [1:0] r2_sel_reg; // @[LVT_Mem.scala 70:27]
  reg [1:0] r3_sel_reg; // @[LVT_Mem.scala 71:27]
  wire  _io_R1_data_T = r1_sel_reg == 2'h0; // @[LVT_Mem.scala 110:45]
  wire  _io_R1_data_T_1 = r1_sel_reg == 2'h1; // @[LVT_Mem.scala 110:79]
  wire  _io_R1_data_T_2 = r1_sel_reg == 2'h2; // @[LVT_Mem.scala 110:113]
  wire  _io_R1_data_T_3 = r1_sel_reg == 2'h3; // @[LVT_Mem.scala 110:147]
  wire [63:0] _io_R1_data_T_4 = _io_R1_data_T_3 ? s4_io_r1data : 64'h0; // @[Mux.scala 101:16]
  wire [63:0] _io_R1_data_T_5 = _io_R1_data_T_2 ? s3_io_r1data : _io_R1_data_T_4; // @[Mux.scala 101:16]
  wire [63:0] _io_R1_data_T_6 = _io_R1_data_T_1 ? s2_io_r1data : _io_R1_data_T_5; // @[Mux.scala 101:16]
  wire  _io_R2_data_T = r2_sel_reg == 2'h0; // @[LVT_Mem.scala 111:45]
  wire  _io_R2_data_T_1 = r2_sel_reg == 2'h1; // @[LVT_Mem.scala 111:79]
  wire  _io_R2_data_T_2 = r2_sel_reg == 2'h2; // @[LVT_Mem.scala 111:113]
  wire  _io_R2_data_T_3 = r2_sel_reg == 2'h3; // @[LVT_Mem.scala 111:147]
  wire [63:0] _io_R2_data_T_4 = _io_R2_data_T_3 ? s4_io_r2data : 64'h0; // @[Mux.scala 101:16]
  wire [63:0] _io_R2_data_T_5 = _io_R2_data_T_2 ? s3_io_r2data : _io_R2_data_T_4; // @[Mux.scala 101:16]
  wire [63:0] _io_R2_data_T_6 = _io_R2_data_T_1 ? s2_io_r2data : _io_R2_data_T_5; // @[Mux.scala 101:16]
  wire  _io_R3_data_T = r3_sel_reg == 2'h0; // @[LVT_Mem.scala 112:45]
  wire  _io_R3_data_T_1 = r3_sel_reg == 2'h1; // @[LVT_Mem.scala 112:79]
  wire  _io_R3_data_T_2 = r3_sel_reg == 2'h2; // @[LVT_Mem.scala 112:113]
  wire  _io_R3_data_T_3 = r3_sel_reg == 2'h3; // @[LVT_Mem.scala 112:147]
  wire [63:0] _io_R3_data_T_4 = _io_R3_data_T_3 ? s4_io_r3data : 64'h0; // @[Mux.scala 101:16]
  wire [63:0] _io_R3_data_T_5 = _io_R3_data_T_2 ? s3_io_r3data : _io_R3_data_T_4; // @[Mux.scala 101:16]
  wire [63:0] _io_R3_data_T_6 = _io_R3_data_T_1 ? s2_io_r3data : _io_R3_data_T_5; // @[Mux.scala 101:16]
  LVT_set s1 ( // @[LVT_Mem.scala 35:18]
    .clock(s1_clock),
    .io_wenable(s1_io_wenable),
    .io_r1enable(s1_io_r1enable),
    .io_r2enable(s1_io_r2enable),
    .io_r3enable(s1_io_r3enable),
    .io_r1addr(s1_io_r1addr),
    .io_r2addr(s1_io_r2addr),
    .io_r3addr(s1_io_r3addr),
    .io_waddr(s1_io_waddr),
    .io_wdata(s1_io_wdata),
    .io_r1data(s1_io_r1data),
    .io_r2data(s1_io_r2data),
    .io_r3data(s1_io_r3data)
  );
  LVT_set s2 ( // @[LVT_Mem.scala 36:18]
    .clock(s2_clock),
    .io_wenable(s2_io_wenable),
    .io_r1enable(s2_io_r1enable),
    .io_r2enable(s2_io_r2enable),
    .io_r3enable(s2_io_r3enable),
    .io_r1addr(s2_io_r1addr),
    .io_r2addr(s2_io_r2addr),
    .io_r3addr(s2_io_r3addr),
    .io_waddr(s2_io_waddr),
    .io_wdata(s2_io_wdata),
    .io_r1data(s2_io_r1data),
    .io_r2data(s2_io_r2data),
    .io_r3data(s2_io_r3data)
  );
  LVT_set s3 ( // @[LVT_Mem.scala 37:18]
    .clock(s3_clock),
    .io_wenable(s3_io_wenable),
    .io_r1enable(s3_io_r1enable),
    .io_r2enable(s3_io_r2enable),
    .io_r3enable(s3_io_r3enable),
    .io_r1addr(s3_io_r1addr),
    .io_r2addr(s3_io_r2addr),
    .io_r3addr(s3_io_r3addr),
    .io_waddr(s3_io_waddr),
    .io_wdata(s3_io_wdata),
    .io_r1data(s3_io_r1data),
    .io_r2data(s3_io_r2data),
    .io_r3data(s3_io_r3data)
  );
  LVT_set s4 ( // @[LVT_Mem.scala 38:18]
    .clock(s4_clock),
    .io_wenable(s4_io_wenable),
    .io_r1enable(s4_io_r1enable),
    .io_r2enable(s4_io_r2enable),
    .io_r3enable(s4_io_r3enable),
    .io_r1addr(s4_io_r1addr),
    .io_r2addr(s4_io_r2addr),
    .io_r3addr(s4_io_r3addr),
    .io_waddr(s4_io_waddr),
    .io_wdata(s4_io_wdata),
    .io_r1data(s4_io_r1data),
    .io_r2data(s4_io_r2data),
    .io_r3data(s4_io_r3data)
  );
  assign LVT_r1_sel_reg_MPORT_en = 1'h1;
  assign LVT_r1_sel_reg_MPORT_addr = io_R1_addr;
  assign LVT_r1_sel_reg_MPORT_data = LVT[LVT_r1_sel_reg_MPORT_addr]; // @[LVT_Mem.scala 32:16]
  assign LVT_r2_sel_reg_MPORT_en = 1'h1;
  assign LVT_r2_sel_reg_MPORT_addr = io_R2_addr;
  assign LVT_r2_sel_reg_MPORT_data = LVT[LVT_r2_sel_reg_MPORT_addr]; // @[LVT_Mem.scala 32:16]
  assign LVT_r3_sel_reg_MPORT_en = 1'h1;
  assign LVT_r3_sel_reg_MPORT_addr = io_R3_addr;
  assign LVT_r3_sel_reg_MPORT_data = LVT[LVT_r3_sel_reg_MPORT_addr]; // @[LVT_Mem.scala 32:16]
  assign LVT_MPORT_data = 2'h0;
  assign LVT_MPORT_addr = io_W1_addr;
  assign LVT_MPORT_mask = 1'h1;
  assign LVT_MPORT_en = io_W1_en;
  assign LVT_MPORT_1_data = 2'h1;
  assign LVT_MPORT_1_addr = io_W2_addr;
  assign LVT_MPORT_1_mask = 1'h1;
  assign LVT_MPORT_1_en = io_W2_en;
  assign LVT_MPORT_2_data = 2'h2;
  assign LVT_MPORT_2_addr = io_W3_addr;
  assign LVT_MPORT_2_mask = 1'h1;
  assign LVT_MPORT_2_en = io_W3_en;
  assign LVT_MPORT_3_data = 2'h3;
  assign LVT_MPORT_3_addr = io_W4_addr;
  assign LVT_MPORT_3_mask = 1'h1;
  assign LVT_MPORT_3_en = io_W4_en;
  assign io_R1_data = _io_R1_data_T ? s1_io_r1data : _io_R1_data_T_6; // @[Mux.scala 101:16]
  assign io_R2_data = _io_R2_data_T ? s1_io_r2data : _io_R2_data_T_6; // @[Mux.scala 101:16]
  assign io_R3_data = _io_R3_data_T ? s1_io_r3data : _io_R3_data_T_6; // @[Mux.scala 101:16]
  assign s1_clock = clock;
  assign s1_io_wenable = io_W1_en; // @[LVT_Mem.scala 55:17]
  assign s1_io_r1enable = io_R1_en; // @[LVT_Mem.scala 93:18]
  assign s1_io_r2enable = io_R2_en; // @[LVT_Mem.scala 98:18]
  assign s1_io_r3enable = io_R3_en; // @[LVT_Mem.scala 103:18]
  assign s1_io_r1addr = io_R1_addr; // @[LVT_Mem.scala 78:16]
  assign s1_io_r2addr = io_R2_addr; // @[LVT_Mem.scala 83:16]
  assign s1_io_r3addr = io_R3_addr; // @[LVT_Mem.scala 88:16]
  assign s1_io_waddr = io_W1_addr; // @[LVT_Mem.scala 63:15]
  assign s1_io_wdata = io_W1_data; // @[LVT_Mem.scala 59:15]
  assign s2_clock = clock;
  assign s2_io_wenable = io_W2_en; // @[LVT_Mem.scala 56:17]
  assign s2_io_r1enable = io_R1_en; // @[LVT_Mem.scala 94:18]
  assign s2_io_r2enable = io_R2_en; // @[LVT_Mem.scala 99:18]
  assign s2_io_r3enable = io_R3_en; // @[LVT_Mem.scala 104:18]
  assign s2_io_r1addr = io_R1_addr; // @[LVT_Mem.scala 79:16]
  assign s2_io_r2addr = io_R2_addr; // @[LVT_Mem.scala 84:16]
  assign s2_io_r3addr = io_R3_addr; // @[LVT_Mem.scala 89:16]
  assign s2_io_waddr = io_W2_addr; // @[LVT_Mem.scala 64:15]
  assign s2_io_wdata = io_W2_data; // @[LVT_Mem.scala 60:15]
  assign s3_clock = clock;
  assign s3_io_wenable = io_W3_en; // @[LVT_Mem.scala 57:17]
  assign s3_io_r1enable = io_R1_en; // @[LVT_Mem.scala 95:18]
  assign s3_io_r2enable = io_R2_en; // @[LVT_Mem.scala 100:18]
  assign s3_io_r3enable = io_R3_en; // @[LVT_Mem.scala 105:18]
  assign s3_io_r1addr = io_R1_addr; // @[LVT_Mem.scala 80:16]
  assign s3_io_r2addr = io_R2_addr; // @[LVT_Mem.scala 85:16]
  assign s3_io_r3addr = io_R3_addr; // @[LVT_Mem.scala 90:16]
  assign s3_io_waddr = io_W3_addr; // @[LVT_Mem.scala 65:15]
  assign s3_io_wdata = io_W3_data; // @[LVT_Mem.scala 61:15]
  assign s4_clock = clock;
  assign s4_io_wenable = io_W4_en; // @[LVT_Mem.scala 58:17]
  assign s4_io_r1enable = io_R1_en; // @[LVT_Mem.scala 96:18]
  assign s4_io_r2enable = io_R2_en; // @[LVT_Mem.scala 101:18]
  assign s4_io_r3enable = io_R3_en; // @[LVT_Mem.scala 106:18]
  assign s4_io_r1addr = io_R1_addr; // @[LVT_Mem.scala 81:16]
  assign s4_io_r2addr = io_R2_addr; // @[LVT_Mem.scala 86:16]
  assign s4_io_r3addr = io_R3_addr; // @[LVT_Mem.scala 91:16]
  assign s4_io_waddr = io_W4_addr; // @[LVT_Mem.scala 66:15]
  assign s4_io_wdata = io_W4_data; // @[LVT_Mem.scala 62:15]
  always @(posedge clock) begin
    if (LVT_MPORT_en & LVT_MPORT_mask) begin
      LVT[LVT_MPORT_addr] <= LVT_MPORT_data; // @[LVT_Mem.scala 32:16]
    end
    if (LVT_MPORT_1_en & LVT_MPORT_1_mask) begin
      LVT[LVT_MPORT_1_addr] <= LVT_MPORT_1_data; // @[LVT_Mem.scala 32:16]
    end
    if (LVT_MPORT_2_en & LVT_MPORT_2_mask) begin
      LVT[LVT_MPORT_2_addr] <= LVT_MPORT_2_data; // @[LVT_Mem.scala 32:16]
    end
    if (LVT_MPORT_3_en & LVT_MPORT_3_mask) begin
      LVT[LVT_MPORT_3_addr] <= LVT_MPORT_3_data; // @[LVT_Mem.scala 32:16]
    end
    if (reset) begin // @[LVT_Mem.scala 69:27]
      r1_sel_reg <= 2'h0; // @[LVT_Mem.scala 69:27]
    end else begin
      r1_sel_reg <= LVT_r1_sel_reg_MPORT_data; // @[LVT_Mem.scala 73:14]
    end
    if (reset) begin // @[LVT_Mem.scala 70:27]
      r2_sel_reg <= 2'h0; // @[LVT_Mem.scala 70:27]
    end else begin
      r2_sel_reg <= LVT_r2_sel_reg_MPORT_data; // @[LVT_Mem.scala 74:14]
    end
    if (reset) begin // @[LVT_Mem.scala 71:27]
      r3_sel_reg <= 2'h0; // @[LVT_Mem.scala 71:27]
    end else begin
      r3_sel_reg <= LVT_r3_sel_reg_MPORT_data; // @[LVT_Mem.scala 75:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    LVT[initvar] = _RAND_0[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  r1_sel_reg = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  r2_sel_reg = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  r3_sel_reg = _RAND_3[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PRF(
  input         clock,
  input         reset,
  input  [5:0]  w1_addr,
  input  [63:0] w1_data,
  input         w1_en,
  input  [5:0]  w2_addr,
  input  [63:0] w2_data,
  input         w2_en,
  input  [5:0]  w3_addr,
  input  [63:0] w3_data,
  input         w3_en,
  input  [5:0]  w4_addr,
  input  [63:0] w4_data,
  input         w4_en,
  input         execRead_valid,
  input  [31:0] execRead_instruction,
  input  [4:0]  execRead_branchmask,
  input  [5:0]  execRead_rs1Addr,
  input  [5:0]  execRead_rs2Addr,
  input  [5:0]  execRead_robAddr,
  input  [5:0]  execRead_prfDest,
  output        toExec_valid,
  output [31:0] toExec_instruction,
  output [4:0]  toExec_branchmask,
  output [5:0]  toExec_rs1Addr,
  output [63:0] toExec_rs1Data,
  output [5:0]  toExec_rs2Addr,
  output [63:0] toExec_rs2Data,
  output [5:0]  toExec_robAddr,
  output [5:0]  toExec_prfDest,
  input         fromStore_valid,
  input  [5:0]  fromStore_rs2Addr,
  output        toStore_valid,
  output [63:0] toStore_rs2Data,
  input         branchCheck_pass,
  input  [4:0]  branchCheck_branchmask,
  input         branchCheck_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  prf_clock; // @[PRF.scala 73:19]
  wire  prf_reset; // @[PRF.scala 73:19]
  wire [5:0] prf_io_R1_addr; // @[PRF.scala 73:19]
  wire [63:0] prf_io_R1_data; // @[PRF.scala 73:19]
  wire  prf_io_R1_en; // @[PRF.scala 73:19]
  wire [5:0] prf_io_R2_addr; // @[PRF.scala 73:19]
  wire [63:0] prf_io_R2_data; // @[PRF.scala 73:19]
  wire  prf_io_R2_en; // @[PRF.scala 73:19]
  wire [5:0] prf_io_R3_addr; // @[PRF.scala 73:19]
  wire [63:0] prf_io_R3_data; // @[PRF.scala 73:19]
  wire  prf_io_R3_en; // @[PRF.scala 73:19]
  wire [5:0] prf_io_W1_addr; // @[PRF.scala 73:19]
  wire [63:0] prf_io_W1_data; // @[PRF.scala 73:19]
  wire  prf_io_W1_en; // @[PRF.scala 73:19]
  wire [5:0] prf_io_W2_addr; // @[PRF.scala 73:19]
  wire [63:0] prf_io_W2_data; // @[PRF.scala 73:19]
  wire  prf_io_W2_en; // @[PRF.scala 73:19]
  wire [5:0] prf_io_W3_addr; // @[PRF.scala 73:19]
  wire [63:0] prf_io_W3_data; // @[PRF.scala 73:19]
  wire  prf_io_W3_en; // @[PRF.scala 73:19]
  wire [5:0] prf_io_W4_addr; // @[PRF.scala 73:19]
  wire [63:0] prf_io_W4_data; // @[PRF.scala 73:19]
  wire  prf_io_W4_en; // @[PRF.scala 73:19]
  reg [5:0] toExec_robAddr_REG; // @[PRF.scala 82:28]
  reg [5:0] toExec_rs1Addr_REG; // @[PRF.scala 83:28]
  reg [5:0] toExec_rs2Addr_REG; // @[PRF.scala 84:28]
  reg [31:0] toExec_instruction_REG; // @[PRF.scala 85:32]
  reg [5:0] toExec_prfDest_REG; // @[PRF.scala 87:28]
  reg  toExec_valid_; // @[PRF.scala 104:29]
  reg [4:0] toExec_mask; // @[PRF.scala 107:28]
  wire [4:0] _T = branchCheck_branchmask & execRead_branchmask; // @[PRF.scala 115:36]
  wire [4:0] _toExec_mask_T = branchCheck_branchmask ^ execRead_branchmask; // @[PRF.scala 116:47]
  reg  toStore_valid_REG_1; // @[PRF.scala 140:27]
  LVT_Mem prf ( // @[PRF.scala 73:19]
    .clock(prf_clock),
    .reset(prf_reset),
    .io_R1_addr(prf_io_R1_addr),
    .io_R1_data(prf_io_R1_data),
    .io_R1_en(prf_io_R1_en),
    .io_R2_addr(prf_io_R2_addr),
    .io_R2_data(prf_io_R2_data),
    .io_R2_en(prf_io_R2_en),
    .io_R3_addr(prf_io_R3_addr),
    .io_R3_data(prf_io_R3_data),
    .io_R3_en(prf_io_R3_en),
    .io_W1_addr(prf_io_W1_addr),
    .io_W1_data(prf_io_W1_data),
    .io_W1_en(prf_io_W1_en),
    .io_W2_addr(prf_io_W2_addr),
    .io_W2_data(prf_io_W2_data),
    .io_W2_en(prf_io_W2_en),
    .io_W3_addr(prf_io_W3_addr),
    .io_W3_data(prf_io_W3_data),
    .io_W3_en(prf_io_W3_en),
    .io_W4_addr(prf_io_W4_addr),
    .io_W4_data(prf_io_W4_data),
    .io_W4_en(prf_io_W4_en)
  );
  assign toExec_valid = toExec_valid_; // @[PRF.scala 136:16]
  assign toExec_instruction = toExec_instruction_REG; // @[PRF.scala 85:22]
  assign toExec_branchmask = toExec_mask; // @[PRF.scala 137:21]
  assign toExec_rs1Addr = toExec_rs1Addr_REG; // @[PRF.scala 83:18]
  assign toExec_rs1Data = prf_io_R1_data; // @[PRF.scala 93:18]
  assign toExec_rs2Addr = toExec_rs2Addr_REG; // @[PRF.scala 84:18]
  assign toExec_rs2Data = prf_io_R2_data; // @[PRF.scala 97:18]
  assign toExec_robAddr = toExec_robAddr_REG; // @[PRF.scala 82:18]
  assign toExec_prfDest = toExec_prfDest_REG; // @[PRF.scala 87:18]
  assign toStore_valid = toStore_valid_REG_1; // @[PRF.scala 140:17]
  assign toStore_rs2Data = prf_io_R3_data; // @[PRF.scala 101:19]
  assign prf_clock = clock;
  assign prf_reset = reset;
  assign prf_io_R1_addr = execRead_rs1Addr; // @[PRF.scala 92:18]
  assign prf_io_R1_en = execRead_valid; // @[PRF.scala 91:16]
  assign prf_io_R2_addr = execRead_rs2Addr; // @[PRF.scala 96:18]
  assign prf_io_R2_en = execRead_valid; // @[PRF.scala 95:16]
  assign prf_io_R3_addr = fromStore_rs2Addr; // @[PRF.scala 100:18]
  assign prf_io_R3_en = fromStore_valid; // @[PRF.scala 99:16]
  assign prf_io_W1_addr = w1_addr; // @[PRF.scala 76:13]
  assign prf_io_W1_data = w1_data; // @[PRF.scala 76:13]
  assign prf_io_W1_en = w1_en; // @[PRF.scala 76:13]
  assign prf_io_W2_addr = w2_addr; // @[PRF.scala 77:13]
  assign prf_io_W2_data = w2_data; // @[PRF.scala 77:13]
  assign prf_io_W2_en = w2_en; // @[PRF.scala 77:13]
  assign prf_io_W3_addr = w3_addr; // @[PRF.scala 78:13]
  assign prf_io_W3_data = w3_data; // @[PRF.scala 78:13]
  assign prf_io_W3_en = w3_en; // @[PRF.scala 78:13]
  assign prf_io_W4_addr = w4_addr; // @[PRF.scala 79:13]
  assign prf_io_W4_data = w4_data; // @[PRF.scala 79:13]
  assign prf_io_W4_en = w4_en; // @[PRF.scala 79:13]
  always @(posedge clock) begin
    toExec_robAddr_REG <= execRead_robAddr; // @[PRF.scala 82:28]
    toExec_rs1Addr_REG <= execRead_rs1Addr; // @[PRF.scala 83:28]
    toExec_rs2Addr_REG <= execRead_rs2Addr; // @[PRF.scala 84:28]
    toExec_instruction_REG <= execRead_instruction; // @[PRF.scala 85:32]
    toExec_prfDest_REG <= execRead_prfDest; // @[PRF.scala 87:28]
    if (reset) begin // @[PRF.scala 104:29]
      toExec_valid_ <= 1'h0; // @[PRF.scala 104:29]
    end else if (branchCheck_valid) begin // @[PRF.scala 110:27]
      if (branchCheck_pass) begin // @[PRF.scala 112:28]
        toExec_valid_ <= execRead_valid; // @[PRF.scala 113:20]
      end else begin
        toExec_valid_ <= _T == 5'h0 & execRead_valid; // @[PRF.scala 122:20]
      end
    end else begin
      toExec_valid_ <= execRead_valid; // @[PRF.scala 129:18]
    end
    if (reset) begin // @[PRF.scala 107:28]
      toExec_mask <= 5'h0; // @[PRF.scala 107:28]
    end else if (branchCheck_valid) begin // @[PRF.scala 110:27]
      if (branchCheck_pass) begin // @[PRF.scala 112:28]
        if (|_T) begin // @[PRF.scala 115:64]
          toExec_mask <= _toExec_mask_T; // @[PRF.scala 116:21]
        end else begin
          toExec_mask <= execRead_branchmask; // @[PRF.scala 114:19]
        end
      end else begin
        toExec_mask <= execRead_branchmask; // @[PRF.scala 123:19]
      end
    end else begin
      toExec_mask <= execRead_branchmask; // @[PRF.scala 130:17]
    end
    if (reset) begin // @[PRF.scala 140:27]
      toStore_valid_REG_1 <= 1'h0; // @[PRF.scala 140:27]
    end else begin
      toStore_valid_REG_1 <= fromStore_valid; // @[PRF.scala 140:27]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  toExec_robAddr_REG = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  toExec_rs1Addr_REG = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  toExec_rs2Addr_REG = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  toExec_instruction_REG = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  toExec_prfDest_REG = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  toExec_valid_ = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  toExec_mask = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  toStore_valid_REG_1 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module soc1_Anon(
  input         clock,
  input         reset,
  output [31:0] iPort_ARADDR,
  output        iPort_ARVALID,
  input         iPort_ARREADY,
  input  [63:0] iPort_RDATA,
  input         iPort_RLAST,
  input         iPort_RVALID,
  output        iPort_RREADY,
  output        debug_probe_arvalid_internal,
  output        debug_probe_cacheMissed,
  output        debug_probe_rready_signal,
  output        debug_probe_cacheFill_valid,
  output        debug_probe_axi_arvalid,
  output        debug_probe_axi_arready,
  output        debug_probe_req_valid,
  output [63:0] debug_probe_req_pc,
  output        fdbg_probe_redirect_bit,
  output        fdbg_probe_fifo_enq_ready,
  output        fdbg_probe_is_fence,
  output        fdbg_probe_handle_fence,
  output [31:0] dPort_AWADDR,
  output        dPort_AWVALID,
  input         dPort_AWREADY,
  output [63:0] dPort_WDATA,
  output        dPort_WLAST,
  output        dPort_WVALID,
  input         dPort_WREADY,
  input  [1:0]  dPort_BRESP,
  input         dPort_BVALID,
  output        dPort_BREADY,
  output [31:0] dPort_ARADDR,
  output        dPort_ARVALID,
  input         dPort_ARREADY,
  input  [63:0] dPort_RDATA,
  input         dPort_RLAST,
  input         dPort_RVALID,
  output        dPort_RREADY,
  output [2:0]  dPort_AWSNOOP,
  output [3:0]  dPort_ARSNOOP,
  input  [3:0]  dPort_RRESP,
  input         dPort_ACVALID,
  output        dPort_ACREADY,
  input  [31:0] dPort_ACADDR,
  input  [3:0]  dPort_ACSNOOP,
  output        dPort_CRVALID,
  input         dPort_CRREADY,
  output [4:0]  dPort_CRRESP,
  output        dPort_CDVALID,
  input         dPort_CDREADY,
  output [63:0] dPort_CDDATA,
  output        dPort_CDLAST,
  output [31:0] peripheral_AWADDR,
  output [7:0]  peripheral_AWLEN,
  output [2:0]  peripheral_AWSIZE,
  output [1:0]  peripheral_AWBURST,
  output [2:0]  peripheral_AWPROT,
  output        peripheral_AWVALID,
  input         peripheral_AWREADY,
  output [31:0] peripheral_WDATA,
  output [3:0]  peripheral_WSTRB,
  output        peripheral_WLAST,
  output        peripheral_WVALID,
  input         peripheral_WREADY,
  input         peripheral_BID,
  input  [1:0]  peripheral_BRESP,
  input         peripheral_BVALID,
  output        peripheral_BREADY,
  output [31:0] peripheral_ARADDR,
  output [7:0]  peripheral_ARLEN,
  output [2:0]  peripheral_ARSIZE,
  output [1:0]  peripheral_ARBURST,
  output [2:0]  peripheral_ARPROT,
  output        peripheral_ARVALID,
  input         peripheral_ARREADY,
  input         peripheral_RID,
  input  [31:0] peripheral_RDATA,
  input  [1:0]  peripheral_RRESP,
  input         peripheral_RLAST,
  input         peripheral_RVALID,
  output        peripheral_RREADY,
  output        core_sample0,
  output        core_sample1,
  input         MTIP
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [95:0] _RAND_47;
  reg [95:0] _RAND_48;
  reg [95:0] _RAND_49;
  reg [95:0] _RAND_50;
  reg [95:0] _RAND_51;
  reg [95:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [95:0] _RAND_62;
  reg [95:0] _RAND_63;
  reg [95:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
`endif // RANDOMIZE_REG_INIT
  wire  icache_clock; // @[core.scala 28:22]
  wire  icache_reset; // @[core.scala 28:22]
  wire  icache_fromFetch_req_ready; // @[core.scala 28:22]
  wire  icache_fromFetch_req_valid; // @[core.scala 28:22]
  wire [63:0] icache_fromFetch_req_bits; // @[core.scala 28:22]
  wire  icache_fromFetch_resp_ready; // @[core.scala 28:22]
  wire  icache_fromFetch_resp_valid; // @[core.scala 28:22]
  wire [31:0] icache_fromFetch_resp_bits; // @[core.scala 28:22]
  wire  icache_updateAllCachelines_ready; // @[core.scala 28:22]
  wire  icache_updateAllCachelines_fired; // @[core.scala 28:22]
  wire  icache_cachelinesUpdatesResp_ready; // @[core.scala 28:22]
  wire  icache_cachelinesUpdatesResp_fired; // @[core.scala 28:22]
  wire [31:0] icache_lowLevelMem_ARADDR; // @[core.scala 28:22]
  wire  icache_lowLevelMem_ARVALID; // @[core.scala 28:22]
  wire  icache_lowLevelMem_ARREADY; // @[core.scala 28:22]
  wire [63:0] icache_lowLevelMem_RDATA; // @[core.scala 28:22]
  wire  icache_lowLevelMem_RLAST; // @[core.scala 28:22]
  wire  icache_lowLevelMem_RVALID; // @[core.scala 28:22]
  wire  icache_lowLevelMem_RREADY; // @[core.scala 28:22]
  wire  icache_debug_probe_arvalid_internal; // @[core.scala 28:22]
  wire  icache_debug_probe_cacheMissed; // @[core.scala 28:22]
  wire  icache_debug_probe_rready_signal; // @[core.scala 28:22]
  wire  icache_debug_probe_cacheFill_valid; // @[core.scala 28:22]
  wire  icache_debug_probe_axi_arvalid; // @[core.scala 28:22]
  wire  icache_debug_probe_axi_arready; // @[core.scala 28:22]
  wire  icache_debug_probe_req_valid; // @[core.scala 28:22]
  wire [63:0] icache_debug_probe_req_pc; // @[core.scala 28:22]
  wire  fetch_clock; // @[core.scala 42:21]
  wire  fetch_reset; // @[core.scala 42:21]
  wire  fetch_cache_req_ready; // @[core.scala 42:21]
  wire  fetch_cache_req_valid; // @[core.scala 42:21]
  wire [63:0] fetch_cache_req_bits; // @[core.scala 42:21]
  wire  fetch_cache_resp_ready; // @[core.scala 42:21]
  wire  fetch_cache_resp_valid; // @[core.scala 42:21]
  wire [31:0] fetch_cache_resp_bits; // @[core.scala 42:21]
  wire  fetch_toDecode_ready; // @[core.scala 42:21]
  wire  fetch_toDecode_fired; // @[core.scala 42:21]
  wire [63:0] fetch_toDecode_pc; // @[core.scala 42:21]
  wire [31:0] fetch_toDecode_instruction; // @[core.scala 42:21]
  wire  fetch_toDecode_expected_valid; // @[core.scala 42:21]
  wire [63:0] fetch_toDecode_expected_pc; // @[core.scala 42:21]
  wire  fetch_toDecode_expected_coherency; // @[core.scala 42:21]
  wire  fetch_branchRes_fired; // @[core.scala 42:21]
  wire  fetch_branchRes_branchTaken; // @[core.scala 42:21]
  wire [63:0] fetch_branchRes_pc; // @[core.scala 42:21]
  wire [63:0] fetch_branchRes_pcAfterBrnach; // @[core.scala 42:21]
  wire  fetch_carryOutFence_ready; // @[core.scala 42:21]
  wire  fetch_carryOutFence_fired; // @[core.scala 42:21]
  wire  fetch_updateAllCachelines_ready; // @[core.scala 42:21]
  wire  fetch_updateAllCachelines_fired; // @[core.scala 42:21]
  wire  fetch_cachelinesUpdatesResp_ready; // @[core.scala 42:21]
  wire  fetch_cachelinesUpdatesResp_fired; // @[core.scala 42:21]
  wire  fetch_fdbg_probe_redirect_bit; // @[core.scala 42:21]
  wire  fetch_fdbg_probe_fifo_enq_ready; // @[core.scala 42:21]
  wire  fetch_fdbg_probe_is_fence; // @[core.scala 42:21]
  wire  fetch_fdbg_probe_handle_fence; // @[core.scala 42:21]
  wire  decode_clock; // @[core.scala 57:22]
  wire  decode_reset; // @[core.scala 57:22]
  wire  decode_fromFetch_ready; // @[core.scala 57:22]
  wire  decode_fromFetch_fired; // @[core.scala 57:22]
  wire [63:0] decode_fromFetch_pc; // @[core.scala 57:22]
  wire [31:0] decode_fromFetch_instruction; // @[core.scala 57:22]
  wire  decode_fromFetch_expected_valid; // @[core.scala 57:22]
  wire [63:0] decode_fromFetch_expected_pc; // @[core.scala 57:22]
  wire  decode_fromFetch_expected_coherency; // @[core.scala 57:22]
  wire  decode_toExec_ready; // @[core.scala 57:22]
  wire  decode_toExec_fired; // @[core.scala 57:22]
  wire [31:0] decode_toExec_instruction; // @[core.scala 57:22]
  wire [63:0] decode_toExec_pc; // @[core.scala 57:22]
  wire [5:0] decode_toExec_PRFDest; // @[core.scala 57:22]
  wire [5:0] decode_toExec_rs1Addr; // @[core.scala 57:22]
  wire  decode_toExec_rs1Ready; // @[core.scala 57:22]
  wire [5:0] decode_toExec_rs2Addr; // @[core.scala 57:22]
  wire  decode_toExec_rs2Ready; // @[core.scala 57:22]
  wire [4:0] decode_toExec_branchMask; // @[core.scala 57:22]
  wire  decode_writeBackResult_fired; // @[core.scala 57:22]
  wire [31:0] decode_writeBackResult_instruction; // @[core.scala 57:22]
  wire [4:0] decode_writeBackResult_rdAddr; // @[core.scala 57:22]
  wire [5:0] decode_writeBackResult_PRFDest; // @[core.scala 57:22]
  wire [63:0] decode_writeBackResult_data; // @[core.scala 57:22]
  wire [5:0] decode_writeAddrPRF_exec1Addr; // @[core.scala 57:22]
  wire [5:0] decode_writeAddrPRF_exec2Addr; // @[core.scala 57:22]
  wire [5:0] decode_writeAddrPRF_exec3Addr; // @[core.scala 57:22]
  wire  decode_writeAddrPRF_exec1Valid; // @[core.scala 57:22]
  wire  decode_writeAddrPRF_exec2Valid; // @[core.scala 57:22]
  wire  decode_writeAddrPRF_exec3Valid; // @[core.scala 57:22]
  wire  decode_jumpAddrWrite_ready; // @[core.scala 57:22]
  wire  decode_jumpAddrWrite_fired; // @[core.scala 57:22]
  wire [5:0] decode_jumpAddrWrite_PRFDest; // @[core.scala 57:22]
  wire [63:0] decode_jumpAddrWrite_linkAddr; // @[core.scala 57:22]
  wire  decode_branchPCs_branchPCReady; // @[core.scala 57:22]
  wire [63:0] decode_branchPCs_branchPC; // @[core.scala 57:22]
  wire  decode_branchPCs_predictedPCReady; // @[core.scala 57:22]
  wire [63:0] decode_branchPCs_predictedPC; // @[core.scala 57:22]
  wire [4:0] decode_branchPCs_branchMask; // @[core.scala 57:22]
  wire  decode_branchEvalIn_fired; // @[core.scala 57:22]
  wire  decode_branchEvalIn_passFail; // @[core.scala 57:22]
  wire [4:0] decode_branchEvalIn_branchMask; // @[core.scala 57:22]
  wire [63:0] decode_branchEvalIn_targetPC; // @[core.scala 57:22]
  wire [63:0] decode_interruptedPC; // @[core.scala 57:22]
  wire  decode_canTakeInterrupt; // @[core.scala 57:22]
  wire  dataQueue_clock; // @[core.scala 73:25]
  wire  dataQueue_reset; // @[core.scala 73:25]
  wire  dataQueue_fromROB_readyNow; // @[core.scala 73:25]
  wire  dataQueue_fromBranch_passOrFail; // @[core.scala 73:25]
  wire [3:0] dataQueue_fromBranch_robAddr; // @[core.scala 73:25]
  wire  dataQueue_fromBranch_valid; // @[core.scala 73:25]
  wire  dataQueue_fromDecode_ready; // @[core.scala 73:25]
  wire  dataQueue_fromDecode_valid; // @[core.scala 73:25]
  wire [5:0] dataQueue_fromDecode_rs2Addr; // @[core.scala 73:25]
  wire [4:0] dataQueue_fromDecode_branchMask; // @[core.scala 73:25]
  wire  dataQueue_toPRF_valid; // @[core.scala 73:25]
  wire [5:0] dataQueue_toPRF_rs2Addr; // @[core.scala 73:25]
  wire  dataQueue_robMapUpdate_valid; // @[core.scala 73:25]
  wire [3:0] dataQueue_robMapUpdate_robAddr; // @[core.scala 73:25]
  wire  rob_clock; // @[core.scala 74:19]
  wire  rob_reset; // @[core.scala 74:19]
  wire  rob_allocate_ready; // @[core.scala 74:19]
  wire  rob_allocate_fired; // @[core.scala 74:19]
  wire [63:0] rob_allocate_pc; // @[core.scala 74:19]
  wire [31:0] rob_allocate_instruction; // @[core.scala 74:19]
  wire [5:0] rob_allocate_prfDest; // @[core.scala 74:19]
  wire [3:0] rob_allocate_robAddr; // @[core.scala 74:19]
  wire  rob_allocate_isReady; // @[core.scala 74:19]
  wire  rob_commit_ready; // @[core.scala 74:19]
  wire  rob_commit_fired; // @[core.scala 74:19]
  wire [5:0] rob_commit_prfDest; // @[core.scala 74:19]
  wire [63:0] rob_commit_pc; // @[core.scala 74:19]
  wire [31:0] rob_commit_instruction; // @[core.scala 74:19]
  wire  rob_commit_exceptionOccurred; // @[core.scala 74:19]
  wire [63:0] rob_commit_mtval; // @[core.scala 74:19]
  wire  rob_commit_isStore; // @[core.scala 74:19]
  wire  rob_commit_is_fence; // @[core.scala 74:19]
  wire [3:0] rob_commit_robAddr; // @[core.scala 74:19]
  wire  rob_branch_valid; // @[core.scala 74:19]
  wire  rob_branch_pass; // @[core.scala 74:19]
  wire [3:0] rob_branch_robAddr; // @[core.scala 74:19]
  wire [3:0] rob_execPorts_0_robAddr; // @[core.scala 74:19]
  wire [63:0] rob_execPorts_0_mtval; // @[core.scala 74:19]
  wire  rob_execPorts_0_valid; // @[core.scala 74:19]
  wire [3:0] rob_execPorts_1_robAddr; // @[core.scala 74:19]
  wire  rob_execPorts_1_valid; // @[core.scala 74:19]
  wire [3:0] rob_execPorts_2_robAddr; // @[core.scala 74:19]
  wire  rob_execPorts_2_valid; // @[core.scala 74:19]
  wire [3:0] rob_execPorts_3_robAddr; // @[core.scala 74:19]
  wire  rob_execPorts_3_valid; // @[core.scala 74:19]
  wire  scheduler_clock; // @[core.scala 75:25]
  wire  scheduler_reset; // @[core.scala 75:25]
  wire  scheduler_allocate_ready; // @[core.scala 75:25]
  wire  scheduler_allocate_fired; // @[core.scala 75:25]
  wire [31:0] scheduler_allocate_instruction; // @[core.scala 75:25]
  wire [4:0] scheduler_allocate_branchMask; // @[core.scala 75:25]
  wire  scheduler_allocate_rs1_ready; // @[core.scala 75:25]
  wire [5:0] scheduler_allocate_rs1_prfAddr; // @[core.scala 75:25]
  wire  scheduler_allocate_rs2_ready; // @[core.scala 75:25]
  wire [5:0] scheduler_allocate_rs2_prfAddr; // @[core.scala 75:25]
  wire [5:0] scheduler_allocate_prfDest; // @[core.scala 75:25]
  wire [3:0] scheduler_allocate_robAddr; // @[core.scala 75:25]
  wire  scheduler_release_ready; // @[core.scala 75:25]
  wire  scheduler_release_fired; // @[core.scala 75:25]
  wire [31:0] scheduler_release_instruction; // @[core.scala 75:25]
  wire [4:0] scheduler_release_branchMask; // @[core.scala 75:25]
  wire [5:0] scheduler_release_rs1prfAddr; // @[core.scala 75:25]
  wire [5:0] scheduler_release_rs2prfAddr; // @[core.scala 75:25]
  wire [5:0] scheduler_release_prfDest; // @[core.scala 75:25]
  wire [3:0] scheduler_release_robAddr; // @[core.scala 75:25]
  wire  scheduler_wakeUpExt_0_valid; // @[core.scala 75:25]
  wire [5:0] scheduler_wakeUpExt_0_prfAddr; // @[core.scala 75:25]
  wire  scheduler_wakeUpExt_1_valid; // @[core.scala 75:25]
  wire [5:0] scheduler_wakeUpExt_1_prfAddr; // @[core.scala 75:25]
  wire  scheduler_branchOps_valid; // @[core.scala 75:25]
  wire [4:0] scheduler_branchOps_branchMask; // @[core.scala 75:25]
  wire  scheduler_branchOps_passed; // @[core.scala 75:25]
  wire  scheduler_memoryReady; // @[core.scala 75:25]
  wire  scheduler_multuplyAndDivideReady; // @[core.scala 75:25]
  wire  scheduler_instrRetired_valid; // @[core.scala 75:25]
  wire [5:0] scheduler_instrRetired_prfAddr; // @[core.scala 75:25]
  wire  memAccess_clock; // @[core.scala 76:25]
  wire  memAccess_reset; // @[core.scala 76:25]
  wire  memAccess_request_valid; // @[core.scala 76:25]
  wire [31:0] memAccess_request_address; // @[core.scala 76:25]
  wire [31:0] memAccess_request_instruction; // @[core.scala 76:25]
  wire [4:0] memAccess_request_branchMask; // @[core.scala 76:25]
  wire [3:0] memAccess_request_robAddr; // @[core.scala 76:25]
  wire [5:0] memAccess_request_prfDest; // @[core.scala 76:25]
  wire [31:0] memAccess_dPort_AWADDR; // @[core.scala 76:25]
  wire  memAccess_dPort_AWVALID; // @[core.scala 76:25]
  wire  memAccess_dPort_AWREADY; // @[core.scala 76:25]
  wire [63:0] memAccess_dPort_WDATA; // @[core.scala 76:25]
  wire  memAccess_dPort_WLAST; // @[core.scala 76:25]
  wire  memAccess_dPort_WVALID; // @[core.scala 76:25]
  wire  memAccess_dPort_WREADY; // @[core.scala 76:25]
  wire [1:0] memAccess_dPort_BRESP; // @[core.scala 76:25]
  wire  memAccess_dPort_BVALID; // @[core.scala 76:25]
  wire  memAccess_dPort_BREADY; // @[core.scala 76:25]
  wire [31:0] memAccess_dPort_ARADDR; // @[core.scala 76:25]
  wire  memAccess_dPort_ARVALID; // @[core.scala 76:25]
  wire  memAccess_dPort_ARREADY; // @[core.scala 76:25]
  wire [63:0] memAccess_dPort_RDATA; // @[core.scala 76:25]
  wire  memAccess_dPort_RLAST; // @[core.scala 76:25]
  wire  memAccess_dPort_RVALID; // @[core.scala 76:25]
  wire  memAccess_dPort_RREADY; // @[core.scala 76:25]
  wire [2:0] memAccess_dPort_AWSNOOP; // @[core.scala 76:25]
  wire [3:0] memAccess_dPort_ARSNOOP; // @[core.scala 76:25]
  wire [3:0] memAccess_dPort_RRESP; // @[core.scala 76:25]
  wire  memAccess_dPort_ACVALID; // @[core.scala 76:25]
  wire  memAccess_dPort_ACREADY; // @[core.scala 76:25]
  wire [31:0] memAccess_dPort_ACADDR; // @[core.scala 76:25]
  wire [3:0] memAccess_dPort_ACSNOOP; // @[core.scala 76:25]
  wire  memAccess_dPort_CRVALID; // @[core.scala 76:25]
  wire  memAccess_dPort_CRREADY; // @[core.scala 76:25]
  wire [4:0] memAccess_dPort_CRRESP; // @[core.scala 76:25]
  wire  memAccess_dPort_CDVALID; // @[core.scala 76:25]
  wire  memAccess_dPort_CDREADY; // @[core.scala 76:25]
  wire [63:0] memAccess_dPort_CDDATA; // @[core.scala 76:25]
  wire  memAccess_dPort_CDLAST; // @[core.scala 76:25]
  wire [31:0] memAccess_peripheral_AWADDR; // @[core.scala 76:25]
  wire [7:0] memAccess_peripheral_AWLEN; // @[core.scala 76:25]
  wire [2:0] memAccess_peripheral_AWSIZE; // @[core.scala 76:25]
  wire [1:0] memAccess_peripheral_AWBURST; // @[core.scala 76:25]
  wire [2:0] memAccess_peripheral_AWPROT; // @[core.scala 76:25]
  wire  memAccess_peripheral_AWVALID; // @[core.scala 76:25]
  wire  memAccess_peripheral_AWREADY; // @[core.scala 76:25]
  wire [31:0] memAccess_peripheral_WDATA; // @[core.scala 76:25]
  wire [3:0] memAccess_peripheral_WSTRB; // @[core.scala 76:25]
  wire  memAccess_peripheral_WLAST; // @[core.scala 76:25]
  wire  memAccess_peripheral_WVALID; // @[core.scala 76:25]
  wire  memAccess_peripheral_WREADY; // @[core.scala 76:25]
  wire [1:0] memAccess_peripheral_BID; // @[core.scala 76:25]
  wire [1:0] memAccess_peripheral_BRESP; // @[core.scala 76:25]
  wire  memAccess_peripheral_BVALID; // @[core.scala 76:25]
  wire  memAccess_peripheral_BREADY; // @[core.scala 76:25]
  wire [31:0] memAccess_peripheral_ARADDR; // @[core.scala 76:25]
  wire [7:0] memAccess_peripheral_ARLEN; // @[core.scala 76:25]
  wire [2:0] memAccess_peripheral_ARSIZE; // @[core.scala 76:25]
  wire [1:0] memAccess_peripheral_ARBURST; // @[core.scala 76:25]
  wire [2:0] memAccess_peripheral_ARPROT; // @[core.scala 76:25]
  wire  memAccess_peripheral_ARVALID; // @[core.scala 76:25]
  wire  memAccess_peripheral_ARREADY; // @[core.scala 76:25]
  wire [1:0] memAccess_peripheral_RID; // @[core.scala 76:25]
  wire [31:0] memAccess_peripheral_RDATA; // @[core.scala 76:25]
  wire [1:0] memAccess_peripheral_RRESP; // @[core.scala 76:25]
  wire  memAccess_peripheral_RLAST; // @[core.scala 76:25]
  wire  memAccess_peripheral_RVALID; // @[core.scala 76:25]
  wire  memAccess_peripheral_RREADY; // @[core.scala 76:25]
  wire  memAccess_responseOut_valid; // @[core.scala 76:25]
  wire [5:0] memAccess_responseOut_prfDest; // @[core.scala 76:25]
  wire [3:0] memAccess_responseOut_robAddr; // @[core.scala 76:25]
  wire [63:0] memAccess_responseOut_result; // @[core.scala 76:25]
  wire [31:0] memAccess_responseOut_instruction; // @[core.scala 76:25]
  wire  memAccess_canAllocate; // @[core.scala 76:25]
  wire  memAccess_writeDataIn_valid; // @[core.scala 76:25]
  wire [63:0] memAccess_writeDataIn_data; // @[core.scala 76:25]
  wire  memAccess_initiateFence; // @[core.scala 76:25]
  wire  memAccess_fenceInstructions_ready; // @[core.scala 76:25]
  wire  memAccess_fenceInstructions_fired; // @[core.scala 76:25]
  wire  memAccess_writeCommit_ready; // @[core.scala 76:25]
  wire  memAccess_writeCommit_fired; // @[core.scala 76:25]
  wire  memAccess_writeInstructionCommit_ready; // @[core.scala 76:25]
  wire  memAccess_writeInstructionCommit_fired; // @[core.scala 76:25]
  wire  memAccess_branchOps_valid; // @[core.scala 76:25]
  wire [4:0] memAccess_branchOps_branchMask; // @[core.scala 76:25]
  wire  memAccess_branchOps_passed; // @[core.scala 76:25]
  wire  memAccess_loadCommit_ready; // @[core.scala 76:25]
  wire  memAccess_loadCommit_valid; // @[core.scala 76:25]
  wire  memAccess_loadCommit_state; // @[core.scala 76:25]
  wire  prf_clock; // @[core.scala 143:19]
  wire  prf_reset; // @[core.scala 143:19]
  wire [5:0] prf_w1_addr; // @[core.scala 143:19]
  wire [63:0] prf_w1_data; // @[core.scala 143:19]
  wire  prf_w1_en; // @[core.scala 143:19]
  wire [5:0] prf_w2_addr; // @[core.scala 143:19]
  wire [63:0] prf_w2_data; // @[core.scala 143:19]
  wire  prf_w2_en; // @[core.scala 143:19]
  wire [5:0] prf_w3_addr; // @[core.scala 143:19]
  wire [63:0] prf_w3_data; // @[core.scala 143:19]
  wire  prf_w3_en; // @[core.scala 143:19]
  wire [5:0] prf_w4_addr; // @[core.scala 143:19]
  wire [63:0] prf_w4_data; // @[core.scala 143:19]
  wire  prf_w4_en; // @[core.scala 143:19]
  wire  prf_execRead_valid; // @[core.scala 143:19]
  wire [31:0] prf_execRead_instruction; // @[core.scala 143:19]
  wire [4:0] prf_execRead_branchmask; // @[core.scala 143:19]
  wire [5:0] prf_execRead_rs1Addr; // @[core.scala 143:19]
  wire [5:0] prf_execRead_rs2Addr; // @[core.scala 143:19]
  wire [5:0] prf_execRead_robAddr; // @[core.scala 143:19]
  wire [5:0] prf_execRead_prfDest; // @[core.scala 143:19]
  wire  prf_toExec_valid; // @[core.scala 143:19]
  wire [31:0] prf_toExec_instruction; // @[core.scala 143:19]
  wire [4:0] prf_toExec_branchmask; // @[core.scala 143:19]
  wire [5:0] prf_toExec_rs1Addr; // @[core.scala 143:19]
  wire [63:0] prf_toExec_rs1Data; // @[core.scala 143:19]
  wire [5:0] prf_toExec_rs2Addr; // @[core.scala 143:19]
  wire [63:0] prf_toExec_rs2Data; // @[core.scala 143:19]
  wire [5:0] prf_toExec_robAddr; // @[core.scala 143:19]
  wire [5:0] prf_toExec_prfDest; // @[core.scala 143:19]
  wire  prf_fromStore_valid; // @[core.scala 143:19]
  wire [5:0] prf_fromStore_rs2Addr; // @[core.scala 143:19]
  wire  prf_toStore_valid; // @[core.scala 143:19]
  wire [63:0] prf_toStore_rs2Data; // @[core.scala 143:19]
  wire  prf_branchCheck_pass; // @[core.scala 143:19]
  wire [4:0] prf_branchCheck_branchmask; // @[core.scala 143:19]
  wire  prf_branchCheck_valid; // @[core.scala 143:19]
  wire  _fetch_toDecode_fired_T_3 = ~decode_fromFetch_expected_valid | decode_fromFetch_expected_pc == fetch_toDecode_pc
    ; // @[core.scala 66:40]
  wire  instructionDecodedReady = 5'h3 == decode_toExec_instruction[6:2] | 5'h5 == decode_toExec_instruction[6:2] | 5'hd
     == decode_toExec_instruction[6:2]; // @[core.scala 101:125]
  wire [6:0] _scheduler_allocate_rs2_ready_T_1 = decode_toExec_instruction[6:0] & 7'h77; // @[core.scala 114:72]
  wire  _GEN_0 = instructionDecodedReady ? 1'h0 : decode_toExec_ready & rob_allocate_ready & scheduler_allocate_ready &
    (decode_toExec_instruction[6:4] != 3'h2 | dataQueue_fromDecode_ready); // @[core.scala 123:{33,60} 103:7]
  reg [4:0] branchEvals_branchMask; // @[core.scala 534:28]
  wire [4:0] _scheduler_allocate_branchMask_T = decode_toExec_branchMask ^ branchEvals_branchMask; // @[core.scala 125:62]
  reg  branchEvals_passed; // @[core.scala 534:28]
  wire  _T = ~branchEvals_passed; // @[core.scala 127:9]
  wire  _GEN_1 = ~branchEvals_passed ? 1'h0 : _GEN_0; // @[core.scala 127:28 128:30]
  wire  _GEN_2 = ~branchEvals_passed ? 1'h0 : decode_toExec_ready & rob_allocate_ready & scheduler_allocate_ready & (
    decode_toExec_instruction[6:4] != 3'h2 | dataQueue_fromDecode_ready); // @[core.scala 127:28 129:24 103:7]
  wire  _GEN_3 = ~branchEvals_passed ? 1'h0 : scheduler_allocate_fired & decode_toExec_instruction[6:4] == 3'h2; // @[core.scala 127:28 122:30 130:32]
  reg  branchEvals_valid; // @[core.scala 534:28]
  wire [5:0] wakeUps_0_prfAddr = scheduler_instrRetired_prfAddr; // @[core.scala 803:20 95:21]
  wire  _GEN_9 = decode_toExec_rs1Addr == wakeUps_0_prfAddr | decode_toExec_rs1Ready; // @[core.scala 112:32 136:{55,86}]
  wire  _GEN_10 = decode_toExec_rs2Addr == wakeUps_0_prfAddr | (7'h13 == _scheduler_allocate_rs2_ready_T_1 |
    decode_toExec_rs2Ready); // @[core.scala 114:32 137:{55,86}]
  wire  wakeUps_0_valid = scheduler_instrRetired_valid; // @[core.scala 804:18 95:21]
  wire  _GEN_11 = wakeUps_0_valid ? _GEN_9 : decode_toExec_rs1Ready; // @[core.scala 135:24 112:32]
  wire  _GEN_12 = wakeUps_0_valid ? _GEN_10 : 7'h13 == _scheduler_allocate_rs2_ready_T_1 | decode_toExec_rs2Ready; // @[core.scala 135:24 114:32]
  wire [5:0] wakeUps_1_prfAddr = memAccess_responseOut_prfDest; // @[core.scala 803:20 95:21]
  wire  _GEN_13 = decode_toExec_rs1Addr == wakeUps_1_prfAddr | _GEN_11; // @[core.scala 136:{55,86}]
  wire  _GEN_14 = decode_toExec_rs2Addr == wakeUps_1_prfAddr | _GEN_12; // @[core.scala 137:{55,86}]
  wire  _T_181 = |memAccess_responseOut_instruction[11:7]; // @[core.scala 798:77]
  wire  wakeUps_1_valid = memAccess_responseOut_valid & |memAccess_responseOut_instruction[11:7]; // @[core.scala 798:33]
  wire  _GEN_15 = wakeUps_1_valid ? _GEN_13 : _GEN_11; // @[core.scala 135:24]
  wire  _GEN_16 = wakeUps_1_valid ? _GEN_14 : _GEN_12; // @[core.scala 135:24]
  reg [5:0] extnMResponse_prfDest; // @[core.scala 235:30]
  wire  _GEN_17 = decode_toExec_rs1Addr == extnMResponse_prfDest | _GEN_15; // @[core.scala 136:{55,86}]
  wire  _GEN_18 = decode_toExec_rs2Addr == extnMResponse_prfDest | _GEN_16; // @[core.scala 137:{55,86}]
  reg  extnMResponse_valid; // @[core.scala 235:30]
  reg [31:0] extnResponseInstruction; // @[core.scala 374:36]
  wire  _T_184 = |extnResponseInstruction[11:7]; // @[core.scala 799:59]
  wire  wakeUps_2_valid = extnMResponse_valid & |extnResponseInstruction[11:7]; // @[core.scala 799:25]
  reg  mExtensionReady; // @[core.scala 141:32]
  wire [3:0] _scheduler_release_fired_T_2 = {scheduler_release_instruction[25],scheduler_release_instruction[6:4]}; // @[Cat.scala 33:92]
  wire  _scheduler_release_fired_T_5 = ~(_scheduler_release_fired_T_2 == 4'hb) | mExtensionReady; // @[core.scala 147:99]
  wire  _GEN_21 = scheduler_release_instruction[1:0] == 2'h0 ? 1'h0 : scheduler_release_fired; // @[core.scala 154:22 156:{57,78}]
  reg  addressGenerationInput_valid; // @[core.scala 164:39]
  reg [63:0] addressGenerationInput_rs1; // @[core.scala 164:39]
  reg [31:0] addressGenerationInput_instruction; // @[core.scala 164:39]
  reg [5:0] addressGenerationInput_prfDest; // @[core.scala 164:39]
  reg [3:0] addressGenerationInput_robAddr; // @[core.scala 164:39]
  reg [4:0] addressGenerationInput_branchMask; // @[core.scala 164:39]
  wire [4:0] _T_9 = prf_toExec_branchmask & branchEvals_branchMask; // @[core.scala 181:33]
  wire  _T_10 = |_T_9; // @[core.scala 181:57]
  wire [4:0] _addressGenerationInput_branchMask_T = prf_toExec_branchmask ^ branchEvals_branchMask; // @[core.scala 182:66]
  wire [4:0] _GEN_22 = |_T_9 ? _addressGenerationInput_branchMask_T : prf_toExec_branchmask; // @[core.scala 178:37 181:62 182:41]
  wire  _T_14 = _T & _T_10; // @[core.scala 184:28]
  wire [4:0] _GEN_24 = branchEvals_valid ? _GEN_22 : prf_toExec_branchmask; // @[core.scala 180:25 178:37]
  reg  memoryRequest_valid; // @[core.scala 187:30]
  reg [31:0] memoryRequest_address; // @[core.scala 187:30]
  reg [31:0] memoryRequest_instruction; // @[core.scala 187:30]
  reg [4:0] memoryRequest_branchMask; // @[core.scala 187:30]
  reg [3:0] memoryRequest_robAddr; // @[core.scala 187:30]
  reg [5:0] memoryRequest_prfDest; // @[core.scala 187:30]
  wire [51:0] _memoryRequest_address_T_2 = addressGenerationInput_instruction[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _memoryRequest_address_T_4 = {_memoryRequest_address_T_2,addressGenerationInput_instruction[31:20]}; // @[Cat.scala 33:92]
  wire [63:0] _memoryRequest_address_T_10 = {_memoryRequest_address_T_2,addressGenerationInput_instruction[31:25],
    addressGenerationInput_instruction[11:7]}; // @[Cat.scala 33:92]
  wire [1:0] _memoryRequest_address_T_13 = {addressGenerationInput_instruction[3],addressGenerationInput_instruction[5]}
    ; // @[Cat.scala 33:92]
  wire [63:0] _GEN_27 = 2'h1 == _memoryRequest_address_T_13 ? _memoryRequest_address_T_10 : _memoryRequest_address_T_4; // @[core.scala 188:{55,55}]
  wire [63:0] _GEN_28 = 2'h2 == _memoryRequest_address_T_13 ? 64'h0 : _GEN_27; // @[core.scala 188:{55,55}]
  wire [63:0] _GEN_29 = 2'h3 == _memoryRequest_address_T_13 ? 64'h0 : _GEN_28; // @[core.scala 188:{55,55}]
  wire [63:0] _memoryRequest_address_T_15 = addressGenerationInput_rs1 + _GEN_29; // @[core.scala 188:55]
  wire [4:0] _T_15 = addressGenerationInput_branchMask & branchEvals_branchMask; // @[core.scala 200:45]
  wire  _T_16 = |_T_15; // @[core.scala 200:69]
  wire [4:0] _memoryRequest_branchMask_T = addressGenerationInput_branchMask ^ branchEvals_branchMask; // @[core.scala 201:69]
  reg  singleCycleArithmeticRequest_valid; // @[core.scala 209:45]
  reg [63:0] singleCycleArithmeticRequest_rs1; // @[core.scala 209:45]
  reg [63:0] singleCycleArithmeticRequest_rs2; // @[core.scala 209:45]
  reg [31:0] singleCycleArithmeticRequest_instruction; // @[core.scala 209:45]
  reg [5:0] singleCycleArithmeticRequest_prfDest; // @[core.scala 209:45]
  reg [3:0] singleCycleArithmeticRequest_robAddr; // @[core.scala 209:45]
  reg [4:0] singleCycleArithmeticRequest_branchMask; // @[core.scala 209:45]
  reg  singleCycleArithmeticResponse_valid; // @[core.scala 219:46]
  reg [63:0] singleCycleArithmeticResponse_result; // @[core.scala 219:46]
  reg [5:0] singleCycleArithmeticResponse_prfDest; // @[core.scala 219:46]
  reg [3:0] singleCycleArithmeticResponse_robAddr; // @[core.scala 219:46]
  reg  extnMRequest_valid; // @[core.scala 226:29]
  reg [63:0] extnMRequest_rs1; // @[core.scala 226:29]
  reg [63:0] extnMRequest_rs2; // @[core.scala 226:29]
  reg [31:0] extnMRequest_instruction; // @[core.scala 226:29]
  reg [5:0] extnMRequest_prfDest; // @[core.scala 226:29]
  reg [3:0] extnMRequest_robAddr; // @[core.scala 226:29]
  reg [4:0] extnMRequest_branchMask; // @[core.scala 226:29]
  reg  extnMServicing_valid; // @[core.scala 228:31]
  reg [31:0] extnMServicing_instruction; // @[core.scala 228:31]
  reg [5:0] extnMServicing_prfDest; // @[core.scala 228:31]
  reg [3:0] extnMServicing_robAddr; // @[core.scala 228:31]
  reg [4:0] extnMServicing_branchMask; // @[core.scala 228:31]
  reg  extnMPartialServicing_valid; // @[core.scala 229:38]
  reg [31:0] extnMPartialServicing_instruction; // @[core.scala 229:38]
  reg [5:0] extnMPartialServicing_prfDest; // @[core.scala 229:38]
  reg [3:0] extnMPartialServicing_robAddr; // @[core.scala 229:38]
  reg [4:0] extnMPartialServicing_branchMask; // @[core.scala 229:38]
  reg [95:0] muls_0; // @[core.scala 230:17]
  reg [95:0] muls_1; // @[core.scala 230:17]
  reg [95:0] muls_2; // @[core.scala 230:17]
  reg [95:0] muls_3; // @[core.scala 230:17]
  reg [95:0] muls_4; // @[core.scala 230:17]
  reg [95:0] muls_5; // @[core.scala 230:17]
  reg [63:0] extnMResponse_result; // @[core.scala 235:30]
  reg [3:0] extnMResponse_robAddr; // @[core.scala 235:30]
  reg  division_request_valid; // @[core.scala 237:25]
  reg [63:0] division_request_rs1; // @[core.scala 237:25]
  reg [63:0] division_request_rs2; // @[core.scala 237:25]
  reg [31:0] division_request_instruction; // @[core.scala 237:25]
  reg [5:0] division_request_prfDest; // @[core.scala 237:25]
  reg [3:0] division_request_robAddr; // @[core.scala 237:25]
  reg [4:0] division_request_branchMask; // @[core.scala 237:25]
  reg [64:0] division_quotient; // @[core.scala 237:25]
  reg [64:0] division_remainder; // @[core.scala 237:25]
  reg [64:0] division_divisor; // @[core.scala 237:25]
  reg [6:0] division_counter; // @[core.scala 237:25]
  reg  fwdBuffers_0_valid; // @[core.scala 246:27]
  reg [5:0] fwdBuffers_0_prfDest; // @[core.scala 246:27]
  reg [63:0] fwdBuffers_0_result; // @[core.scala 246:27]
  reg  fwdBuffers_1_valid; // @[core.scala 246:27]
  reg [5:0] fwdBuffers_1_prfDest; // @[core.scala 246:27]
  reg [63:0] fwdBuffers_1_result; // @[core.scala 246:27]
  wire  _fwdFrom_0_valid_T_1 = |singleCycleArithmeticRequest_instruction[11:7]; // @[core.scala 255:109]
  wire  fwdFrom_0_valid = singleCycleArithmeticRequest_valid & |singleCycleArithmeticRequest_instruction[11:7]; // @[core.scala 255:58]
  wire  _addressGenerationInput_rs1_T_1 = |prf_toExec_instruction[19:15]; // @[core.scala 259:68]
  wire  _addressGenerationInput_rs1_T_3 = fwdFrom_0_valid & singleCycleArithmeticRequest_prfDest == prf_toExec_rs1Addr; // @[core.scala 260:34]
  wire  _addressGenerationInput_rs1_T_5 = fwdBuffers_0_valid & fwdBuffers_0_prfDest == prf_toExec_rs1Addr; // @[core.scala 260:34]
  wire  _addressGenerationInput_rs1_T_7 = fwdBuffers_1_valid & fwdBuffers_1_prfDest == prf_toExec_rs1Addr; // @[core.scala 260:34]
  wire [1:0] _arithmeticResult_arithmetic32_T_56 = {singleCycleArithmeticRequest_instruction[14],
    singleCycleArithmeticRequest_instruction[12]}; // @[Cat.scala 33:92]
  wire [31:0] _arithmeticResult_arithmetic32_T_36 = singleCycleArithmeticRequest_rs1[31:0]; // @[core.scala 275:69]
  wire [31:0] _arithmeticResult_arithmetic32_T_39 = $signed(_arithmeticResult_arithmetic32_T_36) >>>
    singleCycleArithmeticRequest_rs2[4:0]; // @[core.scala 275:90]
  wire [31:0] _arithmeticResult_arithmetic32_T_42 = _arithmeticResult_arithmetic32_T_39[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _arithmeticResult_arithmetic32_T_44 = {_arithmeticResult_arithmetic32_T_42,
    _arithmeticResult_arithmetic32_T_39}; // @[Cat.scala 33:92]
  wire [31:0] _arithmeticResult_arithmetic32_T_47 = singleCycleArithmeticRequest_rs1[31:0] >>
    singleCycleArithmeticRequest_rs2[4:0]; // @[core.scala 275:122]
  wire [31:0] _arithmeticResult_arithmetic32_T_50 = _arithmeticResult_arithmetic32_T_47[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _arithmeticResult_arithmetic32_T_52 = {_arithmeticResult_arithmetic32_T_50,
    _arithmeticResult_arithmetic32_T_47}; // @[Cat.scala 33:92]
  wire [63:0] _arithmeticResult_arithmetic32_T_53 = singleCycleArithmeticRequest_instruction[30] ?
    _arithmeticResult_arithmetic32_T_44 : _arithmeticResult_arithmetic32_T_52; // @[core.scala 275:20]
  wire [94:0] _GEN_250 = {{31'd0}, singleCycleArithmeticRequest_rs1}; // @[core.scala 274:34]
  wire [94:0] _arithmeticResult_arithmetic32_T_27 = _GEN_250 << singleCycleArithmeticRequest_rs2[4:0]; // @[core.scala 274:34]
  wire [31:0] _arithmeticResult_arithmetic32_T_30 = _arithmeticResult_arithmetic32_T_27[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _arithmeticResult_arithmetic32_T_32 = {_arithmeticResult_arithmetic32_T_30,
    _arithmeticResult_arithmetic32_T_27[31:0]}; // @[Cat.scala 33:92]
  wire [1:0] _arithmeticResult_arithmetic32_T_2 = {singleCycleArithmeticRequest_instruction[30],
    singleCycleArithmeticRequest_instruction[5]}; // @[Cat.scala 33:92]
  wire  _arithmeticResult_arithmetic32_T_3 = _arithmeticResult_arithmetic32_T_2 == 2'h3; // @[core.scala 272:58]
  wire [63:0] _arithmeticResult_arithmetic32_T_5 = singleCycleArithmeticRequest_rs1 - singleCycleArithmeticRequest_rs2; // @[core.scala 272:87]
  wire [31:0] _arithmeticResult_arithmetic32_T_8 = _arithmeticResult_arithmetic32_T_5[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _arithmeticResult_arithmetic32_T_10 = {_arithmeticResult_arithmetic32_T_8,
    _arithmeticResult_arithmetic32_T_5[31:0]}; // @[Cat.scala 33:92]
  wire [63:0] _arithmeticResult_arithmetic32_T_12 = singleCycleArithmeticRequest_rs1 + singleCycleArithmeticRequest_rs2; // @[core.scala 272:111]
  wire [31:0] _arithmeticResult_arithmetic32_T_15 = _arithmeticResult_arithmetic32_T_12[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _arithmeticResult_arithmetic32_T_17 = {_arithmeticResult_arithmetic32_T_15,
    _arithmeticResult_arithmetic32_T_12[31:0]}; // @[Cat.scala 33:92]
  wire [63:0] _arithmeticResult_arithmetic32_T_18 = _arithmeticResult_arithmetic32_T_2 == 2'h3 ?
    _arithmeticResult_arithmetic32_T_10 : _arithmeticResult_arithmetic32_T_17; // @[core.scala 272:20]
  wire [63:0] _GEN_36 = 2'h1 == _arithmeticResult_arithmetic32_T_56 ? _arithmeticResult_arithmetic32_T_32 :
    _arithmeticResult_arithmetic32_T_18; // @[core.scala 291:{8,8}]
  wire [63:0] _GEN_37 = 2'h2 == _arithmeticResult_arithmetic32_T_56 ? _arithmeticResult_arithmetic32_T_32 : _GEN_36; // @[core.scala 291:{8,8}]
  wire [63:0] _GEN_38 = 2'h3 == _arithmeticResult_arithmetic32_T_56 ? _arithmeticResult_arithmetic32_T_53 : _GEN_37; // @[core.scala 291:{8,8}]
  wire [63:0] _arithmeticResult_arithmetic64_T_26 = singleCycleArithmeticRequest_rs1 & singleCycleArithmeticRequest_rs2; // @[core.scala 289:22]
  wire [126:0] _arithmeticResult_arithmetic64_WIRE_7 = {{63'd0}, _arithmeticResult_arithmetic64_T_26}; // @[core.scala 281:{43,43}]
  wire [63:0] _arithmeticResult_arithmetic64_T_25 = singleCycleArithmeticRequest_rs1 | singleCycleArithmeticRequest_rs2; // @[core.scala 288:22]
  wire [126:0] _arithmeticResult_arithmetic64_WIRE_6 = {{63'd0}, _arithmeticResult_arithmetic64_T_25}; // @[core.scala 281:{43,43}]
  wire [63:0] _arithmeticResult_arithmetic64_T_21 = $signed(singleCycleArithmeticRequest_rs1) >>>
    singleCycleArithmeticRequest_rs2[5:0]; // @[core.scala 287:71]
  wire [63:0] _arithmeticResult_arithmetic64_T_23 = singleCycleArithmeticRequest_rs1 >> singleCycleArithmeticRequest_rs2
    [5:0]; // @[core.scala 287:84]
  wire [63:0] _arithmeticResult_arithmetic64_T_24 = singleCycleArithmeticRequest_instruction[30] ?
    _arithmeticResult_arithmetic64_T_21 : _arithmeticResult_arithmetic64_T_23; // @[core.scala 287:20]
  wire [126:0] _arithmeticResult_arithmetic64_WIRE_5 = {{63'd0}, _arithmeticResult_arithmetic64_T_24}; // @[core.scala 281:{43,43}]
  wire [63:0] _arithmeticResult_arithmetic64_T_15 = singleCycleArithmeticRequest_rs1 ^ singleCycleArithmeticRequest_rs2; // @[core.scala 286:22]
  wire [126:0] _arithmeticResult_arithmetic64_WIRE_4 = {{63'd0}, _arithmeticResult_arithmetic64_T_15}; // @[core.scala 281:{43,43}]
  wire  _arithmeticResult_arithmetic64_T_14 = singleCycleArithmeticRequest_rs1 < singleCycleArithmeticRequest_rs2; // @[core.scala 285:22]
  wire [126:0] _arithmeticResult_arithmetic64_WIRE_3 = {{126'd0}, _arithmeticResult_arithmetic64_T_14}; // @[core.scala 281:{43,43}]
  wire  _arithmeticResult_arithmetic64_T_13 = $signed(singleCycleArithmeticRequest_rs1) < $signed(
    singleCycleArithmeticRequest_rs2); // @[core.scala 284:29]
  wire [126:0] _arithmeticResult_arithmetic64_WIRE_2 = {{126'd0}, _arithmeticResult_arithmetic64_T_13}; // @[core.scala 281:{43,43}]
  wire [126:0] _GEN_252 = {{63'd0}, singleCycleArithmeticRequest_rs1}; // @[core.scala 283:22]
  wire [126:0] _arithmeticResult_arithmetic64_T_10 = _GEN_252 << singleCycleArithmeticRequest_rs2[5:0]; // @[core.scala 283:22]
  wire [63:0] _arithmeticResult_arithmetic64_T_8 = _arithmeticResult_arithmetic32_T_3 ?
    _arithmeticResult_arithmetic32_T_5 : _arithmeticResult_arithmetic32_T_12; // @[core.scala 282:20]
  wire [126:0] _arithmeticResult_arithmetic64_WIRE_0 = {{63'd0}, _arithmeticResult_arithmetic64_T_8}; // @[core.scala 281:{43,43}]
  wire [126:0] _GEN_40 = 3'h1 == singleCycleArithmeticRequest_instruction[14:12] ? _arithmeticResult_arithmetic64_T_10
     : _arithmeticResult_arithmetic64_WIRE_0; // @[core.scala 291:{8,8}]
  wire [126:0] _GEN_41 = 3'h2 == singleCycleArithmeticRequest_instruction[14:12] ? _arithmeticResult_arithmetic64_WIRE_2
     : _GEN_40; // @[core.scala 291:{8,8}]
  wire [126:0] _GEN_42 = 3'h3 == singleCycleArithmeticRequest_instruction[14:12] ? _arithmeticResult_arithmetic64_WIRE_3
     : _GEN_41; // @[core.scala 291:{8,8}]
  wire [126:0] _GEN_43 = 3'h4 == singleCycleArithmeticRequest_instruction[14:12] ? _arithmeticResult_arithmetic64_WIRE_4
     : _GEN_42; // @[core.scala 291:{8,8}]
  wire [126:0] _GEN_44 = 3'h5 == singleCycleArithmeticRequest_instruction[14:12] ? _arithmeticResult_arithmetic64_WIRE_5
     : _GEN_43; // @[core.scala 291:{8,8}]
  wire [126:0] _GEN_45 = 3'h6 == singleCycleArithmeticRequest_instruction[14:12] ? _arithmeticResult_arithmetic64_WIRE_6
     : _GEN_44; // @[core.scala 291:{8,8}]
  wire [126:0] _GEN_46 = 3'h7 == singleCycleArithmeticRequest_instruction[14:12] ? _arithmeticResult_arithmetic64_WIRE_7
     : _GEN_45; // @[core.scala 291:{8,8}]
  wire [126:0] arithmeticResult = singleCycleArithmeticRequest_instruction[3] ? {{63'd0}, _GEN_38} : _GEN_46; // @[core.scala 291:8]
  wire [63:0] fwdFrom_0_result = arithmeticResult[63:0]; // @[core.scala 252:33 293:21]
  wire [51:0] _arithmeticImm_T_2 = prf_toExec_instruction[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 77:12]
  wire [63:0] arithmeticImm = {_arithmeticImm_T_2,prf_toExec_instruction[31:20]}; // @[Cat.scala 33:92]
  wire [2:0] _singleCycleArithmeticRequest_valid_T_1 = prf_toExec_instruction[4:2] & 3'h5; // @[core.scala 298:91]
  wire  _singleCycleArithmeticRequest_rs2_T_5 = fwdFrom_0_valid & singleCycleArithmeticRequest_prfDest ==
    prf_toExec_rs2Addr; // @[core.scala 307:34]
  wire  _singleCycleArithmeticRequest_rs2_T_7 = fwdBuffers_0_valid & fwdBuffers_0_prfDest == prf_toExec_rs2Addr; // @[core.scala 307:34]
  wire  _singleCycleArithmeticRequest_rs2_T_9 = fwdBuffers_1_valid & fwdBuffers_1_prfDest == prf_toExec_rs2Addr; // @[core.scala 307:34]
  wire [63:0] _singleCycleArithmeticRequest_rs2_T_10 = _singleCycleArithmeticRequest_rs2_T_9 ? fwdBuffers_1_result :
    prf_toExec_rs2Data; // @[Mux.scala 101:16]
  wire [4:0] _T_30 = branchEvals_branchMask & singleCycleArithmeticRequest_branchMask; // @[core.scala 326:53]
  wire [4:0] _extnMRequest_valid_T_1 = prf_toExec_instruction[6:2] & 5'h1d; // @[core.scala 332:75]
  wire  _GEN_54 = _T_14 ? 1'h0 : prf_toExec_valid & 5'hc == _extnMRequest_valid_T_1 & prf_toExec_instruction[25]; // @[core.scala 332:22 339:83 340:26]
  wire  _GEN_56 = branchEvals_valid ? _GEN_54 : prf_toExec_valid & 5'hc == _extnMRequest_valid_T_1 &
    prf_toExec_instruction[25]; // @[core.scala 332:22 335:25]
  wire [32:0] _partialMuls32x32_T_7 = {extnMRequest_rs1[63],extnMRequest_rs1[63:32]}; // @[core.scala 355:57]
  wire [32:0] _partialMuls32x32_T_10 = {1'h0,extnMRequest_rs2[31:0]}; // @[core.scala 355:105]
  wire [32:0] _partialMuls32x32_T_15 = {1'h0,extnMRequest_rs1[31:0]}; // @[core.scala 357:44]
  wire [32:0] _partialMuls32x32_T_19 = {extnMRequest_rs2[63],extnMRequest_rs2[63:32]}; // @[core.scala 357:105]
  wire [32:0] _partialMuls32x32_T_28 = {1'h0,extnMRequest_rs2[63:32]}; // @[core.scala 359:106]
  wire [31:0] _partialMuls32x32_T_30 = extnMRequest_rs1[63:32]; // @[core.scala 360:30]
  wire [31:0] _partialMuls32x32_T_32 = extnMRequest_rs2[63:32]; // @[core.scala 360:64]
  wire [31:0] _partialMuls32x32_T_34 = extnMRequest_rs1[31:0]; // @[core.scala 361:29]
  wire [31:0] _partialMuls32x32_T_36 = extnMRequest_rs2[31:0]; // @[core.scala 361:62]
  reg [63:0] narrowMuls_0; // @[core.scala 363:23]
  reg [63:0] narrowMuls_1; // @[core.scala 363:23]
  reg [63:0] narrowMuls_2; // @[core.scala 363:23]
  reg [63:0] narrowMuls_3; // @[core.scala 363:23]
  reg [63:0] narrowMuls_4; // @[core.scala 363:23]
  reg [63:0] narrowMuls_5; // @[core.scala 363:23]
  reg [63:0] narrowMuls_6; // @[core.scala 363:23]
  reg [63:0] narrowMuls_7; // @[core.scala 363:23]
  reg [63:0] narrowMuls_8; // @[core.scala 363:23]
  wire [65:0] _T_39 = $signed(_partialMuls32x32_T_7) * $signed(_partialMuls32x32_T_10); // @[core.scala 364:41]
  wire [65:0] _T_40 = $signed(_partialMuls32x32_T_15) * $signed(_partialMuls32x32_T_19); // @[core.scala 364:41]
  wire [65:0] _T_41 = $signed(_partialMuls32x32_T_7) * $signed(_partialMuls32x32_T_28); // @[core.scala 364:41]
  wire [95:0] _muls_0_T = {narrowMuls_1,32'h0}; // @[Cat.scala 33:92]
  wire [95:0] _GEN_94 = {{32'd0}, narrowMuls_0}; // @[core.scala 367:29]
  wire [95:0] _muls_1_T = {narrowMuls_5,32'h0}; // @[Cat.scala 33:92]
  wire [95:0] _GEN_108 = {{32'd0}, narrowMuls_3}; // @[core.scala 368:28]
  wire [95:0] _muls_2_T = {narrowMuls_6,32'h0}; // @[Cat.scala 33:92]
  wire [31:0] _muls_3_T_2 = narrowMuls_4[63] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [95:0] _muls_3_T_3 = {_muls_3_T_2,narrowMuls_4}; // @[Cat.scala 33:92]
  wire [95:0] _muls_3_T_4 = {narrowMuls_7,32'h0}; // @[Cat.scala 33:92]
  wire [95:0] _muls_4_T = {narrowMuls_2,32'h0}; // @[Cat.scala 33:92]
  wire [31:0] _extnMResponse_result_T_4 = muls_5[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _extnMResponse_result_T_6 = {_extnMResponse_result_T_4,muls_5[31:0]}; // @[Cat.scala 33:92]
  wire [31:0] _extnMResponse_result_T_9 = muls_4[95] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [127:0] _extnMResponse_result_T_10 = {_extnMResponse_result_T_9,muls_4}; // @[Cat.scala 33:92]
  wire [127:0] _extnMResponse_result_T_11 = {muls_3,32'h0}; // @[Cat.scala 33:92]
  wire [127:0] _extnMResponse_result_T_13 = _extnMResponse_result_T_10 + _extnMResponse_result_T_11; // @[core.scala 379:42]
  wire [127:0] _extnMResponse_result_T_27 = {muls_2,32'h0}; // @[Cat.scala 33:92]
  wire [127:0] _extnMResponse_result_T_29 = _extnMResponse_result_T_10 + _extnMResponse_result_T_27; // @[core.scala 381:42]
  wire [127:0] _extnMResponse_result_T_31 = {muls_1,32'h0}; // @[Cat.scala 33:92]
  wire [127:0] _GEN_144 = {{32'd0}, muls_0}; // @[core.scala 382:14]
  wire [127:0] _extnMResponse_result_T_33 = _GEN_144 + _extnMResponse_result_T_31; // @[core.scala 382:14]
  wire [63:0] _GEN_58 = 2'h1 == extnMServicing_instruction[13:12] ? _extnMResponse_result_T_13[127:64] :
    _extnMResponse_result_T_13[63:0]; // @[core.scala 377:{30,30}]
  wire [63:0] _GEN_59 = 2'h2 == extnMServicing_instruction[13:12] ? _extnMResponse_result_T_29[127:64] : _GEN_58; // @[core.scala 377:{30,30}]
  wire [63:0] _GEN_60 = 2'h3 == extnMServicing_instruction[13:12] ? _extnMResponse_result_T_33[127:64] : _GEN_59; // @[core.scala 377:{30,30}]
  wire [63:0] _extnMResponse_result_T_36 = extnMServicing_instruction[3] ? _extnMResponse_result_T_6 : _GEN_60; // @[core.scala 377:30]
  wire [63:0] _GEN_61 = extnMServicing_valid & (~(|extnMServicing_instruction[24:20]) | ~(|extnMServicing_instruction[19
    :15])) ? 64'h0 : _extnMResponse_result_T_36; // @[core.scala 384:118 377:24 385:26]
  wire [4:0] _T_55 = extnMRequest_branchMask ^ branchEvals_branchMask; // @[core.scala 392:103]
  wire [4:0] _T_56 = extnMRequest_branchMask & branchEvals_branchMask; // @[core.scala 392:130]
  wire  _T_57 = |_T_56; // @[core.scala 392:154]
  wire [4:0] _T_58 = extnMPartialServicing_branchMask ^ branchEvals_branchMask; // @[core.scala 392:103]
  wire [4:0] _T_59 = extnMPartialServicing_branchMask & branchEvals_branchMask; // @[core.scala 392:130]
  wire  _T_60 = |_T_59; // @[core.scala 392:154]
  wire [4:0] _T_64 = extnMServicing_branchMask & branchEvals_branchMask; // @[core.scala 398:93]
  wire  _T_67 = |_T_64; // @[core.scala 398:123]
  wire  _GEN_67 = _T_67 & extnMServicing_valid ? 1'h0 : extnMServicing_valid; // @[core.scala 400:{101,107} 388:23]
  reg [4:0] divBranchMask; // @[core.scala 404:26]
  wire [4:0] _T_74 = {scheduler_release_instruction[25],scheduler_release_instruction[14],scheduler_release_instruction[
    6:4]}; // @[Cat.scala 33:92]
  wire  _T_75 = _T_74 == 5'h1b; // @[core.scala 406:115]
  wire  _T_76 = scheduler_release_fired & _T_75; // @[core.scala 405:32]
  wire [4:0] _mExtensionReady_T = branchEvals_branchMask & scheduler_release_branchMask; // @[core.scala 408:77]
  wire  _mExtensionReady_T_2 = branchEvals_valid & |_mExtensionReady_T; // @[core.scala 408:52]
  wire [4:0] _divBranchMask_T_3 = scheduler_release_branchMask ^ branchEvals_branchMask; // @[core.scala 410:133]
  wire [4:0] _divBranchMask_T_4 = _mExtensionReady_T_2 ? _divBranchMask_T_3 : scheduler_release_branchMask; // @[core.scala 410:25]
  wire  _GEN_77 = _T_76 ? branchEvals_valid & |_mExtensionReady_T & _T : mExtensionReady; // @[core.scala 406:132 408:21 141:32]
  wire [4:0] _GEN_78 = _T_76 ? _divBranchMask_T_4 : divBranchMask; // @[core.scala 406:132 410:19 404:26]
  wire [4:0] _T_78 = branchEvals_branchMask & divBranchMask; // @[core.scala 413:51]
  wire [4:0] _divBranchMask_T_5 = divBranchMask ^ branchEvals_branchMask; // @[core.scala 415:40]
  wire  _GEN_80 = _T | _GEN_77; // @[core.scala 417:31 418:25]
  wire  _GEN_82 = branchEvals_valid & |_T_78 ? _GEN_80 : _GEN_77; // @[core.scala 413:73]
  wire  _GEN_84 = ~mExtensionReady ? _GEN_82 : _GEN_77; // @[core.scala 412:26]
  wire  _GEN_85 = extnMResponse_valid & extnResponseInstruction[14] | _GEN_84; // @[core.scala 422:{67,85}]
  wire [64:0] _division_remainder_T_2 = {division_remainder[63:0],division_quotient[64]}; // @[Cat.scala 33:92]
  wire [64:0] _division_remainder_T_6 = 65'h0 - division_divisor; // @[core.scala 424:134]
  wire [64:0] _division_remainder_T_7 = division_remainder[64] ? division_divisor : _division_remainder_T_6; // @[core.scala 424:84]
  wire [64:0] _division_remainder_T_9 = _division_remainder_T_2 + _division_remainder_T_7; // @[core.scala 424:79]
  wire  _division_quotient_T_12 = ~_division_remainder_T_9[64]; // @[core.scala 425:54]
  wire [64:0] _division_quotient_T_13 = {division_quotient[63:0],_division_quotient_T_12}; // @[Cat.scala 33:92]
  wire [6:0] _division_counter_T_1 = division_counter - 7'h1; // @[core.scala 426:40]
  wire [64:0] _division_divisor_T_1 = {33'h0,extnMRequest_rs2[31:0]}; // @[Cat.scala 33:92]
  wire [64:0] _division_quotient_T_15 = {33'h0,extnMRequest_rs1[31:0]}; // @[Cat.scala 33:92]
  wire [64:0] _GEN_86 = extnMRequest_instruction[3] ? _division_divisor_T_1 : {{1'd0}, extnMRequest_rs2}; // @[core.scala 430:22 432:46 433:24]
  wire [64:0] _GEN_87 = extnMRequest_instruction[3] ? _division_quotient_T_15 : {{1'd0}, extnMRequest_rs1}; // @[core.scala 431:23 432:46 434:25]
  wire [63:0] _division_quotient_T_17 = 64'h0 - extnMRequest_rs1; // @[core.scala 441:79]
  wire [64:0] _division_quotient_T_19 = {1'h0,_division_quotient_T_17}; // @[Cat.scala 33:92]
  wire [64:0] _GEN_88 = extnMRequest_rs1[63] ? _division_quotient_T_19 : _GEN_87; // @[core.scala 441:{41,61}]
  wire [63:0] _division_divisor_T_3 = 64'h0 - extnMRequest_rs2; // @[core.scala 442:78]
  wire [64:0] _division_divisor_T_5 = {1'h0,_division_divisor_T_3}; // @[Cat.scala 33:92]
  wire [64:0] _GEN_89 = extnMRequest_rs2[63] ? _division_divisor_T_5 : _GEN_86; // @[core.scala 442:{41,60}]
  wire [31:0] _division_quotient_T_22 = 32'h0 - extnMRequest_rs1[31:0]; // @[core.scala 444:82]
  wire [64:0] _division_quotient_T_24 = {33'h0,_division_quotient_T_22}; // @[Cat.scala 33:92]
  wire [31:0] _division_divisor_T_8 = 32'h0 - extnMRequest_rs2[31:0]; // @[core.scala 445:81]
  wire [64:0] _division_divisor_T_10 = {33'h0,_division_divisor_T_8}; // @[Cat.scala 33:92]
  wire  _GEN_101 = extnMRequest_valid & extnMRequest_instruction[14] ? extnMRequest_valid : division_request_valid; // @[core.scala 428:67 437:22 237:25]
  wire [4:0] _GEN_107 = extnMRequest_valid & extnMRequest_instruction[14] ? extnMRequest_branchMask :
    division_request_branchMask; // @[core.scala 428:67 437:22 237:25]
  wire  _extnMResponse_result_quotient32_T_6 = ~(division_quotient == 65'h1ffffffffffffffff); // @[core.scala 453:99]
  wire [64:0] _extnMResponse_result_quotient32_T_9 = 65'h0 - division_quotient; // @[core.scala 453:125]
  wire [31:0] extnMResponse_result_quotient32 = (division_request_rs1[31] ^ division_request_rs2[31]) & ~(
    division_quotient == 65'h1ffffffffffffffff) ? _extnMResponse_result_quotient32_T_9[31:0] : division_quotient[31:0]; // @[core.scala 453:27]
  wire [64:0] _extnMResponse_result_remainder64Unsigned_T_3 = division_remainder + division_divisor; // @[core.scala 454:87]
  wire [64:0] extnMResponse_result_remainder64Unsigned = division_remainder[64] ?
    _extnMResponse_result_remainder64Unsigned_T_3 : division_remainder; // @[core.scala 454:36]
  wire [64:0] _extnMResponse_result_remainder32Signed_T_3 = 65'h0 - extnMResponse_result_remainder64Unsigned; // @[core.scala 455:70]
  wire [64:0] extnMResponse_result_remainder32Signed = division_request_rs1[31] ?
    _extnMResponse_result_remainder32Signed_T_3 : extnMResponse_result_remainder64Unsigned; // @[core.scala 455:34]
  wire [64:0] _extnMResponse_result_T_47 = (division_request_rs1[63] ^ division_request_rs2[63]) &
    _extnMResponse_result_quotient32_T_6 ? _extnMResponse_result_quotient32_T_9 : division_quotient; // @[core.scala 458:10]
  wire [64:0] _extnMResponse_result_T_52 = division_request_rs1[63] ? _extnMResponse_result_remainder32Signed_T_3 :
    extnMResponse_result_remainder64Unsigned; // @[core.scala 460:10]
  wire [31:0] _extnMResponse_result_T_55 = extnMResponse_result_quotient32[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _extnMResponse_result_T_57 = {_extnMResponse_result_T_55,extnMResponse_result_quotient32}; // @[Cat.scala 33:92]
  wire [31:0] _extnMResponse_result_T_60 = division_quotient[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _extnMResponse_result_T_62 = {_extnMResponse_result_T_60,division_quotient[31:0]}; // @[Cat.scala 33:92]
  wire [31:0] _extnMResponse_result_T_65 = extnMResponse_result_remainder32Signed[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _extnMResponse_result_T_67 = {_extnMResponse_result_T_65,extnMResponse_result_remainder32Signed[31:0]}; // @[Cat.scala 33:92]
  wire [31:0] _extnMResponse_result_T_70 = extnMResponse_result_remainder64Unsigned[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _extnMResponse_result_T_72 = {_extnMResponse_result_T_70,extnMResponse_result_remainder64Unsigned[31:0]}; // @[Cat.scala 33:92]
  wire [2:0] _extnMResponse_result_T_75 = {division_request_instruction[3],division_request_instruction[13:12]}; // @[Cat.scala 33:92]
  wire [64:0] _GEN_110 = 3'h1 == _extnMResponse_result_T_75 ? division_quotient : _extnMResponse_result_T_47; // @[core.scala 452:{26,26}]
  wire [64:0] _GEN_111 = 3'h2 == _extnMResponse_result_T_75 ? _extnMResponse_result_T_52 : _GEN_110; // @[core.scala 452:{26,26}]
  wire [64:0] _GEN_112 = 3'h3 == _extnMResponse_result_T_75 ? extnMResponse_result_remainder64Unsigned : _GEN_111; // @[core.scala 452:{26,26}]
  wire [64:0] _extnMResponse_result_WIRE_1_4 = {{1'd0}, _extnMResponse_result_T_57}; // @[core.scala 457:{14,14}]
  wire [64:0] _GEN_113 = 3'h4 == _extnMResponse_result_T_75 ? _extnMResponse_result_WIRE_1_4 : _GEN_112; // @[core.scala 452:{26,26}]
  wire [64:0] _extnMResponse_result_WIRE_1_5 = {{1'd0}, _extnMResponse_result_T_62}; // @[core.scala 457:{14,14}]
  wire [64:0] _GEN_114 = 3'h5 == _extnMResponse_result_T_75 ? _extnMResponse_result_WIRE_1_5 : _GEN_113; // @[core.scala 452:{26,26}]
  wire [64:0] _extnMResponse_result_WIRE_1_6 = {{1'd0}, _extnMResponse_result_T_67}; // @[core.scala 457:{14,14}]
  wire [64:0] _GEN_115 = 3'h6 == _extnMResponse_result_T_75 ? _extnMResponse_result_WIRE_1_6 : _GEN_114; // @[core.scala 452:{26,26}]
  wire [64:0] _extnMResponse_result_WIRE_1_7 = {{1'd0}, _extnMResponse_result_T_72}; // @[core.scala 457:{14,14}]
  wire [64:0] _GEN_116 = 3'h7 == _extnMResponse_result_T_75 ? _extnMResponse_result_WIRE_1_7 : _GEN_115; // @[core.scala 452:{26,26}]
  wire [4:0] _T_106 = division_request_branchMask & branchEvals_branchMask; // @[core.scala 475:41]
  wire  _T_107 = |_T_106; // @[core.scala 475:65]
  wire [64:0] _GEN_120 = division_request_valid & ~(|division_counter) ? _GEN_116 : {{1'd0}, _GEN_61}; // @[core.scala 450:57 452:26]
  wire  _GEN_124 = division_request_valid & ~(|division_counter) ? 1'h0 : _GEN_101; // @[core.scala 450:57 473:28]
  wire  _GEN_126 = _T & _T_57 ? 1'h0 : _GEN_124; // @[core.scala 482:{112,87}]
  wire [4:0] _division_request_branchMask_T_1 = division_request_branchMask ^ branchEvals_branchMask; // @[core.scala 484:130]
  reg  branchPCs_0_valid; // @[core.scala 500:26]
  reg [63:0] branchPCs_0_pc; // @[core.scala 500:26]
  reg [4:0] branchPCs_0_branchMask; // @[core.scala 500:26]
  reg  branchPCs_1_valid; // @[core.scala 500:26]
  reg [63:0] branchPCs_1_pc; // @[core.scala 500:26]
  reg [4:0] branchPCs_1_branchMask; // @[core.scala 500:26]
  reg  branchPCs_2_valid; // @[core.scala 500:26]
  reg [63:0] branchPCs_2_pc; // @[core.scala 500:26]
  reg [4:0] branchPCs_2_branchMask; // @[core.scala 500:26]
  reg  branchPCs_3_valid; // @[core.scala 500:26]
  reg [63:0] branchPCs_3_pc; // @[core.scala 500:26]
  reg [4:0] branchPCs_3_branchMask; // @[core.scala 500:26]
  reg  predictedPCs_0_valid; // @[core.scala 507:29]
  reg [63:0] predictedPCs_0_pc; // @[core.scala 507:29]
  reg  predictedPCs_1_valid; // @[core.scala 507:29]
  reg [63:0] predictedPCs_1_pc; // @[core.scala 507:29]
  reg  predictedPCs_2_valid; // @[core.scala 507:29]
  reg [63:0] predictedPCs_2_pc; // @[core.scala 507:29]
  reg  predictedPCs_3_valid; // @[core.scala 507:29]
  reg [63:0] predictedPCs_3_pc; // @[core.scala 507:29]
  reg  branchInstruction_valid; // @[core.scala 512:34]
  reg [63:0] branchInstruction_rs1; // @[core.scala 512:34]
  reg [63:0] branchInstruction_rs2; // @[core.scala 512:34]
  reg [3:0] branchInstruction_robAddr; // @[core.scala 512:34]
  reg [31:0] branchInstruction_instruction; // @[core.scala 512:34]
  reg [63:0] branchInstruction_immediate; // @[core.scala 512:34]
  wire [63:0] _branchInstruction_immediate_T_6 = {_arithmeticImm_T_2,prf_toExec_instruction[7],prf_toExec_instruction[30
    :25],prf_toExec_instruction[11:8],1'h0}; // @[Cat.scala 33:92]
  wire [43:0] _branchInstruction_immediate_T_14 = prf_toExec_instruction[31] ? 44'hfffffffffff : 44'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _branchInstruction_immediate_T_18 = {_branchInstruction_immediate_T_14,prf_toExec_instruction[19:12],
    prf_toExec_instruction[20],prf_toExec_instruction[30:21],1'h0}; // @[Cat.scala 33:92]
  reg [3:0] branchEvals_robAddr; // @[core.scala 534:28]
  reg [63:0] branchEvals_nextPC; // @[core.scala 534:28]
  wire [5:0] _GEN_140 = prf_toExec_valid & prf_toExec_instruction[6:5] == 2'h3 ? prf_toExec_robAddr : {{2'd0},
    branchInstruction_robAddr}; // @[core.scala 546:71 554:31 512:34]
  wire [4:0] _T_128 = branchEvals_branchMask & prf_toExec_branchmask; // @[core.scala 562:53]
  wire  _coherentLoadInvalid_T_5 = ~(|rob_commit_instruction[6:2]); // @[core.scala 568:141]
  wire  coherentLoadInvalid = ~memAccess_loadCommit_state & memAccess_loadCommit_valid & rob_commit_ready & ~(|
    rob_commit_instruction[6:2]); // @[core.scala 568:107]
  wire [3:0] _branchEvals_robAddr_T_1 = rob_commit_robAddr - 4'h1; // @[core.scala 572:68]
  wire [63:0] branchTaken_rs1 = |branchInstruction_instruction[19:15] ? branchInstruction_rs1 : 64'h0; // @[core.scala 583:18]
  wire [63:0] branchTaken_rs2 = |branchInstruction_instruction[24:20] ? branchInstruction_rs2 : 64'h0; // @[core.scala 584:18]
  wire  branchTaken_conditionEval_0 = branchTaken_rs1 == branchTaken_rs2; // @[core.scala 588:41]
  wire [63:0] _branchTaken_conditionEval_T_2 = |branchInstruction_instruction[19:15] ? branchInstruction_rs1 : 64'h0; // @[core.scala 588:67]
  wire [63:0] _branchTaken_conditionEval_T_3 = |branchInstruction_instruction[24:20] ? branchInstruction_rs2 : 64'h0; // @[core.scala 588:80]
  wire  branchTaken_conditionEval_4 = $signed(_branchTaken_conditionEval_T_2) < $signed(_branchTaken_conditionEval_T_3); // @[core.scala 588:74]
  wire  branchTaken_conditionEval_6 = branchTaken_rs1 < branchTaken_rs2; // @[core.scala 588:92]
  wire  branchTaken_conditionEval_1 = ~branchTaken_conditionEval_0; // @[core.scala 588:125]
  wire  branchTaken_conditionEval_5 = ~branchTaken_conditionEval_4; // @[core.scala 588:125]
  wire  branchTaken_conditionEval_7 = ~branchTaken_conditionEval_6; // @[core.scala 588:125]
  wire  nextCorrectPC_conditionEval_0 = branchInstruction_rs1 == branchInstruction_rs2; // @[core.scala 608:11]
  wire  nextCorrectPC_conditionEval_1 = branchInstruction_rs1 != branchInstruction_rs2; // @[core.scala 609:11]
  wire  nextCorrectPC_conditionEval_4 = $signed(branchInstruction_rs1) < $signed(branchInstruction_rs2); // @[core.scala 612:18]
  wire  nextCorrectPC_conditionEval_5 = $signed(branchInstruction_rs1) >= $signed(branchInstruction_rs2); // @[core.scala 613:18]
  wire  nextCorrectPC_conditionEval_6 = branchInstruction_rs1 < branchInstruction_rs2; // @[core.scala 614:11]
  wire  nextCorrectPC_conditionEval_7 = branchInstruction_rs1 >= branchInstruction_rs2; // @[core.scala 615:11]
  wire [63:0] _nextCorrectPC_T_2 = branchPCs_0_pc + branchInstruction_immediate; // @[core.scala 619:50]
  wire [63:0] _nextCorrectPC_T_4 = branchPCs_0_pc + 64'h4; // @[core.scala 619:66]
  wire  _GEN_149 = 3'h1 == branchInstruction_instruction[14:12] ? nextCorrectPC_conditionEval_1 :
    nextCorrectPC_conditionEval_0; // @[core.scala 619:{10,10}]
  wire  _GEN_150 = 3'h2 == branchInstruction_instruction[14:12] ? 1'h0 : _GEN_149; // @[core.scala 619:{10,10}]
  wire  _GEN_151 = 3'h3 == branchInstruction_instruction[14:12] ? 1'h0 : _GEN_150; // @[core.scala 619:{10,10}]
  wire  _GEN_152 = 3'h4 == branchInstruction_instruction[14:12] ? nextCorrectPC_conditionEval_4 : _GEN_151; // @[core.scala 619:{10,10}]
  wire  _GEN_153 = 3'h5 == branchInstruction_instruction[14:12] ? nextCorrectPC_conditionEval_5 : _GEN_152; // @[core.scala 619:{10,10}]
  wire  _GEN_154 = 3'h6 == branchInstruction_instruction[14:12] ? nextCorrectPC_conditionEval_6 : _GEN_153; // @[core.scala 619:{10,10}]
  wire  _GEN_155 = 3'h7 == branchInstruction_instruction[14:12] ? nextCorrectPC_conditionEval_7 : _GEN_154; // @[core.scala 619:{10,10}]
  wire [63:0] _nextCorrectPC_T_5 = _GEN_155 ? _nextCorrectPC_T_2 : _nextCorrectPC_T_4; // @[core.scala 619:10]
  wire [63:0] _nextCorrectPC_T_7 = branchInstruction_rs1 + branchInstruction_immediate; // @[core.scala 620:11]
  wire [63:0] _GEN_157 = 2'h1 == branchInstruction_instruction[3:2] ? _nextCorrectPC_T_7 : _nextCorrectPC_T_5; // @[core.scala 627:{28,28}]
  wire [63:0] _GEN_158 = 2'h2 == branchInstruction_instruction[3:2] ? 64'h0 : _GEN_157; // @[core.scala 627:{28,28}]
  wire [63:0] _GEN_159 = 2'h3 == branchInstruction_instruction[3:2] ? _nextCorrectPC_T_2 : _GEN_158; // @[core.scala 627:{28,28}]
  wire  _branchEvals_passed_T_2 = coherentLoadInvalid ? 1'h0 : predictedPCs_0_valid & _GEN_159 == predictedPCs_0_pc; // @[core.scala 629:28]
  wire  _T_133 = branchPCs_0_valid & branchPCs_1_valid; // @[core.scala 635:46]
  wire  _T_134 = branchPCs_0_valid & branchPCs_1_valid & branchPCs_2_valid; // @[core.scala 635:46]
  wire [63:0] _GEN_161 = ~branchPCs_0_valid ? decode_branchPCs_branchPC : branchPCs_0_pc; // @[core.scala 636:82 638:12 500:26]
  wire [4:0] _GEN_162 = ~branchPCs_0_valid ? decode_branchPCs_branchMask : branchPCs_0_branchMask; // @[core.scala 636:82 639:20 500:26]
  wire  _T_138 = ~branchPCs_1_valid; // @[core.scala 636:70]
  wire [63:0] _GEN_164 = branchPCs_0_valid & ~branchPCs_1_valid ? decode_branchPCs_branchPC : branchPCs_1_pc; // @[core.scala 636:82 638:12 500:26]
  wire [4:0] _GEN_165 = branchPCs_0_valid & ~branchPCs_1_valid ? decode_branchPCs_branchMask : branchPCs_1_branchMask; // @[core.scala 636:82 639:20 500:26]
  wire  _T_140 = ~branchPCs_2_valid; // @[core.scala 636:70]
  wire [63:0] _GEN_167 = _T_133 & ~branchPCs_2_valid ? decode_branchPCs_branchPC : branchPCs_2_pc; // @[core.scala 636:82 638:12 500:26]
  wire [4:0] _GEN_168 = _T_133 & ~branchPCs_2_valid ? decode_branchPCs_branchMask : branchPCs_2_branchMask; // @[core.scala 636:82 639:20 500:26]
  wire  _T_142 = ~branchPCs_3_valid; // @[core.scala 636:70]
  wire  _T_145 = branchEvals_valid & _T; // @[core.scala 641:24]
  wire  entry_1_valid = branchPCs_1_valid | decode_branchPCs_branchPCReady & (_T_138 & branchPCs_0_valid); // @[core.scala 647:32]
  wire  entry_2_valid = branchPCs_2_valid | decode_branchPCs_branchPCReady & (_T_140 & _T_133); // @[core.scala 647:32]
  wire  entry_3_valid = branchPCs_3_valid | decode_branchPCs_branchPCReady & (_T_142 & _T_134); // @[core.scala 647:32]
  wire  _T_151 = predictedPCs_0_valid & predictedPCs_1_valid; // @[core.scala 659:49]
  wire  _T_152 = predictedPCs_0_valid & predictedPCs_1_valid & predictedPCs_2_valid; // @[core.scala 659:49]
  wire [63:0] _GEN_193 = ~predictedPCs_0_valid ? decode_branchPCs_predictedPC : predictedPCs_0_pc; // @[core.scala 660:82 662:12 507:29]
  wire  _T_156 = ~predictedPCs_1_valid; // @[core.scala 660:70]
  wire [63:0] _GEN_195 = predictedPCs_0_valid & ~predictedPCs_1_valid ? decode_branchPCs_predictedPC : predictedPCs_1_pc
    ; // @[core.scala 660:82 662:12 507:29]
  wire  _T_158 = ~predictedPCs_2_valid; // @[core.scala 660:70]
  wire [63:0] _GEN_197 = _T_151 & ~predictedPCs_2_valid ? decode_branchPCs_predictedPC : predictedPCs_2_pc; // @[core.scala 660:82 662:12 507:29]
  wire  _T_160 = ~predictedPCs_3_valid; // @[core.scala 660:70]
  wire  entry_5_valid = predictedPCs_1_valid | decode_branchPCs_predictedPCReady & (_T_156 & predictedPCs_0_valid); // @[core.scala 670:32]
  wire  entry_6_valid = predictedPCs_2_valid | decode_branchPCs_predictedPCReady & (_T_158 & _T_151); // @[core.scala 670:32]
  wire  entry_7_valid = predictedPCs_3_valid | decode_branchPCs_predictedPCReady & (_T_160 & _T_152); // @[core.scala 670:32]
  reg  coherentLoadInvalidReg; // @[core.scala 708:39]
  wire  _GEN_215 = 3'h1 == branchInstruction_instruction[14:12] ? branchTaken_conditionEval_1 :
    branchTaken_conditionEval_0; // @[core.scala 712:{31,31}]
  wire  _GEN_216 = 3'h2 == branchInstruction_instruction[14:12] ? branchTaken_conditionEval_0 : _GEN_215; // @[core.scala 712:{31,31}]
  wire  _GEN_217 = 3'h3 == branchInstruction_instruction[14:12] ? branchTaken_conditionEval_1 : _GEN_216; // @[core.scala 712:{31,31}]
  wire  _GEN_218 = 3'h4 == branchInstruction_instruction[14:12] ? branchTaken_conditionEval_4 : _GEN_217; // @[core.scala 712:{31,31}]
  wire  _GEN_219 = 3'h5 == branchInstruction_instruction[14:12] ? branchTaken_conditionEval_5 : _GEN_218; // @[core.scala 712:{31,31}]
  wire  _GEN_220 = 3'h6 == branchInstruction_instruction[14:12] ? branchTaken_conditionEval_6 : _GEN_219; // @[core.scala 712:{31,31}]
  wire  _memAccess_writeInstructionCommit_fired_T_1 = rob_commit_instruction[6:4] == 3'h2; // @[core.scala 728:117]
  reg [63:0] rob_execPorts_0_mtval_REG; // @[core.scala 758:36]
  reg  REG; // @[core.scala 779:129]
  reg [5:0] prf_fromStore_rs2Addr_REG; // @[core.scala 815:43]
  reg [5:0] prf_fromStore_rs2Addr_REG_1; // @[core.scala 815:35]
  reg  prf_fromStore_valid_REG; // @[core.scala 816:41]
  reg  prf_fromStore_valid_REG_1; // @[core.scala 816:33]
  wire  _memAccess_initiateFence_T = rob_commit_fired & rob_commit_is_fence; // @[core.scala 858:47]
  reg [1:0] fenceState_state; // @[core.scala 862:27]
  reg [4:0] fenceState_branchMask; // @[core.scala 862:27]
  wire [19:0] _T_188 = fetch_toDecode_instruction[19:0] & 20'hfefff; // @[core.scala 871:72]
  wire [19:0] _T_195 = decode_toExec_instruction[19:0] & 20'hfefff; // @[core.scala 880:76]
  wire [1:0] _GEN_223 = decode_toExec_fired & _T_195 == 20'hf ? 2'h2 : fenceState_state; // @[core.scala 880:119 881:26 862:27]
  wire  _GEN_225 = _T_145 | rob_commit_fired & rob_commit_is_fence; // @[core.scala 858:27 876:54 878:33]
  wire [4:0] _T_199 = branchEvals_branchMask & fenceState_branchMask; // @[core.scala 886:57]
  wire  _T_201 = branchEvals_valid & |_T_199; // @[core.scala 886:30]
  wire [4:0] _fenceState_branchMask_T = fenceState_branchMask ^ branchEvals_branchMask; // @[core.scala 894:57]
  wire [4:0] _GEN_228 = _T_201 & branchEvals_passed ? _fenceState_branchMask_T : fenceState_branchMask; // @[core.scala 893:115 862:27 894:31]
  wire  _GEN_229 = rob_commit_fired & rob_commit_is_fence | rob_commit_fired & rob_commit_is_fence; // @[core.scala 858:27 890:59 891:33]
  wire [1:0] _GEN_230 = _memAccess_initiateFence_T ? 2'h0 : fenceState_state; // @[core.scala 890:59 892:26 862:27]
  wire [4:0] _GEN_231 = _memAccess_initiateFence_T ? fenceState_branchMask : _GEN_228; // @[core.scala 862:27 890:59]
  wire  _GEN_232 = branchEvals_valid & |_T_199 & _T | _GEN_229; // @[core.scala 886:110 888:33]
  wire [1:0] _GEN_233 = branchEvals_valid & |_T_199 & _T ? 2'h0 : _GEN_230; // @[core.scala 886:110 889:26]
  wire  _GEN_235 = 2'h2 == fenceState_state ? _GEN_232 : rob_commit_fired & rob_commit_is_fence; // @[core.scala 858:27 869:28]
  wire  _GEN_238 = 2'h1 == fenceState_state ? _GEN_225 : _GEN_235; // @[core.scala 869:28]
  wire  _GEN_242 = 2'h0 == fenceState_state ? rob_commit_fired & rob_commit_is_fence : _GEN_238; // @[core.scala 858:27 869:28]
  wire  _GEN_244 = _T_145 & fetch_cachelinesUpdatesResp_ready | _GEN_242; // @[core.scala 917:85 918:29]
  reg  REG_1; // @[core.scala 920:15]
  reg [2:0] branchCounter; // @[core.scala 1033:30]
  wire  _branchCounter_T_2 = decode_fromFetch_fired & decode_fromFetch_instruction[6:4] == 3'h6; // @[core.scala 1037:29]
  wire [2:0] _GEN_247 = {{2'd0}, _branchCounter_T_2}; // @[core.scala 1034:34]
  wire [3:0] _branchCounter_T_3 = branchCounter + _GEN_247; // @[core.scala 1034:34]
  wire [3:0] _GEN_248 = {{3'd0}, branchEvals_valid}; // @[core.scala 1037:81]
  wire [4:0] _branchCounter_T_4 = _branchCounter_T_3 - _GEN_248; // @[core.scala 1037:81]
  wire [4:0] _GEN_267 = _T_145 ? 5'h0 : _branchCounter_T_4; // @[core.scala 1034:17 1040:50 1043:19]
  reg [3:0] lastBranchExecRob; // @[core.scala 1047:30]
  reg [63:0] lastBranchExecPC; // @[core.scala 1048:29]
  reg [63:0] lastBranchExecPC_REG; // @[core.scala 1051:32]
  reg  lastRetiredSystem; // @[core.scala 1067:34]
  reg [1:0] interruptInjectStatus; // @[core.scala 1070:38]
  wire  _T_231 = |branchCounter; // @[core.scala 1081:60]
  wire [1:0] _GEN_272 = branchInstruction_valid & branchInstruction_instruction[6:0] == 7'h63 ? 2'h2 :
    interruptInjectStatus; // @[core.scala 1082:135 1070:38 1083:79]
  wire  _GEN_273 = branchInstruction_valid & branchInstruction_instruction[6:0] == 7'h63 ? 1'h0 :
    _branchEvals_passed_T_2; // @[core.scala 1082:135 1086:76 629:22]
  wire [1:0] _GEN_274 = decode_fromFetch_fired ? 2'h0 : interruptInjectStatus; // @[core.scala 1096:110 1070:38 1096:86]
  wire [63:0] _GEN_275 = fetch_toDecode_instruction[6:0] != 7'hf & fetch_toDecode_instruction[6:0] != 7'h73 ? 64'h80000073
     : {{32'd0}, fetch_toDecode_instruction}; // @[core.scala 1089:162 1091:86 70:32]
  wire [1:0] _GEN_276 = fetch_toDecode_instruction[6:0] != 7'hf & fetch_toDecode_instruction[6:0] != 7'h73 ? _GEN_274 :
    interruptInjectStatus; // @[core.scala 1089:162 1070:38]
  wire [1:0] _GEN_277 = |branchCounter ? _GEN_272 : _GEN_276; // @[core.scala 1081:65]
  wire  _GEN_278 = |branchCounter ? _GEN_273 : _branchEvals_passed_T_2; // @[core.scala 1081:65 629:22]
  wire [63:0] _GEN_279 = |branchCounter ? {{32'd0}, fetch_toDecode_instruction} : _GEN_275; // @[core.scala 1081:65 70:32]
  wire [1:0] _GEN_280 = ~branchEvals_valid ? _GEN_277 : interruptInjectStatus; // @[core.scala 1070:38 1080:58]
  wire [63:0] _GEN_282 = ~branchEvals_valid ? _GEN_279 : {{32'd0}, fetch_toDecode_instruction}; // @[core.scala 1080:58 70:32]
  wire [63:0] _GEN_285 = decode_canTakeInterrupt ? _GEN_282 : {{32'd0}, fetch_toDecode_instruction}; // @[core.scala 1079:56 70:32]
  wire [1:0] _GEN_286 = decode_writeBackResult_fired ? 2'h0 : interruptInjectStatus; // @[core.scala 1070:38 1110:{44,68}]
  wire [63:0] _GEN_287 = rob_commit_robAddr == lastBranchExecRob ? 64'h80000073 : {{32'd0}, rob_commit_instruction}; // @[core.scala 1106:54 1108:44 719:38]
  wire [1:0] _GEN_288 = rob_commit_robAddr == lastBranchExecRob ? _GEN_286 : interruptInjectStatus; // @[core.scala 1070:38 1106:54]
  wire [63:0] _GEN_289 = 2'h3 == interruptInjectStatus ? _GEN_287 : {{32'd0}, rob_commit_instruction}; // @[core.scala 1071:33 719:38]
  wire [1:0] _GEN_290 = 2'h3 == interruptInjectStatus ? _GEN_288 : interruptInjectStatus; // @[core.scala 1071:33 1070:38]
  wire [63:0] _GEN_292 = 2'h2 == interruptInjectStatus ? {{32'd0}, rob_commit_instruction} : _GEN_289; // @[core.scala 1071:33 719:38]
  wire [63:0] _GEN_295 = 2'h1 == interruptInjectStatus ? _GEN_285 : {{32'd0}, fetch_toDecode_instruction}; // @[core.scala 1071:33 70:32]
  wire [63:0] _GEN_296 = 2'h1 == interruptInjectStatus ? {{32'd0}, rob_commit_instruction} : _GEN_292; // @[core.scala 1071:33 719:38]
  wire [63:0] _GEN_299 = 2'h0 == interruptInjectStatus ? {{32'd0}, fetch_toDecode_instruction} : _GEN_295; // @[core.scala 1071:33 70:32]
  wire [63:0] _GEN_300 = 2'h0 == interruptInjectStatus ? {{32'd0}, rob_commit_instruction} : _GEN_296; // @[core.scala 1071:33 719:38]
  wire [4:0] _GEN_249 = reset ? 5'h0 : _GEN_267; // @[core.scala 1033:{30,30}]
  iCache icache ( // @[core.scala 28:22]
    .clock(icache_clock),
    .reset(icache_reset),
    .fromFetch_req_ready(icache_fromFetch_req_ready),
    .fromFetch_req_valid(icache_fromFetch_req_valid),
    .fromFetch_req_bits(icache_fromFetch_req_bits),
    .fromFetch_resp_ready(icache_fromFetch_resp_ready),
    .fromFetch_resp_valid(icache_fromFetch_resp_valid),
    .fromFetch_resp_bits(icache_fromFetch_resp_bits),
    .updateAllCachelines_ready(icache_updateAllCachelines_ready),
    .updateAllCachelines_fired(icache_updateAllCachelines_fired),
    .cachelinesUpdatesResp_ready(icache_cachelinesUpdatesResp_ready),
    .cachelinesUpdatesResp_fired(icache_cachelinesUpdatesResp_fired),
    .lowLevelMem_ARADDR(icache_lowLevelMem_ARADDR),
    .lowLevelMem_ARVALID(icache_lowLevelMem_ARVALID),
    .lowLevelMem_ARREADY(icache_lowLevelMem_ARREADY),
    .lowLevelMem_RDATA(icache_lowLevelMem_RDATA),
    .lowLevelMem_RLAST(icache_lowLevelMem_RLAST),
    .lowLevelMem_RVALID(icache_lowLevelMem_RVALID),
    .lowLevelMem_RREADY(icache_lowLevelMem_RREADY),
    .debug_probe_arvalid_internal(icache_debug_probe_arvalid_internal),
    .debug_probe_cacheMissed(icache_debug_probe_cacheMissed),
    .debug_probe_rready_signal(icache_debug_probe_rready_signal),
    .debug_probe_cacheFill_valid(icache_debug_probe_cacheFill_valid),
    .debug_probe_axi_arvalid(icache_debug_probe_axi_arvalid),
    .debug_probe_axi_arready(icache_debug_probe_axi_arready),
    .debug_probe_req_valid(icache_debug_probe_req_valid),
    .debug_probe_req_pc(icache_debug_probe_req_pc)
  );
  fetch fetch ( // @[core.scala 42:21]
    .clock(fetch_clock),
    .reset(fetch_reset),
    .cache_req_ready(fetch_cache_req_ready),
    .cache_req_valid(fetch_cache_req_valid),
    .cache_req_bits(fetch_cache_req_bits),
    .cache_resp_ready(fetch_cache_resp_ready),
    .cache_resp_valid(fetch_cache_resp_valid),
    .cache_resp_bits(fetch_cache_resp_bits),
    .toDecode_ready(fetch_toDecode_ready),
    .toDecode_fired(fetch_toDecode_fired),
    .toDecode_pc(fetch_toDecode_pc),
    .toDecode_instruction(fetch_toDecode_instruction),
    .toDecode_expected_valid(fetch_toDecode_expected_valid),
    .toDecode_expected_pc(fetch_toDecode_expected_pc),
    .toDecode_expected_coherency(fetch_toDecode_expected_coherency),
    .branchRes_fired(fetch_branchRes_fired),
    .branchRes_branchTaken(fetch_branchRes_branchTaken),
    .branchRes_pc(fetch_branchRes_pc),
    .branchRes_pcAfterBrnach(fetch_branchRes_pcAfterBrnach),
    .carryOutFence_ready(fetch_carryOutFence_ready),
    .carryOutFence_fired(fetch_carryOutFence_fired),
    .updateAllCachelines_ready(fetch_updateAllCachelines_ready),
    .updateAllCachelines_fired(fetch_updateAllCachelines_fired),
    .cachelinesUpdatesResp_ready(fetch_cachelinesUpdatesResp_ready),
    .cachelinesUpdatesResp_fired(fetch_cachelinesUpdatesResp_fired),
    .fdbg_probe_redirect_bit(fetch_fdbg_probe_redirect_bit),
    .fdbg_probe_fifo_enq_ready(fetch_fdbg_probe_fifo_enq_ready),
    .fdbg_probe_is_fence(fetch_fdbg_probe_is_fence),
    .fdbg_probe_handle_fence(fetch_fdbg_probe_handle_fence)
  );
  core_Anon decode ( // @[core.scala 57:22]
    .clock(decode_clock),
    .reset(decode_reset),
    .fromFetch_ready(decode_fromFetch_ready),
    .fromFetch_fired(decode_fromFetch_fired),
    .fromFetch_pc(decode_fromFetch_pc),
    .fromFetch_instruction(decode_fromFetch_instruction),
    .fromFetch_expected_valid(decode_fromFetch_expected_valid),
    .fromFetch_expected_pc(decode_fromFetch_expected_pc),
    .fromFetch_expected_coherency(decode_fromFetch_expected_coherency),
    .toExec_ready(decode_toExec_ready),
    .toExec_fired(decode_toExec_fired),
    .toExec_instruction(decode_toExec_instruction),
    .toExec_pc(decode_toExec_pc),
    .toExec_PRFDest(decode_toExec_PRFDest),
    .toExec_rs1Addr(decode_toExec_rs1Addr),
    .toExec_rs1Ready(decode_toExec_rs1Ready),
    .toExec_rs2Addr(decode_toExec_rs2Addr),
    .toExec_rs2Ready(decode_toExec_rs2Ready),
    .toExec_branchMask(decode_toExec_branchMask),
    .writeBackResult_fired(decode_writeBackResult_fired),
    .writeBackResult_instruction(decode_writeBackResult_instruction),
    .writeBackResult_rdAddr(decode_writeBackResult_rdAddr),
    .writeBackResult_PRFDest(decode_writeBackResult_PRFDest),
    .writeBackResult_data(decode_writeBackResult_data),
    .writeAddrPRF_exec1Addr(decode_writeAddrPRF_exec1Addr),
    .writeAddrPRF_exec2Addr(decode_writeAddrPRF_exec2Addr),
    .writeAddrPRF_exec3Addr(decode_writeAddrPRF_exec3Addr),
    .writeAddrPRF_exec1Valid(decode_writeAddrPRF_exec1Valid),
    .writeAddrPRF_exec2Valid(decode_writeAddrPRF_exec2Valid),
    .writeAddrPRF_exec3Valid(decode_writeAddrPRF_exec3Valid),
    .jumpAddrWrite_ready(decode_jumpAddrWrite_ready),
    .jumpAddrWrite_fired(decode_jumpAddrWrite_fired),
    .jumpAddrWrite_PRFDest(decode_jumpAddrWrite_PRFDest),
    .jumpAddrWrite_linkAddr(decode_jumpAddrWrite_linkAddr),
    .branchPCs_branchPCReady(decode_branchPCs_branchPCReady),
    .branchPCs_branchPC(decode_branchPCs_branchPC),
    .branchPCs_predictedPCReady(decode_branchPCs_predictedPCReady),
    .branchPCs_predictedPC(decode_branchPCs_predictedPC),
    .branchPCs_branchMask(decode_branchPCs_branchMask),
    .branchEvalIn_fired(decode_branchEvalIn_fired),
    .branchEvalIn_passFail(decode_branchEvalIn_passFail),
    .branchEvalIn_branchMask(decode_branchEvalIn_branchMask),
    .branchEvalIn_targetPC(decode_branchEvalIn_targetPC),
    .interruptedPC(decode_interruptedPC),
    .canTakeInterrupt(decode_canTakeInterrupt)
  );
  storeDataIssue dataQueue ( // @[core.scala 73:25]
    .clock(dataQueue_clock),
    .reset(dataQueue_reset),
    .fromROB_readyNow(dataQueue_fromROB_readyNow),
    .fromBranch_passOrFail(dataQueue_fromBranch_passOrFail),
    .fromBranch_robAddr(dataQueue_fromBranch_robAddr),
    .fromBranch_valid(dataQueue_fromBranch_valid),
    .fromDecode_ready(dataQueue_fromDecode_ready),
    .fromDecode_valid(dataQueue_fromDecode_valid),
    .fromDecode_rs2Addr(dataQueue_fromDecode_rs2Addr),
    .fromDecode_branchMask(dataQueue_fromDecode_branchMask),
    .toPRF_valid(dataQueue_toPRF_valid),
    .toPRF_rs2Addr(dataQueue_toPRF_rs2Addr),
    .robMapUpdate_valid(dataQueue_robMapUpdate_valid),
    .robMapUpdate_robAddr(dataQueue_robMapUpdate_robAddr)
  );
  rob rob ( // @[core.scala 74:19]
    .clock(rob_clock),
    .reset(rob_reset),
    .allocate_ready(rob_allocate_ready),
    .allocate_fired(rob_allocate_fired),
    .allocate_pc(rob_allocate_pc),
    .allocate_instruction(rob_allocate_instruction),
    .allocate_prfDest(rob_allocate_prfDest),
    .allocate_robAddr(rob_allocate_robAddr),
    .allocate_isReady(rob_allocate_isReady),
    .commit_ready(rob_commit_ready),
    .commit_fired(rob_commit_fired),
    .commit_prfDest(rob_commit_prfDest),
    .commit_pc(rob_commit_pc),
    .commit_instruction(rob_commit_instruction),
    .commit_exceptionOccurred(rob_commit_exceptionOccurred),
    .commit_mtval(rob_commit_mtval),
    .commit_isStore(rob_commit_isStore),
    .commit_is_fence(rob_commit_is_fence),
    .commit_robAddr(rob_commit_robAddr),
    .branch_valid(rob_branch_valid),
    .branch_pass(rob_branch_pass),
    .branch_robAddr(rob_branch_robAddr),
    .execPorts_0_robAddr(rob_execPorts_0_robAddr),
    .execPorts_0_mtval(rob_execPorts_0_mtval),
    .execPorts_0_valid(rob_execPorts_0_valid),
    .execPorts_1_robAddr(rob_execPorts_1_robAddr),
    .execPorts_1_valid(rob_execPorts_1_valid),
    .execPorts_2_robAddr(rob_execPorts_2_robAddr),
    .execPorts_2_valid(rob_execPorts_2_valid),
    .execPorts_3_robAddr(rob_execPorts_3_robAddr),
    .execPorts_3_valid(rob_execPorts_3_valid)
  );
  scheduler scheduler ( // @[core.scala 75:25]
    .clock(scheduler_clock),
    .reset(scheduler_reset),
    .allocate_ready(scheduler_allocate_ready),
    .allocate_fired(scheduler_allocate_fired),
    .allocate_instruction(scheduler_allocate_instruction),
    .allocate_branchMask(scheduler_allocate_branchMask),
    .allocate_rs1_ready(scheduler_allocate_rs1_ready),
    .allocate_rs1_prfAddr(scheduler_allocate_rs1_prfAddr),
    .allocate_rs2_ready(scheduler_allocate_rs2_ready),
    .allocate_rs2_prfAddr(scheduler_allocate_rs2_prfAddr),
    .allocate_prfDest(scheduler_allocate_prfDest),
    .allocate_robAddr(scheduler_allocate_robAddr),
    .release_ready(scheduler_release_ready),
    .release_fired(scheduler_release_fired),
    .release_instruction(scheduler_release_instruction),
    .release_branchMask(scheduler_release_branchMask),
    .release_rs1prfAddr(scheduler_release_rs1prfAddr),
    .release_rs2prfAddr(scheduler_release_rs2prfAddr),
    .release_prfDest(scheduler_release_prfDest),
    .release_robAddr(scheduler_release_robAddr),
    .wakeUpExt_0_valid(scheduler_wakeUpExt_0_valid),
    .wakeUpExt_0_prfAddr(scheduler_wakeUpExt_0_prfAddr),
    .wakeUpExt_1_valid(scheduler_wakeUpExt_1_valid),
    .wakeUpExt_1_prfAddr(scheduler_wakeUpExt_1_prfAddr),
    .branchOps_valid(scheduler_branchOps_valid),
    .branchOps_branchMask(scheduler_branchOps_branchMask),
    .branchOps_passed(scheduler_branchOps_passed),
    .memoryReady(scheduler_memoryReady),
    .multuplyAndDivideReady(scheduler_multuplyAndDivideReady),
    .instrRetired_valid(scheduler_instrRetired_valid),
    .instrRetired_prfAddr(scheduler_instrRetired_prfAddr)
  );
  core_Anon_1 memAccess ( // @[core.scala 76:25]
    .clock(memAccess_clock),
    .reset(memAccess_reset),
    .request_valid(memAccess_request_valid),
    .request_address(memAccess_request_address),
    .request_instruction(memAccess_request_instruction),
    .request_branchMask(memAccess_request_branchMask),
    .request_robAddr(memAccess_request_robAddr),
    .request_prfDest(memAccess_request_prfDest),
    .dPort_AWADDR(memAccess_dPort_AWADDR),
    .dPort_AWVALID(memAccess_dPort_AWVALID),
    .dPort_AWREADY(memAccess_dPort_AWREADY),
    .dPort_WDATA(memAccess_dPort_WDATA),
    .dPort_WLAST(memAccess_dPort_WLAST),
    .dPort_WVALID(memAccess_dPort_WVALID),
    .dPort_WREADY(memAccess_dPort_WREADY),
    .dPort_BRESP(memAccess_dPort_BRESP),
    .dPort_BVALID(memAccess_dPort_BVALID),
    .dPort_BREADY(memAccess_dPort_BREADY),
    .dPort_ARADDR(memAccess_dPort_ARADDR),
    .dPort_ARVALID(memAccess_dPort_ARVALID),
    .dPort_ARREADY(memAccess_dPort_ARREADY),
    .dPort_RDATA(memAccess_dPort_RDATA),
    .dPort_RLAST(memAccess_dPort_RLAST),
    .dPort_RVALID(memAccess_dPort_RVALID),
    .dPort_RREADY(memAccess_dPort_RREADY),
    .dPort_AWSNOOP(memAccess_dPort_AWSNOOP),
    .dPort_ARSNOOP(memAccess_dPort_ARSNOOP),
    .dPort_RRESP(memAccess_dPort_RRESP),
    .dPort_ACVALID(memAccess_dPort_ACVALID),
    .dPort_ACREADY(memAccess_dPort_ACREADY),
    .dPort_ACADDR(memAccess_dPort_ACADDR),
    .dPort_ACSNOOP(memAccess_dPort_ACSNOOP),
    .dPort_CRVALID(memAccess_dPort_CRVALID),
    .dPort_CRREADY(memAccess_dPort_CRREADY),
    .dPort_CRRESP(memAccess_dPort_CRRESP),
    .dPort_CDVALID(memAccess_dPort_CDVALID),
    .dPort_CDREADY(memAccess_dPort_CDREADY),
    .dPort_CDDATA(memAccess_dPort_CDDATA),
    .dPort_CDLAST(memAccess_dPort_CDLAST),
    .peripheral_AWADDR(memAccess_peripheral_AWADDR),
    .peripheral_AWLEN(memAccess_peripheral_AWLEN),
    .peripheral_AWSIZE(memAccess_peripheral_AWSIZE),
    .peripheral_AWBURST(memAccess_peripheral_AWBURST),
    .peripheral_AWPROT(memAccess_peripheral_AWPROT),
    .peripheral_AWVALID(memAccess_peripheral_AWVALID),
    .peripheral_AWREADY(memAccess_peripheral_AWREADY),
    .peripheral_WDATA(memAccess_peripheral_WDATA),
    .peripheral_WSTRB(memAccess_peripheral_WSTRB),
    .peripheral_WLAST(memAccess_peripheral_WLAST),
    .peripheral_WVALID(memAccess_peripheral_WVALID),
    .peripheral_WREADY(memAccess_peripheral_WREADY),
    .peripheral_BID(memAccess_peripheral_BID),
    .peripheral_BRESP(memAccess_peripheral_BRESP),
    .peripheral_BVALID(memAccess_peripheral_BVALID),
    .peripheral_BREADY(memAccess_peripheral_BREADY),
    .peripheral_ARADDR(memAccess_peripheral_ARADDR),
    .peripheral_ARLEN(memAccess_peripheral_ARLEN),
    .peripheral_ARSIZE(memAccess_peripheral_ARSIZE),
    .peripheral_ARBURST(memAccess_peripheral_ARBURST),
    .peripheral_ARPROT(memAccess_peripheral_ARPROT),
    .peripheral_ARVALID(memAccess_peripheral_ARVALID),
    .peripheral_ARREADY(memAccess_peripheral_ARREADY),
    .peripheral_RID(memAccess_peripheral_RID),
    .peripheral_RDATA(memAccess_peripheral_RDATA),
    .peripheral_RRESP(memAccess_peripheral_RRESP),
    .peripheral_RLAST(memAccess_peripheral_RLAST),
    .peripheral_RVALID(memAccess_peripheral_RVALID),
    .peripheral_RREADY(memAccess_peripheral_RREADY),
    .responseOut_valid(memAccess_responseOut_valid),
    .responseOut_prfDest(memAccess_responseOut_prfDest),
    .responseOut_robAddr(memAccess_responseOut_robAddr),
    .responseOut_result(memAccess_responseOut_result),
    .responseOut_instruction(memAccess_responseOut_instruction),
    .canAllocate(memAccess_canAllocate),
    .writeDataIn_valid(memAccess_writeDataIn_valid),
    .writeDataIn_data(memAccess_writeDataIn_data),
    .initiateFence(memAccess_initiateFence),
    .fenceInstructions_ready(memAccess_fenceInstructions_ready),
    .fenceInstructions_fired(memAccess_fenceInstructions_fired),
    .writeCommit_ready(memAccess_writeCommit_ready),
    .writeCommit_fired(memAccess_writeCommit_fired),
    .writeInstructionCommit_ready(memAccess_writeInstructionCommit_ready),
    .writeInstructionCommit_fired(memAccess_writeInstructionCommit_fired),
    .branchOps_valid(memAccess_branchOps_valid),
    .branchOps_branchMask(memAccess_branchOps_branchMask),
    .branchOps_passed(memAccess_branchOps_passed),
    .loadCommit_ready(memAccess_loadCommit_ready),
    .loadCommit_valid(memAccess_loadCommit_valid),
    .loadCommit_state(memAccess_loadCommit_state)
  );
  PRF prf ( // @[core.scala 143:19]
    .clock(prf_clock),
    .reset(prf_reset),
    .w1_addr(prf_w1_addr),
    .w1_data(prf_w1_data),
    .w1_en(prf_w1_en),
    .w2_addr(prf_w2_addr),
    .w2_data(prf_w2_data),
    .w2_en(prf_w2_en),
    .w3_addr(prf_w3_addr),
    .w3_data(prf_w3_data),
    .w3_en(prf_w3_en),
    .w4_addr(prf_w4_addr),
    .w4_data(prf_w4_data),
    .w4_en(prf_w4_en),
    .execRead_valid(prf_execRead_valid),
    .execRead_instruction(prf_execRead_instruction),
    .execRead_branchmask(prf_execRead_branchmask),
    .execRead_rs1Addr(prf_execRead_rs1Addr),
    .execRead_rs2Addr(prf_execRead_rs2Addr),
    .execRead_robAddr(prf_execRead_robAddr),
    .execRead_prfDest(prf_execRead_prfDest),
    .toExec_valid(prf_toExec_valid),
    .toExec_instruction(prf_toExec_instruction),
    .toExec_branchmask(prf_toExec_branchmask),
    .toExec_rs1Addr(prf_toExec_rs1Addr),
    .toExec_rs1Data(prf_toExec_rs1Data),
    .toExec_rs2Addr(prf_toExec_rs2Addr),
    .toExec_rs2Data(prf_toExec_rs2Data),
    .toExec_robAddr(prf_toExec_robAddr),
    .toExec_prfDest(prf_toExec_prfDest),
    .fromStore_valid(prf_fromStore_valid),
    .fromStore_rs2Addr(prf_fromStore_rs2Addr),
    .toStore_valid(prf_toStore_valid),
    .toStore_rs2Data(prf_toStore_rs2Data),
    .branchCheck_pass(prf_branchCheck_pass),
    .branchCheck_branchmask(prf_branchCheck_branchmask),
    .branchCheck_valid(prf_branchCheck_valid)
  );
  assign iPort_ARADDR = icache_lowLevelMem_ARADDR; // @[core.scala 31:9]
  assign iPort_ARVALID = icache_lowLevelMem_ARVALID; // @[core.scala 31:9]
  assign iPort_RREADY = icache_lowLevelMem_RREADY; // @[core.scala 31:9]
  assign debug_probe_arvalid_internal = icache_debug_probe_arvalid_internal; // @[core.scala 35:9]
  assign debug_probe_cacheMissed = icache_debug_probe_cacheMissed; // @[core.scala 35:9]
  assign debug_probe_rready_signal = icache_debug_probe_rready_signal; // @[core.scala 35:9]
  assign debug_probe_cacheFill_valid = icache_debug_probe_cacheFill_valid; // @[core.scala 35:9]
  assign debug_probe_axi_arvalid = icache_debug_probe_axi_arvalid; // @[core.scala 35:9]
  assign debug_probe_axi_arready = icache_debug_probe_axi_arready; // @[core.scala 35:9]
  assign debug_probe_req_valid = icache_debug_probe_req_valid; // @[core.scala 35:9]
  assign debug_probe_req_pc = icache_debug_probe_req_pc; // @[core.scala 35:9]
  assign fdbg_probe_redirect_bit = fetch_fdbg_probe_redirect_bit; // @[core.scala 50:8]
  assign fdbg_probe_fifo_enq_ready = fetch_fdbg_probe_fifo_enq_ready; // @[core.scala 50:8]
  assign fdbg_probe_is_fence = fetch_fdbg_probe_is_fence; // @[core.scala 50:8]
  assign fdbg_probe_handle_fence = fetch_fdbg_probe_handle_fence; // @[core.scala 50:8]
  assign dPort_AWADDR = memAccess_dPort_AWADDR; // @[core.scala 846:9]
  assign dPort_AWVALID = memAccess_dPort_AWVALID; // @[core.scala 846:9]
  assign dPort_WDATA = memAccess_dPort_WDATA; // @[core.scala 846:9]
  assign dPort_WLAST = memAccess_dPort_WLAST; // @[core.scala 846:9]
  assign dPort_WVALID = memAccess_dPort_WVALID; // @[core.scala 846:9]
  assign dPort_BREADY = memAccess_dPort_BREADY; // @[core.scala 846:9]
  assign dPort_ARADDR = memAccess_dPort_ARADDR; // @[core.scala 846:9]
  assign dPort_ARVALID = memAccess_dPort_ARVALID; // @[core.scala 846:9]
  assign dPort_RREADY = memAccess_dPort_RREADY; // @[core.scala 846:9]
  assign dPort_AWSNOOP = memAccess_dPort_AWSNOOP; // @[core.scala 846:9]
  assign dPort_ARSNOOP = memAccess_dPort_ARSNOOP; // @[core.scala 846:9]
  assign dPort_ACREADY = memAccess_dPort_ACREADY; // @[core.scala 846:9]
  assign dPort_CRVALID = memAccess_dPort_CRVALID; // @[core.scala 846:9]
  assign dPort_CRRESP = memAccess_dPort_CRRESP; // @[core.scala 846:9]
  assign dPort_CDVALID = memAccess_dPort_CDVALID; // @[core.scala 846:9]
  assign dPort_CDDATA = memAccess_dPort_CDDATA; // @[core.scala 846:9]
  assign dPort_CDLAST = memAccess_dPort_CDLAST; // @[core.scala 846:9]
  assign peripheral_AWADDR = memAccess_peripheral_AWADDR; // @[core.scala 847:14]
  assign peripheral_AWLEN = memAccess_peripheral_AWLEN; // @[core.scala 847:14]
  assign peripheral_AWSIZE = memAccess_peripheral_AWSIZE; // @[core.scala 847:14]
  assign peripheral_AWBURST = memAccess_peripheral_AWBURST; // @[core.scala 847:14]
  assign peripheral_AWPROT = memAccess_peripheral_AWPROT; // @[core.scala 847:14]
  assign peripheral_AWVALID = memAccess_peripheral_AWVALID; // @[core.scala 847:14]
  assign peripheral_WDATA = memAccess_peripheral_WDATA; // @[core.scala 847:14]
  assign peripheral_WSTRB = memAccess_peripheral_WSTRB; // @[core.scala 847:14]
  assign peripheral_WLAST = memAccess_peripheral_WLAST; // @[core.scala 847:14]
  assign peripheral_WVALID = memAccess_peripheral_WVALID; // @[core.scala 847:14]
  assign peripheral_BREADY = memAccess_peripheral_BREADY; // @[core.scala 847:14]
  assign peripheral_ARADDR = memAccess_peripheral_ARADDR; // @[core.scala 847:14]
  assign peripheral_ARLEN = memAccess_peripheral_ARLEN; // @[core.scala 847:14]
  assign peripheral_ARSIZE = memAccess_peripheral_ARSIZE; // @[core.scala 847:14]
  assign peripheral_ARBURST = memAccess_peripheral_ARBURST; // @[core.scala 847:14]
  assign peripheral_ARPROT = memAccess_peripheral_ARPROT; // @[core.scala 847:14]
  assign peripheral_ARVALID = memAccess_peripheral_ARVALID; // @[core.scala 847:14]
  assign peripheral_RREADY = memAccess_peripheral_RREADY; // @[core.scala 847:14]
  assign core_sample0 = decode_fromFetch_expected_valid; // @[core.scala 995:16]
  assign core_sample1 = decode_fromFetch_expected_pc[30]; // @[core.scala 996:47]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_fromFetch_req_valid = fetch_cache_req_valid; // @[core.scala 44:24]
  assign icache_fromFetch_req_bits = {32'h0,fetch_cache_req_bits[31:0]}; // @[Cat.scala 33:92]
  assign icache_fromFetch_resp_ready = fetch_cache_resp_ready; // @[core.scala 46:20]
  assign icache_updateAllCachelines_fired = memAccess_fenceInstructions_ready & icache_updateAllCachelines_ready; // @[core.scala 901:45]
  assign icache_cachelinesUpdatesResp_fired = icache_cachelinesUpdatesResp_ready & fetch_cachelinesUpdatesResp_ready; // @[core.scala 911:46]
  assign icache_lowLevelMem_ARREADY = iPort_ARREADY; // @[core.scala 31:9]
  assign icache_lowLevelMem_RDATA = iPort_RDATA; // @[core.scala 31:9]
  assign icache_lowLevelMem_RLAST = iPort_RLAST; // @[core.scala 31:9]
  assign icache_lowLevelMem_RVALID = iPort_RVALID; // @[core.scala 31:9]
  assign fetch_clock = clock;
  assign fetch_reset = reset;
  assign fetch_cache_req_ready = icache_fromFetch_req_ready; // @[core.scala 44:24]
  assign fetch_cache_resp_valid = icache_fromFetch_resp_valid; // @[core.scala 46:20]
  assign fetch_cache_resp_bits = icache_fromFetch_resp_bits; // @[core.scala 46:20]
  assign fetch_toDecode_fired = ~(interruptInjectStatus == 2'h0 | interruptInjectStatus == 2'h1 & ~_T_231) ? 1'h0 :
    decode_fromFetch_ready & fetch_toDecode_ready & _fetch_toDecode_fired_T_3; // @[core.scala 1114:126 1116:26 65:7]
  assign fetch_toDecode_expected_valid = decode_fromFetch_expected_valid; // @[core.scala 69:27]
  assign fetch_toDecode_expected_pc = decode_fromFetch_expected_pc; // @[core.scala 69:27]
  assign fetch_toDecode_expected_coherency = decode_fromFetch_expected_coherency; // @[core.scala 69:27]
  assign fetch_branchRes_fired = branchEvals_valid & ~coherentLoadInvalidReg; // @[core.scala 716:71]
  assign fetch_branchRes_branchTaken = 3'h7 == branchInstruction_instruction[14:12] ? branchTaken_conditionEval_7 :
    _GEN_220; // @[core.scala 712:{31,31}]
  assign fetch_branchRes_pc = branchPCs_0_pc; // @[core.scala 714:22]
  assign fetch_branchRes_pcAfterBrnach = branchEvals_nextPC; // @[core.scala 715:33]
  assign fetch_carryOutFence_fired = fetch_carryOutFence_ready; // @[core.scala 903:29]
  assign fetch_updateAllCachelines_fired = fetch_updateAllCachelines_ready; // @[core.scala 908:35]
  assign fetch_cachelinesUpdatesResp_fired = icache_cachelinesUpdatesResp_ready & fetch_cachelinesUpdatesResp_ready; // @[core.scala 911:46]
  assign decode_clock = clock;
  assign decode_reset = reset;
  assign decode_fromFetch_fired = ~(interruptInjectStatus == 2'h0 | interruptInjectStatus == 2'h1 & ~_T_231) ? 1'h0 :
    decode_fromFetch_ready & fetch_toDecode_ready & _fetch_toDecode_fired_T_3; // @[core.scala 1114:126 1117:28 65:7]
  assign decode_fromFetch_pc = fetch_toDecode_pc; // @[core.scala 71:23]
  assign decode_fromFetch_instruction = _GEN_299[31:0];
  assign decode_toExec_fired = decode_toExec_ready & rob_allocate_ready & scheduler_allocate_ready & (
    decode_toExec_instruction[6:4] != 3'h2 | dataQueue_fromDecode_ready); // @[core.scala 103:81]
  assign decode_writeBackResult_fired = (~_coherentLoadInvalid_T_5 | ~coherentLoadInvalid & memAccess_loadCommit_valid)
     & rob_commit_ready & (memAccess_writeInstructionCommit_ready | rob_commit_instruction[6:4] != 3'h2); // @[core.scala 725:160]
  assign decode_writeBackResult_instruction = _GEN_300[31:0];
  assign decode_writeBackResult_rdAddr = rob_commit_instruction[11:7]; // @[core.scala 721:58]
  assign decode_writeBackResult_PRFDest = rob_commit_prfDest; // @[core.scala 718:34]
  assign decode_writeBackResult_data = rob_commit_mtval; // @[core.scala 915:31]
  assign decode_writeAddrPRF_exec1Addr = scheduler_instrRetired_prfAddr; // @[core.scala 736:33]
  assign decode_writeAddrPRF_exec2Addr = memAccess_responseOut_prfDest; // @[core.scala 738:33]
  assign decode_writeAddrPRF_exec3Addr = extnMResponse_prfDest; // @[core.scala 739:33]
  assign decode_writeAddrPRF_exec1Valid = scheduler_instrRetired_valid; // @[core.scala 737:34]
  assign decode_writeAddrPRF_exec2Valid = memAccess_responseOut_valid & _T_181; // @[core.scala 740:65]
  assign decode_writeAddrPRF_exec3Valid = extnMResponse_valid & _T_184; // @[core.scala 741:57]
  assign decode_jumpAddrWrite_fired = decode_jumpAddrWrite_ready; // @[core.scala 807:30]
  assign decode_branchEvalIn_fired = branchEvals_valid; // @[core.scala 746:58]
  assign decode_branchEvalIn_passFail = branchEvals_passed; // @[core.scala 744:32]
  assign decode_branchEvalIn_branchMask = branchEvals_branchMask; // @[core.scala 743:34]
  assign decode_branchEvalIn_targetPC = branchEvals_nextPC; // @[core.scala 745:32]
  assign decode_interruptedPC = lastBranchExecPC; // @[core.scala 1053:24]
  assign dataQueue_clock = clock;
  assign dataQueue_reset = reset;
  assign dataQueue_fromROB_readyNow = memAccess_writeCommit_fired; // @[core.scala 826:30]
  assign dataQueue_fromBranch_passOrFail = branchEvals_passed; // @[core.scala 542:20 89:23]
  assign dataQueue_fromBranch_robAddr = branchEvals_robAddr; // @[core.scala 819:32]
  assign dataQueue_fromBranch_valid = branchEvals_valid; // @[core.scala 541:19 89:23]
  assign dataQueue_fromDecode_valid = branchEvals_valid ? _GEN_3 : scheduler_allocate_fired & decode_toExec_instruction[
    6:4] == 3'h2; // @[core.scala 124:25 122:30]
  assign dataQueue_fromDecode_rs2Addr = decode_toExec_rs2Addr; // @[core.scala 120:32]
  assign dataQueue_fromDecode_branchMask = branchEvals_valid ? _scheduler_allocate_branchMask_T :
    decode_toExec_branchMask; // @[core.scala 124:25 118:35 126:36]
  assign dataQueue_robMapUpdate_valid = rob_allocate_fired; // @[core.scala 824:32]
  assign dataQueue_robMapUpdate_robAddr = rob_allocate_robAddr; // @[core.scala 823:34]
  assign rob_clock = clock;
  assign rob_reset = reset;
  assign rob_allocate_fired = branchEvals_valid ? _GEN_2 : decode_toExec_ready & rob_allocate_ready &
    scheduler_allocate_ready & (decode_toExec_instruction[6:4] != 3'h2 | dataQueue_fromDecode_ready); // @[core.scala 124:25 103:7]
  assign rob_allocate_pc = decode_toExec_pc; // @[core.scala 106:19]
  assign rob_allocate_instruction = decode_toExec_instruction; // @[core.scala 107:28]
  assign rob_allocate_prfDest = decode_toExec_PRFDest; // @[core.scala 108:24]
  assign rob_allocate_isReady = 5'h3 == decode_toExec_instruction[6:2] | 5'h5 == decode_toExec_instruction[6:2] | 5'hd
     == decode_toExec_instruction[6:2]; // @[core.scala 101:125]
  assign rob_commit_fired = (~_coherentLoadInvalid_T_5 | ~coherentLoadInvalid & memAccess_loadCommit_valid) &
    rob_commit_ready & (memAccess_writeInstructionCommit_ready | rob_commit_instruction[6:4] != 3'h2); // @[core.scala 725:160]
  assign rob_branch_valid = branchEvals_valid; // @[core.scala 750:20]
  assign rob_branch_pass = branchEvals_passed; // @[core.scala 748:19]
  assign rob_branch_robAddr = branchEvals_robAddr; // @[core.scala 749:22]
  assign rob_execPorts_0_robAddr = singleCycleArithmeticResponse_robAddr; // @[core.scala 774:22]
  assign rob_execPorts_0_mtval = rob_execPorts_0_mtval_REG; // @[core.scala 758:26]
  assign rob_execPorts_0_valid = singleCycleArithmeticResponse_valid; // @[core.scala 775:20]
  assign rob_execPorts_1_robAddr = branchEvals_robAddr; // @[core.scala 774:22]
  assign rob_execPorts_1_valid = branchEvals_valid; // @[core.scala 775:20]
  assign rob_execPorts_2_robAddr = memAccess_responseOut_robAddr; // @[core.scala 774:22]
  assign rob_execPorts_2_valid = memAccess_responseOut_valid; // @[core.scala 775:20]
  assign rob_execPorts_3_robAddr = extnMResponse_robAddr; // @[core.scala 774:22]
  assign rob_execPorts_3_valid = extnMResponse_valid; // @[core.scala 775:20]
  assign scheduler_clock = clock;
  assign scheduler_reset = reset;
  assign scheduler_allocate_fired = branchEvals_valid ? _GEN_1 : _GEN_0; // @[core.scala 124:25]
  assign scheduler_allocate_instruction = decode_toExec_instruction; // @[core.scala 110:34]
  assign scheduler_allocate_branchMask = branchEvals_valid ? _scheduler_allocate_branchMask_T : decode_toExec_branchMask
    ; // @[core.scala 124:25 111:33 125:34]
  assign scheduler_allocate_rs1_ready = wakeUps_2_valid ? _GEN_17 : _GEN_15; // @[core.scala 135:24]
  assign scheduler_allocate_rs1_prfAddr = decode_toExec_rs1Addr; // @[core.scala 113:34]
  assign scheduler_allocate_rs2_ready = wakeUps_2_valid ? _GEN_18 : _GEN_16; // @[core.scala 135:24]
  assign scheduler_allocate_rs2_prfAddr = decode_toExec_rs2Addr; // @[core.scala 115:34]
  assign scheduler_allocate_prfDest = decode_toExec_PRFDest; // @[core.scala 116:30]
  assign scheduler_allocate_robAddr = rob_allocate_robAddr; // @[core.scala 117:30]
  assign scheduler_release_fired = scheduler_release_ready & _scheduler_release_fired_T_5; // @[core.scala 145:29]
  assign scheduler_wakeUpExt_0_valid = memAccess_responseOut_valid & |memAccess_responseOut_instruction[11:7]; // @[core.scala 798:33]
  assign scheduler_wakeUpExt_0_prfAddr = memAccess_responseOut_prfDest; // @[core.scala 803:20 95:21]
  assign scheduler_wakeUpExt_1_valid = extnMResponse_valid & |extnResponseInstruction[11:7]; // @[core.scala 799:25]
  assign scheduler_wakeUpExt_1_prfAddr = extnMResponse_prfDest; // @[core.scala 803:20 95:21]
  assign scheduler_branchOps_valid = branchEvals_valid; // @[core.scala 541:19 89:23]
  assign scheduler_branchOps_branchMask = branchEvals_branchMask; // @[core.scala 89:23 543:24]
  assign scheduler_branchOps_passed = branchEvals_passed; // @[core.scala 542:20 89:23]
  assign scheduler_memoryReady = memAccess_canAllocate; // @[core.scala 752:25]
  assign scheduler_multuplyAndDivideReady = mExtensionReady; // @[core.scala 753:36]
  assign memAccess_clock = clock;
  assign memAccess_reset = reset;
  assign memAccess_request_valid = memoryRequest_valid; // @[core.scala 206:21]
  assign memAccess_request_address = memoryRequest_address; // @[core.scala 206:21]
  assign memAccess_request_instruction = memoryRequest_instruction; // @[core.scala 206:21]
  assign memAccess_request_branchMask = memoryRequest_branchMask; // @[core.scala 206:21]
  assign memAccess_request_robAddr = memoryRequest_robAddr; // @[core.scala 206:21]
  assign memAccess_request_prfDest = memoryRequest_prfDest; // @[core.scala 206:21]
  assign memAccess_dPort_AWREADY = dPort_AWREADY; // @[core.scala 846:9]
  assign memAccess_dPort_WREADY = dPort_WREADY; // @[core.scala 846:9]
  assign memAccess_dPort_BRESP = dPort_BRESP; // @[core.scala 846:9]
  assign memAccess_dPort_BVALID = dPort_BVALID; // @[core.scala 846:9]
  assign memAccess_dPort_ARREADY = dPort_ARREADY; // @[core.scala 846:9]
  assign memAccess_dPort_RDATA = dPort_RDATA; // @[core.scala 846:9]
  assign memAccess_dPort_RLAST = dPort_RLAST; // @[core.scala 846:9]
  assign memAccess_dPort_RVALID = dPort_RVALID; // @[core.scala 846:9]
  assign memAccess_dPort_RRESP = dPort_RRESP; // @[core.scala 846:9]
  assign memAccess_dPort_ACVALID = dPort_ACVALID; // @[core.scala 846:9]
  assign memAccess_dPort_ACADDR = dPort_ACADDR; // @[core.scala 846:9]
  assign memAccess_dPort_ACSNOOP = dPort_ACSNOOP; // @[core.scala 846:9]
  assign memAccess_dPort_CRREADY = dPort_CRREADY; // @[core.scala 846:9]
  assign memAccess_dPort_CDREADY = dPort_CDREADY; // @[core.scala 846:9]
  assign memAccess_peripheral_AWREADY = peripheral_AWREADY; // @[core.scala 847:14]
  assign memAccess_peripheral_WREADY = peripheral_WREADY; // @[core.scala 847:14]
  assign memAccess_peripheral_BID = {{1'd0}, peripheral_BID}; // @[core.scala 847:14]
  assign memAccess_peripheral_BRESP = peripheral_BRESP; // @[core.scala 847:14]
  assign memAccess_peripheral_BVALID = peripheral_BVALID; // @[core.scala 847:14]
  assign memAccess_peripheral_ARREADY = peripheral_ARREADY; // @[core.scala 847:14]
  assign memAccess_peripheral_RID = {{1'd0}, peripheral_RID}; // @[core.scala 847:14]
  assign memAccess_peripheral_RDATA = peripheral_RDATA; // @[core.scala 847:14]
  assign memAccess_peripheral_RRESP = peripheral_RRESP; // @[core.scala 847:14]
  assign memAccess_peripheral_RLAST = peripheral_RLAST; // @[core.scala 847:14]
  assign memAccess_peripheral_RVALID = peripheral_RVALID; // @[core.scala 847:14]
  assign memAccess_writeDataIn_valid = prf_toStore_valid; // @[core.scala 829:31]
  assign memAccess_writeDataIn_data = prf_toStore_rs2Data; // @[core.scala 828:30]
  assign memAccess_initiateFence = REG_1 | _GEN_244; // @[core.scala 920:131 921:29]
  assign memAccess_fenceInstructions_fired = memAccess_fenceInstructions_ready & icache_updateAllCachelines_ready; // @[core.scala 901:45]
  assign memAccess_writeCommit_fired = memAccess_writeCommit_ready & _memAccess_writeInstructionCommit_fired_T_1; // @[core.scala 831:62]
  assign memAccess_writeInstructionCommit_fired = memAccess_writeInstructionCommit_ready & rob_commit_instruction[6:4]
     == 3'h2 & rob_commit_fired; // @[core.scala 728:132]
  assign memAccess_branchOps_valid = branchEvals_valid; // @[core.scala 541:19 89:23]
  assign memAccess_branchOps_branchMask = branchEvals_branchMask; // @[core.scala 89:23 543:24]
  assign memAccess_branchOps_passed = branchEvals_passed; // @[core.scala 542:20 89:23]
  assign memAccess_loadCommit_ready = _coherentLoadInvalid_T_5 & rob_commit_ready; // @[core.scala 731:71]
  assign prf_clock = clock;
  assign prf_reset = reset;
  assign prf_w1_addr = singleCycleArithmeticResponse_prfDest; // @[core.scala 786:20]
  assign prf_w1_data = singleCycleArithmeticResponse_result; // @[core.scala 787:20]
  assign prf_w1_en = singleCycleArithmeticResponse_valid & REG; // @[core.scala 779:119]
  assign prf_w2_addr = decode_jumpAddrWrite_PRFDest; // @[core.scala 786:20]
  assign prf_w2_data = decode_jumpAddrWrite_linkAddr; // @[core.scala 787:20]
  assign prf_w2_en = decode_jumpAddrWrite_ready; // @[core.scala 788:18]
  assign prf_w3_addr = memAccess_responseOut_prfDest; // @[core.scala 786:20]
  assign prf_w3_data = memAccess_responseOut_result; // @[core.scala 787:20]
  assign prf_w3_en = memAccess_responseOut_valid & _T_181; // @[core.scala 781:95]
  assign prf_w4_addr = extnMResponse_prfDest; // @[core.scala 786:20]
  assign prf_w4_data = extnMResponse_result; // @[core.scala 787:20]
  assign prf_w4_en = extnMResponse_valid & _T_184; // @[core.scala 782:71]
  assign prf_execRead_valid = scheduler_release_instruction[4:2] == 3'h2 ? 1'h0 : _GEN_21; // @[core.scala 926:{63,84}]
  assign prf_execRead_instruction = scheduler_release_instruction; // @[core.scala 149:28]
  assign prf_execRead_branchmask = scheduler_release_branchMask; // @[core.scala 150:27]
  assign prf_execRead_rs1Addr = scheduler_release_rs1prfAddr; // @[core.scala 151:24]
  assign prf_execRead_rs2Addr = scheduler_release_rs2prfAddr; // @[core.scala 152:24]
  assign prf_execRead_robAddr = {{2'd0}, scheduler_release_robAddr}; // @[core.scala 153:24]
  assign prf_execRead_prfDest = scheduler_release_prfDest; // @[core.scala 155:24]
  assign prf_fromStore_valid = prf_fromStore_valid_REG_1; // @[core.scala 816:23]
  assign prf_fromStore_rs2Addr = prf_fromStore_rs2Addr_REG_1; // @[core.scala 815:25]
  assign prf_branchCheck_pass = branchEvals_passed; // @[core.scala 542:20 89:23]
  assign prf_branchCheck_branchmask = branchEvals_branchMask; // @[core.scala 89:23 543:24]
  assign prf_branchCheck_valid = branchEvals_valid; // @[core.scala 541:19 89:23]
  always @(posedge clock) begin
    if (coherentLoadInvalid) begin // @[core.scala 573:32]
      branchEvals_branchMask <= 5'h10;
    end else begin
      branchEvals_branchMask <= branchPCs_0_branchMask;
    end
    if (2'h0 == interruptInjectStatus) begin // @[core.scala 1071:33]
      branchEvals_passed <= _branchEvals_passed_T_2; // @[core.scala 629:22]
    end else if (2'h1 == interruptInjectStatus) begin // @[core.scala 1071:33]
      if (decode_canTakeInterrupt) begin // @[core.scala 1079:56]
        if (~branchEvals_valid) begin // @[core.scala 1080:58]
          branchEvals_passed <= _GEN_278;
        end else begin
          branchEvals_passed <= _branchEvals_passed_T_2; // @[core.scala 629:22]
        end
      end else begin
        branchEvals_passed <= _branchEvals_passed_T_2; // @[core.scala 629:22]
      end
    end else begin
      branchEvals_passed <= _branchEvals_passed_T_2; // @[core.scala 629:22]
    end
    if (reset) begin // @[core.scala 534:28]
      branchEvals_valid <= 1'h0; // @[core.scala 534:28]
    end else if (branchEvals_valid) begin // @[core.scala 575:25]
      if (_T) begin // @[core.scala 577:29]
        branchEvals_valid <= 1'h0; // @[core.scala 578:25]
      end else begin
        branchEvals_valid <= coherentLoadInvalid | branchInstruction_valid; // @[core.scala 571:21]
      end
    end else begin
      branchEvals_valid <= coherentLoadInvalid | branchInstruction_valid; // @[core.scala 571:21]
    end
    if (division_request_valid & ~(|division_counter)) begin // @[core.scala 450:57]
      extnMResponse_prfDest <= division_request_prfDest; // @[core.scala 451:27]
    end else begin
      extnMResponse_prfDest <= extnMServicing_prfDest; // @[core.scala 376:25]
    end
    if (reset) begin // @[core.scala 235:30]
      extnMResponse_valid <= 1'h0; // @[core.scala 235:30]
    end else if (division_request_valid & ~(|division_counter)) begin // @[core.scala 450:57]
      if (branchEvals_valid) begin // @[core.scala 474:27]
        if (|_T_106 & _T) begin // @[core.scala 475:91]
          extnMResponse_valid <= 1'h0; // @[core.scala 475:113]
        end else begin
          extnMResponse_valid <= division_request_valid; // @[core.scala 471:25]
        end
      end else begin
        extnMResponse_valid <= division_request_valid; // @[core.scala 471:25]
      end
    end else if (branchEvals_valid) begin // @[core.scala 391:25]
      if (_T) begin // @[core.scala 397:29]
        extnMResponse_valid <= _GEN_67;
      end else begin
        extnMResponse_valid <= extnMServicing_valid; // @[core.scala 388:23]
      end
    end else begin
      extnMResponse_valid <= extnMServicing_valid; // @[core.scala 388:23]
    end
    if (division_request_valid & ~(|division_counter)) begin // @[core.scala 450:57]
      extnResponseInstruction <= division_request_instruction; // @[core.scala 472:29]
    end else begin
      extnResponseInstruction <= extnMServicing_instruction; // @[core.scala 389:27]
    end
    mExtensionReady <= reset | _GEN_85; // @[core.scala 141:{32,32}]
    if (reset) begin // @[core.scala 164:39]
      addressGenerationInput_valid <= 1'h0; // @[core.scala 164:39]
    end else if (branchEvals_valid) begin // @[core.scala 180:25]
      if (_T & _T_10) begin // @[core.scala 184:83]
        addressGenerationInput_valid <= 1'h0; // @[core.scala 184:114]
      end else begin
        addressGenerationInput_valid <= prf_toExec_valid & ~(prf_toExec_instruction[6] | prf_toExec_instruction[4]); // @[core.scala 173:32]
      end
    end else begin
      addressGenerationInput_valid <= prf_toExec_valid & ~(prf_toExec_instruction[6] | prf_toExec_instruction[4]); // @[core.scala 173:32]
    end
    if (|prf_toExec_instruction[19:15]) begin // @[core.scala 259:36]
      if (_addressGenerationInput_rs1_T_3) begin // @[Mux.scala 101:16]
        addressGenerationInput_rs1 <= fwdFrom_0_result;
      end else if (_addressGenerationInput_rs1_T_5) begin // @[Mux.scala 101:16]
        addressGenerationInput_rs1 <= fwdBuffers_0_result;
      end else if (_addressGenerationInput_rs1_T_7) begin // @[Mux.scala 101:16]
        addressGenerationInput_rs1 <= fwdBuffers_1_result;
      end else begin
        addressGenerationInput_rs1 <= prf_toExec_rs1Data;
      end
    end else begin
      addressGenerationInput_rs1 <= 64'h0;
    end
    addressGenerationInput_instruction <= prf_toExec_instruction; // @[core.scala 175:38]
    addressGenerationInput_prfDest <= prf_toExec_prfDest; // @[core.scala 176:34]
    addressGenerationInput_robAddr <= prf_toExec_robAddr[3:0]; // @[core.scala 177:34]
    if (branchEvals_valid) begin // @[core.scala 180:25]
      if (|_T_9) begin // @[core.scala 181:62]
        addressGenerationInput_branchMask <= _addressGenerationInput_branchMask_T; // @[core.scala 182:41]
      end else begin
        addressGenerationInput_branchMask <= prf_toExec_branchmask; // @[core.scala 178:37]
      end
    end else begin
      addressGenerationInput_branchMask <= prf_toExec_branchmask; // @[core.scala 178:37]
    end
    if (reset) begin // @[core.scala 187:30]
      memoryRequest_valid <= 1'h0; // @[core.scala 187:30]
    end else if (branchEvals_valid) begin // @[core.scala 199:25]
      if (_T & _T_16) begin // @[core.scala 203:95]
        memoryRequest_valid <= 1'h0; // @[core.scala 203:117]
      end else begin
        memoryRequest_valid <= addressGenerationInput_valid; // @[core.scala 197:23]
      end
    end else begin
      memoryRequest_valid <= addressGenerationInput_valid; // @[core.scala 197:23]
    end
    memoryRequest_address <= _memoryRequest_address_T_15[31:0]; // @[core.scala 188:25]
    memoryRequest_instruction <= addressGenerationInput_instruction; // @[core.scala 194:29]
    if (branchEvals_valid) begin // @[core.scala 199:25]
      if (|_T_15) begin // @[core.scala 200:74]
        memoryRequest_branchMask <= _memoryRequest_branchMask_T; // @[core.scala 201:32]
      end else begin
        memoryRequest_branchMask <= addressGenerationInput_branchMask; // @[core.scala 193:28]
      end
    end else begin
      memoryRequest_branchMask <= addressGenerationInput_branchMask; // @[core.scala 193:28]
    end
    memoryRequest_robAddr <= addressGenerationInput_robAddr; // @[core.scala 196:25]
    memoryRequest_prfDest <= addressGenerationInput_prfDest; // @[core.scala 195:25]
    if (reset) begin // @[core.scala 209:45]
      singleCycleArithmeticRequest_valid <= 1'h0; // @[core.scala 209:45]
    end else if (branchEvals_valid) begin // @[core.scala 310:25]
      if (_T_14) begin // @[core.scala 314:83]
        singleCycleArithmeticRequest_valid <= 1'h0; // @[core.scala 315:42]
      end else begin
        singleCycleArithmeticRequest_valid <= prf_toExec_valid & 3'h4 == _singleCycleArithmeticRequest_valid_T_1 & (
          prf_toExec_instruction[6] | ~prf_toExec_instruction[5] | ~prf_toExec_instruction[25]); // @[core.scala 298:38]
      end
    end else begin
      singleCycleArithmeticRequest_valid <= prf_toExec_valid & 3'h4 == _singleCycleArithmeticRequest_valid_T_1 & (
        prf_toExec_instruction[6] | ~prf_toExec_instruction[5] | ~prf_toExec_instruction[25]); // @[core.scala 298:38]
    end
    if (_addressGenerationInput_rs1_T_1) begin // @[core.scala 303:42]
      if (_addressGenerationInput_rs1_T_3) begin // @[Mux.scala 101:16]
        singleCycleArithmeticRequest_rs1 <= fwdFrom_0_result;
      end else if (_addressGenerationInput_rs1_T_5) begin // @[Mux.scala 101:16]
        singleCycleArithmeticRequest_rs1 <= fwdBuffers_0_result;
      end else if (_addressGenerationInput_rs1_T_7) begin // @[Mux.scala 101:16]
        singleCycleArithmeticRequest_rs1 <= fwdBuffers_1_result;
      end else begin
        singleCycleArithmeticRequest_rs1 <= prf_toExec_rs1Data;
      end
    end else begin
      singleCycleArithmeticRequest_rs1 <= 64'h0;
    end
    if (prf_toExec_instruction[5]) begin // @[core.scala 306:42]
      if (|prf_toExec_instruction[24:20]) begin // @[core.scala 306:80]
        if (_singleCycleArithmeticRequest_rs2_T_5) begin // @[Mux.scala 101:16]
          singleCycleArithmeticRequest_rs2 <= fwdFrom_0_result;
        end else if (_singleCycleArithmeticRequest_rs2_T_7) begin // @[Mux.scala 101:16]
          singleCycleArithmeticRequest_rs2 <= fwdBuffers_0_result;
        end else begin
          singleCycleArithmeticRequest_rs2 <= _singleCycleArithmeticRequest_rs2_T_10;
        end
      end else begin
        singleCycleArithmeticRequest_rs2 <= 64'h0;
      end
    end else begin
      singleCycleArithmeticRequest_rs2 <= arithmeticImm;
    end
    singleCycleArithmeticRequest_instruction <= prf_toExec_instruction; // @[core.scala 300:44]
    singleCycleArithmeticRequest_prfDest <= prf_toExec_prfDest; // @[core.scala 301:40]
    singleCycleArithmeticRequest_robAddr <= prf_toExec_robAddr[3:0]; // @[core.scala 302:40]
    if (branchEvals_valid) begin // @[core.scala 310:25]
      if (|_T_9) begin // @[core.scala 181:62]
        singleCycleArithmeticRequest_branchMask <= _addressGenerationInput_branchMask_T; // @[core.scala 182:41]
      end else begin
        singleCycleArithmeticRequest_branchMask <= prf_toExec_branchmask; // @[core.scala 178:37]
      end
    end else begin
      singleCycleArithmeticRequest_branchMask <= prf_toExec_branchmask; // @[core.scala 299:43]
    end
    if (reset) begin // @[core.scala 219:46]
      singleCycleArithmeticResponse_valid <= 1'h0; // @[core.scala 219:46]
    end else if (branchEvals_valid) begin // @[core.scala 325:25]
      if (_T & |_T_30) begin // @[core.scala 326:101]
        singleCycleArithmeticResponse_valid <= 1'h0; // @[core.scala 327:43]
      end else begin
        singleCycleArithmeticResponse_valid <= singleCycleArithmeticRequest_valid; // @[core.scala 323:39]
      end
    end else begin
      singleCycleArithmeticResponse_valid <= singleCycleArithmeticRequest_valid; // @[core.scala 323:39]
    end
    singleCycleArithmeticResponse_result <= arithmeticResult[63:0]; // @[core.scala 321:40]
    singleCycleArithmeticResponse_prfDest <= singleCycleArithmeticRequest_prfDest; // @[core.scala 320:41]
    singleCycleArithmeticResponse_robAddr <= singleCycleArithmeticRequest_robAddr; // @[core.scala 322:41]
    if (reset) begin // @[core.scala 226:29]
      extnMRequest_valid <= 1'h0; // @[core.scala 226:29]
    end else if (branchEvals_valid) begin // @[core.scala 391:25]
      if (_T) begin // @[core.scala 397:29]
        if (_T_10 & prf_toExec_valid) begin // @[core.scala 400:101]
          extnMRequest_valid <= 1'h0; // @[core.scala 400:107]
        end else begin
          extnMRequest_valid <= _GEN_56;
        end
      end else begin
        extnMRequest_valid <= _GEN_56;
      end
    end else begin
      extnMRequest_valid <= _GEN_56;
    end
    if (_addressGenerationInput_rs1_T_3) begin // @[Mux.scala 101:16]
      extnMRequest_rs1 <= fwdFrom_0_result;
    end else if (_addressGenerationInput_rs1_T_5) begin // @[Mux.scala 101:16]
      extnMRequest_rs1 <= fwdBuffers_0_result;
    end else if (_addressGenerationInput_rs1_T_7) begin // @[Mux.scala 101:16]
      extnMRequest_rs1 <= fwdBuffers_1_result;
    end else begin
      extnMRequest_rs1 <= prf_toExec_rs1Data;
    end
    if (_singleCycleArithmeticRequest_rs2_T_5) begin // @[Mux.scala 101:16]
      extnMRequest_rs2 <= fwdFrom_0_result;
    end else if (_singleCycleArithmeticRequest_rs2_T_7) begin // @[Mux.scala 101:16]
      extnMRequest_rs2 <= fwdBuffers_0_result;
    end else if (_singleCycleArithmeticRequest_rs2_T_9) begin // @[Mux.scala 101:16]
      extnMRequest_rs2 <= fwdBuffers_1_result;
    end else begin
      extnMRequest_rs2 <= prf_toExec_rs2Data;
    end
    extnMRequest_instruction <= prf_toExec_instruction; // @[core.scala 334:28]
    extnMRequest_prfDest <= prf_toExec_prfDest; // @[core.scala 343:24]
    extnMRequest_robAddr <= prf_toExec_robAddr[3:0]; // @[core.scala 344:24]
    if (branchEvals_valid) begin // @[core.scala 391:25]
      if (_T_10) begin // @[core.scala 394:73]
        extnMRequest_branchMask <= _addressGenerationInput_branchMask_T; // @[core.scala 395:11]
      end else begin
        extnMRequest_branchMask <= _GEN_24;
      end
    end else begin
      extnMRequest_branchMask <= _GEN_24;
    end
    if (reset) begin // @[core.scala 228:31]
      extnMServicing_valid <= 1'h0; // @[core.scala 228:31]
    end else if (branchEvals_valid) begin // @[core.scala 391:25]
      if (_T) begin // @[core.scala 397:29]
        if (_T_57 & extnMRequest_valid) begin // @[core.scala 400:101]
          extnMServicing_valid <= 1'h0; // @[core.scala 400:107]
        end else begin
          extnMServicing_valid <= extnMPartialServicing_valid; // @[core.scala 232:18]
        end
      end else begin
        extnMServicing_valid <= extnMPartialServicing_valid; // @[core.scala 232:18]
      end
    end else begin
      extnMServicing_valid <= extnMPartialServicing_valid; // @[core.scala 232:18]
    end
    extnMServicing_instruction <= extnMPartialServicing_instruction; // @[core.scala 232:18]
    extnMServicing_prfDest <= extnMPartialServicing_prfDest; // @[core.scala 232:18]
    extnMServicing_robAddr <= extnMPartialServicing_robAddr; // @[core.scala 232:18]
    if (branchEvals_valid) begin // @[core.scala 391:25]
      if (_T_60) begin // @[core.scala 394:73]
        extnMServicing_branchMask <= _T_58; // @[core.scala 395:11]
      end else begin
        extnMServicing_branchMask <= extnMPartialServicing_branchMask; // @[core.scala 232:18]
      end
    end else begin
      extnMServicing_branchMask <= extnMPartialServicing_branchMask; // @[core.scala 232:18]
    end
    if (reset) begin // @[core.scala 229:38]
      extnMPartialServicing_valid <= 1'h0; // @[core.scala 229:38]
    end else if (extnMRequest_instruction[14]) begin // @[core.scala 233:45]
      extnMPartialServicing_valid <= 1'h0; // @[core.scala 233:75]
    end else begin
      extnMPartialServicing_valid <= extnMRequest_valid; // @[core.scala 231:25]
    end
    extnMPartialServicing_instruction <= extnMRequest_instruction; // @[core.scala 231:25]
    extnMPartialServicing_prfDest <= extnMRequest_prfDest; // @[core.scala 231:25]
    extnMPartialServicing_robAddr <= extnMRequest_robAddr; // @[core.scala 231:25]
    if (branchEvals_valid) begin // @[core.scala 391:25]
      if (_T_57) begin // @[core.scala 394:73]
        extnMPartialServicing_branchMask <= _T_55; // @[core.scala 395:11]
      end else begin
        extnMPartialServicing_branchMask <= extnMRequest_branchMask; // @[core.scala 231:25]
      end
    end else begin
      extnMPartialServicing_branchMask <= extnMRequest_branchMask; // @[core.scala 231:25]
    end
    muls_0 <= _GEN_94 + _muls_0_T; // @[core.scala 367:29]
    muls_1 <= _GEN_108 + _muls_1_T; // @[core.scala 368:28]
    muls_2 <= _GEN_108 + _muls_2_T; // @[core.scala 369:28]
    muls_3 <= _muls_3_T_3 + _muls_3_T_4; // @[core.scala 370:62]
    muls_4 <= _GEN_94 + _muls_4_T; // @[core.scala 371:28]
    muls_5 <= {{32'd0}, narrowMuls_8}; // @[core.scala 372:11]
    extnMResponse_result <= _GEN_120[63:0];
    if (division_request_valid & ~(|division_counter)) begin // @[core.scala 450:57]
      extnMResponse_robAddr <= division_request_robAddr; // @[core.scala 470:27]
    end else begin
      extnMResponse_robAddr <= extnMServicing_robAddr; // @[core.scala 387:25]
    end
    if (reset) begin // @[core.scala 237:25]
      division_request_valid <= 1'h0; // @[core.scala 237:25]
    end else if (branchEvals_valid) begin // @[core.scala 479:25]
      if (_T & _T_107) begin // @[core.scala 485:89]
        division_request_valid <= 1'h0; // @[core.scala 485:114]
      end else if (extnMRequest_valid) begin // @[core.scala 480:30]
        division_request_valid <= _GEN_126;
      end else begin
        division_request_valid <= _GEN_124;
      end
    end else begin
      division_request_valid <= _GEN_124;
    end
    if (extnMRequest_valid & extnMRequest_instruction[14]) begin // @[core.scala 428:67]
      division_request_rs1 <= extnMRequest_rs1; // @[core.scala 437:22]
    end
    if (extnMRequest_valid & extnMRequest_instruction[14]) begin // @[core.scala 428:67]
      division_request_rs2 <= extnMRequest_rs2; // @[core.scala 437:22]
    end
    if (extnMRequest_valid & extnMRequest_instruction[14]) begin // @[core.scala 428:67]
      division_request_instruction <= extnMRequest_instruction; // @[core.scala 437:22]
    end
    if (extnMRequest_valid & extnMRequest_instruction[14]) begin // @[core.scala 428:67]
      division_request_prfDest <= extnMRequest_prfDest; // @[core.scala 437:22]
    end
    if (extnMRequest_valid & extnMRequest_instruction[14]) begin // @[core.scala 428:67]
      division_request_robAddr <= extnMRequest_robAddr; // @[core.scala 437:22]
    end
    if (branchEvals_valid) begin // @[core.scala 479:25]
      if (_T_107) begin // @[core.scala 484:69]
        division_request_branchMask <= _division_request_branchMask_T_1; // @[core.scala 484:99]
      end else if (extnMRequest_valid) begin // @[core.scala 480:30]
        if (_T_57) begin // @[core.scala 481:67]
          division_request_branchMask <= _T_55; // @[core.scala 481:97]
        end else begin
          division_request_branchMask <= _GEN_107;
        end
      end else begin
        division_request_branchMask <= _GEN_107;
      end
    end else begin
      division_request_branchMask <= _GEN_107;
    end
    if (extnMRequest_valid & extnMRequest_instruction[14]) begin // @[core.scala 428:67]
      if (~extnMRequest_instruction[12]) begin // @[core.scala 439:47]
        if (extnMRequest_instruction[3]) begin // @[core.scala 443:48]
          if (extnMRequest_rs1[31]) begin // @[core.scala 444:43]
            division_quotient <= _division_quotient_T_24; // @[core.scala 444:63]
          end else begin
            division_quotient <= _GEN_88;
          end
        end else begin
          division_quotient <= _GEN_88;
        end
      end else begin
        division_quotient <= _GEN_87;
      end
    end else begin
      division_quotient <= _division_quotient_T_13; // @[core.scala 425:21]
    end
    if (extnMRequest_valid & extnMRequest_instruction[14]) begin // @[core.scala 428:67]
      division_remainder <= 65'h0; // @[core.scala 436:24]
    end else begin
      division_remainder <= _division_remainder_T_9; // @[core.scala 424:22]
    end
    if (extnMRequest_valid & extnMRequest_instruction[14]) begin // @[core.scala 428:67]
      if (~extnMRequest_instruction[12]) begin // @[core.scala 439:47]
        if (extnMRequest_instruction[3]) begin // @[core.scala 443:48]
          if (extnMRequest_rs2[31]) begin // @[core.scala 445:43]
            division_divisor <= _division_divisor_T_10; // @[core.scala 445:62]
          end else begin
            division_divisor <= _GEN_89;
          end
        end else begin
          division_divisor <= _GEN_89;
        end
      end else begin
        division_divisor <= _GEN_86;
      end
    end
    if (extnMRequest_valid & extnMRequest_instruction[14]) begin // @[core.scala 428:67]
      division_counter <= 7'h41; // @[core.scala 429:22]
    end else begin
      division_counter <= _division_counter_T_1; // @[core.scala 426:20]
    end
    if (reset) begin // @[core.scala 246:27]
      fwdBuffers_0_valid <= 1'h0; // @[core.scala 246:27]
    end else begin
      fwdBuffers_0_valid <= fwdFrom_0_valid; // @[core.scala 490:64]
    end
    fwdBuffers_0_prfDest <= singleCycleArithmeticRequest_prfDest; // @[core.scala 252:33 256:22]
    fwdBuffers_0_result <= arithmeticResult[63:0]; // @[core.scala 252:33 293:21]
    if (reset) begin // @[core.scala 246:27]
      fwdBuffers_1_valid <= 1'h0; // @[core.scala 246:27]
    end else begin
      fwdBuffers_1_valid <= fwdBuffers_0_valid; // @[core.scala 490:64]
    end
    fwdBuffers_1_prfDest <= fwdBuffers_0_prfDest; // @[core.scala 252:33 253:14]
    fwdBuffers_1_result <= fwdBuffers_0_result; // @[core.scala 252:33 253:14]
    narrowMuls_0 <= extnMRequest_rs1[31:0] * extnMRequest_rs2[31:0]; // @[core.scala 353:29]
    narrowMuls_1 <= extnMRequest_rs1[63:32] * extnMRequest_rs2[31:0]; // @[core.scala 354:30]
    narrowMuls_2 <= _T_39[63:0]; // @[core.scala 364:80]
    narrowMuls_3 <= extnMRequest_rs1[31:0] * extnMRequest_rs2[63:32]; // @[core.scala 356:29]
    narrowMuls_4 <= _T_40[63:0]; // @[core.scala 364:80]
    narrowMuls_5 <= extnMRequest_rs1[63:32] * extnMRequest_rs2[63:32]; // @[core.scala 358:30]
    narrowMuls_6 <= _T_41[63:0]; // @[core.scala 364:80]
    narrowMuls_7 <= $signed(_partialMuls32x32_T_30) * $signed(_partialMuls32x32_T_32); // @[core.scala 364:41]
    narrowMuls_8 <= $signed(_partialMuls32x32_T_34) * $signed(_partialMuls32x32_T_36); // @[core.scala 364:41]
    if (~mExtensionReady) begin // @[core.scala 412:26]
      if (branchEvals_valid & |_T_78) begin // @[core.scala 413:73]
        if (branchEvals_passed) begin // @[core.scala 414:30]
          divBranchMask <= _divBranchMask_T_5; // @[core.scala 415:23]
        end else begin
          divBranchMask <= _GEN_78;
        end
      end else begin
        divBranchMask <= _GEN_78;
      end
    end else begin
      divBranchMask <= _GEN_78;
    end
    if (reset) begin // @[core.scala 500:26]
      branchPCs_0_valid <= 1'h0; // @[core.scala 500:26]
    end else if (branchEvals_valid & _T) begin // @[core.scala 641:46]
      branchPCs_0_valid <= 1'h0; // @[core.scala 642:32]
    end else if (branchInstruction_valid) begin // @[core.scala 643:39]
      branchPCs_0_valid <= entry_1_valid; // @[core.scala 654:40]
    end else if (~branchPCs_0_valid) begin // @[core.scala 636:82]
      branchPCs_0_valid <= decode_branchPCs_branchPCReady; // @[core.scala 637:15]
    end
    if (branchEvals_valid & _T) begin // @[core.scala 641:46]
      branchPCs_0_pc <= _GEN_161;
    end else if (branchInstruction_valid) begin // @[core.scala 643:39]
      if (branchPCs_1_valid) begin // @[core.scala 648:22]
        branchPCs_0_pc <= branchPCs_1_pc;
      end else begin
        branchPCs_0_pc <= decode_branchPCs_branchPC;
      end
    end else begin
      branchPCs_0_pc <= _GEN_161;
    end
    if (branchEvals_valid & _T) begin // @[core.scala 641:46]
      branchPCs_0_branchMask <= _GEN_162;
    end else if (branchInstruction_valid) begin // @[core.scala 643:39]
      if (branchPCs_1_valid) begin // @[core.scala 649:30]
        branchPCs_0_branchMask <= branchPCs_1_branchMask;
      end else begin
        branchPCs_0_branchMask <= decode_branchPCs_branchMask;
      end
    end else begin
      branchPCs_0_branchMask <= _GEN_162;
    end
    if (reset) begin // @[core.scala 500:26]
      branchPCs_1_valid <= 1'h0; // @[core.scala 500:26]
    end else if (branchEvals_valid & _T) begin // @[core.scala 641:46]
      branchPCs_1_valid <= 1'h0; // @[core.scala 642:32]
    end else if (branchInstruction_valid) begin // @[core.scala 643:39]
      branchPCs_1_valid <= entry_2_valid; // @[core.scala 654:40]
    end else if (branchPCs_0_valid & ~branchPCs_1_valid) begin // @[core.scala 636:82]
      branchPCs_1_valid <= decode_branchPCs_branchPCReady; // @[core.scala 637:15]
    end
    if (branchEvals_valid & _T) begin // @[core.scala 641:46]
      branchPCs_1_pc <= _GEN_164;
    end else if (branchInstruction_valid) begin // @[core.scala 643:39]
      if (branchPCs_2_valid) begin // @[core.scala 648:22]
        branchPCs_1_pc <= branchPCs_2_pc;
      end else begin
        branchPCs_1_pc <= decode_branchPCs_branchPC;
      end
    end else begin
      branchPCs_1_pc <= _GEN_164;
    end
    if (branchEvals_valid & _T) begin // @[core.scala 641:46]
      branchPCs_1_branchMask <= _GEN_165;
    end else if (branchInstruction_valid) begin // @[core.scala 643:39]
      if (branchPCs_2_valid) begin // @[core.scala 649:30]
        branchPCs_1_branchMask <= branchPCs_2_branchMask;
      end else begin
        branchPCs_1_branchMask <= decode_branchPCs_branchMask;
      end
    end else begin
      branchPCs_1_branchMask <= _GEN_165;
    end
    if (reset) begin // @[core.scala 500:26]
      branchPCs_2_valid <= 1'h0; // @[core.scala 500:26]
    end else if (branchEvals_valid & _T) begin // @[core.scala 641:46]
      branchPCs_2_valid <= 1'h0; // @[core.scala 642:32]
    end else if (branchInstruction_valid) begin // @[core.scala 643:39]
      branchPCs_2_valid <= entry_3_valid; // @[core.scala 654:40]
    end else if (_T_133 & ~branchPCs_2_valid) begin // @[core.scala 636:82]
      branchPCs_2_valid <= decode_branchPCs_branchPCReady; // @[core.scala 637:15]
    end
    if (branchEvals_valid & _T) begin // @[core.scala 641:46]
      branchPCs_2_pc <= _GEN_167;
    end else if (branchInstruction_valid) begin // @[core.scala 643:39]
      if (branchPCs_3_valid) begin // @[core.scala 648:22]
        branchPCs_2_pc <= branchPCs_3_pc;
      end else begin
        branchPCs_2_pc <= decode_branchPCs_branchPC;
      end
    end else begin
      branchPCs_2_pc <= _GEN_167;
    end
    if (branchEvals_valid & _T) begin // @[core.scala 641:46]
      branchPCs_2_branchMask <= _GEN_168;
    end else if (branchInstruction_valid) begin // @[core.scala 643:39]
      if (branchPCs_3_valid) begin // @[core.scala 649:30]
        branchPCs_2_branchMask <= branchPCs_3_branchMask;
      end else begin
        branchPCs_2_branchMask <= decode_branchPCs_branchMask;
      end
    end else begin
      branchPCs_2_branchMask <= _GEN_168;
    end
    if (reset) begin // @[core.scala 500:26]
      branchPCs_3_valid <= 1'h0; // @[core.scala 500:26]
    end else if (branchEvals_valid & _T) begin // @[core.scala 641:46]
      branchPCs_3_valid <= 1'h0; // @[core.scala 642:32]
    end else if (branchInstruction_valid) begin // @[core.scala 643:39]
      branchPCs_3_valid <= 1'h0; // @[core.scala 655:41]
    end else if (_T_134 & ~branchPCs_3_valid) begin // @[core.scala 636:82]
      branchPCs_3_valid <= decode_branchPCs_branchPCReady; // @[core.scala 637:15]
    end
    if (_T_134 & ~branchPCs_3_valid) begin // @[core.scala 636:82]
      branchPCs_3_pc <= decode_branchPCs_branchPC; // @[core.scala 638:12]
    end
    if (_T_134 & ~branchPCs_3_valid) begin // @[core.scala 636:82]
      branchPCs_3_branchMask <= decode_branchPCs_branchMask; // @[core.scala 639:20]
    end
    if (reset) begin // @[core.scala 507:29]
      predictedPCs_0_valid <= 1'h0; // @[core.scala 507:29]
    end else if (_T_145) begin // @[core.scala 664:46]
      predictedPCs_0_valid <= 1'h0; // @[core.scala 665:35]
    end else if (branchInstruction_valid) begin // @[core.scala 666:39]
      predictedPCs_0_valid <= entry_5_valid; // @[core.scala 676:40]
    end else if (~predictedPCs_0_valid) begin // @[core.scala 660:82]
      predictedPCs_0_valid <= decode_branchPCs_predictedPCReady; // @[core.scala 661:15]
    end
    if (_T_145) begin // @[core.scala 664:46]
      predictedPCs_0_pc <= _GEN_193;
    end else if (branchInstruction_valid) begin // @[core.scala 666:39]
      if (predictedPCs_1_valid) begin // @[core.scala 671:22]
        predictedPCs_0_pc <= predictedPCs_1_pc;
      end else begin
        predictedPCs_0_pc <= decode_branchPCs_predictedPC;
      end
    end else begin
      predictedPCs_0_pc <= _GEN_193;
    end
    if (reset) begin // @[core.scala 507:29]
      predictedPCs_1_valid <= 1'h0; // @[core.scala 507:29]
    end else if (_T_145) begin // @[core.scala 664:46]
      predictedPCs_1_valid <= 1'h0; // @[core.scala 665:35]
    end else if (branchInstruction_valid) begin // @[core.scala 666:39]
      predictedPCs_1_valid <= entry_6_valid; // @[core.scala 676:40]
    end else if (predictedPCs_0_valid & ~predictedPCs_1_valid) begin // @[core.scala 660:82]
      predictedPCs_1_valid <= decode_branchPCs_predictedPCReady; // @[core.scala 661:15]
    end
    if (_T_145) begin // @[core.scala 664:46]
      predictedPCs_1_pc <= _GEN_195;
    end else if (branchInstruction_valid) begin // @[core.scala 666:39]
      if (predictedPCs_2_valid) begin // @[core.scala 671:22]
        predictedPCs_1_pc <= predictedPCs_2_pc;
      end else begin
        predictedPCs_1_pc <= decode_branchPCs_predictedPC;
      end
    end else begin
      predictedPCs_1_pc <= _GEN_195;
    end
    if (reset) begin // @[core.scala 507:29]
      predictedPCs_2_valid <= 1'h0; // @[core.scala 507:29]
    end else if (_T_145) begin // @[core.scala 664:46]
      predictedPCs_2_valid <= 1'h0; // @[core.scala 665:35]
    end else if (branchInstruction_valid) begin // @[core.scala 666:39]
      predictedPCs_2_valid <= entry_7_valid; // @[core.scala 676:40]
    end else if (_T_151 & ~predictedPCs_2_valid) begin // @[core.scala 660:82]
      predictedPCs_2_valid <= decode_branchPCs_predictedPCReady; // @[core.scala 661:15]
    end
    if (_T_145) begin // @[core.scala 664:46]
      predictedPCs_2_pc <= _GEN_197;
    end else if (branchInstruction_valid) begin // @[core.scala 666:39]
      if (predictedPCs_3_valid) begin // @[core.scala 671:22]
        predictedPCs_2_pc <= predictedPCs_3_pc;
      end else begin
        predictedPCs_2_pc <= decode_branchPCs_predictedPC;
      end
    end else begin
      predictedPCs_2_pc <= _GEN_197;
    end
    if (reset) begin // @[core.scala 507:29]
      predictedPCs_3_valid <= 1'h0; // @[core.scala 507:29]
    end else if (_T_145) begin // @[core.scala 664:46]
      predictedPCs_3_valid <= 1'h0; // @[core.scala 665:35]
    end else if (branchInstruction_valid) begin // @[core.scala 666:39]
      predictedPCs_3_valid <= 1'h0; // @[core.scala 677:44]
    end else if (_T_152 & ~predictedPCs_3_valid) begin // @[core.scala 660:82]
      predictedPCs_3_valid <= decode_branchPCs_predictedPCReady; // @[core.scala 661:15]
    end
    if (_T_152 & ~predictedPCs_3_valid) begin // @[core.scala 660:82]
      predictedPCs_3_pc <= decode_branchPCs_predictedPC; // @[core.scala 662:12]
    end
    if (reset) begin // @[core.scala 512:34]
      branchInstruction_valid <= 1'h0; // @[core.scala 512:34]
    end else if (branchEvals_valid) begin // @[core.scala 558:25]
      if (_T & |_T_128) begin // @[core.scala 562:83]
        branchInstruction_valid <= 1'h0; // @[core.scala 563:31]
      end else begin
        branchInstruction_valid <= prf_toExec_valid & prf_toExec_instruction[6:4] == 3'h6; // @[core.scala 545:27]
      end
    end else begin
      branchInstruction_valid <= prf_toExec_valid & prf_toExec_instruction[6:4] == 3'h6; // @[core.scala 545:27]
    end
    if (prf_toExec_valid & prf_toExec_instruction[6:5] == 2'h3) begin // @[core.scala 546:71]
      if (_addressGenerationInput_rs1_T_3) begin // @[Mux.scala 101:16]
        branchInstruction_rs1 <= fwdFrom_0_result;
      end else if (_addressGenerationInput_rs1_T_5) begin // @[Mux.scala 101:16]
        branchInstruction_rs1 <= fwdBuffers_0_result;
      end else if (_addressGenerationInput_rs1_T_7) begin // @[Mux.scala 101:16]
        branchInstruction_rs1 <= fwdBuffers_1_result;
      end else begin
        branchInstruction_rs1 <= prf_toExec_rs1Data;
      end
    end
    if (prf_toExec_valid & prf_toExec_instruction[6:5] == 2'h3) begin // @[core.scala 546:71]
      if (_singleCycleArithmeticRequest_rs2_T_5) begin // @[Mux.scala 101:16]
        branchInstruction_rs2 <= fwdFrom_0_result;
      end else if (_singleCycleArithmeticRequest_rs2_T_7) begin // @[Mux.scala 101:16]
        branchInstruction_rs2 <= fwdBuffers_0_result;
      end else if (_singleCycleArithmeticRequest_rs2_T_9) begin // @[Mux.scala 101:16]
        branchInstruction_rs2 <= fwdBuffers_1_result;
      end else begin
        branchInstruction_rs2 <= prf_toExec_rs2Data;
      end
    end
    branchInstruction_robAddr <= _GEN_140[3:0];
    if (prf_toExec_valid & prf_toExec_instruction[6:5] == 2'h3) begin // @[core.scala 546:71]
      branchInstruction_instruction <= prf_toExec_instruction; // @[core.scala 555:35]
    end
    if (2'h3 == prf_toExec_instruction[3:2]) begin // @[core.scala 523:31]
      branchInstruction_immediate <= _branchInstruction_immediate_T_18; // @[core.scala 523:31]
    end else if (2'h2 == prf_toExec_instruction[3:2]) begin // @[core.scala 523:31]
      branchInstruction_immediate <= 64'h0; // @[core.scala 523:31]
    end else if (2'h1 == prf_toExec_instruction[3:2]) begin // @[core.scala 523:31]
      branchInstruction_immediate <= arithmeticImm; // @[core.scala 523:31]
    end else begin
      branchInstruction_immediate <= _branchInstruction_immediate_T_6;
    end
    if (coherentLoadInvalid) begin // @[core.scala 572:29]
      branchEvals_robAddr <= _branchEvals_robAddr_T_1;
    end else begin
      branchEvals_robAddr <= branchInstruction_robAddr;
    end
    if (coherentLoadInvalid) begin // @[core.scala 627:28]
      branchEvals_nextPC <= rob_commit_pc;
    end else if (2'h3 == branchInstruction_instruction[3:2]) begin // @[core.scala 627:28]
      branchEvals_nextPC <= _nextCorrectPC_T_2; // @[core.scala 627:28]
    end else if (2'h2 == branchInstruction_instruction[3:2]) begin // @[core.scala 627:28]
      branchEvals_nextPC <= 64'h0; // @[core.scala 627:28]
    end else if (2'h1 == branchInstruction_instruction[3:2]) begin // @[core.scala 627:28]
      branchEvals_nextPC <= _nextCorrectPC_T_7; // @[core.scala 627:28]
    end else begin
      branchEvals_nextPC <= _nextCorrectPC_T_5;
    end
    coherentLoadInvalidReg <= ~memAccess_loadCommit_state & memAccess_loadCommit_valid & rob_commit_ready & ~(|
      rob_commit_instruction[6:2]); // @[core.scala 568:107]
    rob_execPorts_0_mtval_REG <= singleCycleArithmeticRequest_rs1; // @[core.scala 758:36]
    if (reset) begin // @[core.scala 779:129]
      REG <= 1'h0; // @[core.scala 779:129]
    end else begin
      REG <= _fwdFrom_0_valid_T_1 & singleCycleArithmeticRequest_instruction[6:2] != 5'h1c; // @[core.scala 779:129]
    end
    prf_fromStore_rs2Addr_REG <= dataQueue_toPRF_rs2Addr; // @[core.scala 815:43]
    prf_fromStore_rs2Addr_REG_1 <= prf_fromStore_rs2Addr_REG; // @[core.scala 815:35]
    if (reset) begin // @[core.scala 816:41]
      prf_fromStore_valid_REG <= 1'h0; // @[core.scala 816:41]
    end else begin
      prf_fromStore_valid_REG <= dataQueue_toPRF_valid & dataQueue_fromROB_readyNow; // @[core.scala 816:41]
    end
    if (reset) begin // @[core.scala 816:33]
      prf_fromStore_valid_REG_1 <= 1'h0; // @[core.scala 816:33]
    end else begin
      prf_fromStore_valid_REG_1 <= prf_fromStore_valid_REG; // @[core.scala 816:33]
    end
    if (reset) begin // @[core.scala 862:27]
      fenceState_state <= 2'h0; // @[core.scala 862:27]
    end else if (2'h0 == fenceState_state) begin // @[core.scala 869:28]
      if (fetch_toDecode_fired & _T_188 == 20'hf) begin // @[core.scala 871:115]
        fenceState_state <= 2'h1; // @[core.scala 872:26]
      end
    end else if (2'h1 == fenceState_state) begin // @[core.scala 869:28]
      if (_T_145) begin // @[core.scala 876:54]
        fenceState_state <= 2'h0; // @[core.scala 879:26]
      end else begin
        fenceState_state <= _GEN_223;
      end
    end else if (2'h2 == fenceState_state) begin // @[core.scala 869:28]
      fenceState_state <= _GEN_233;
    end
    if (!(2'h0 == fenceState_state)) begin // @[core.scala 869:28]
      if (2'h1 == fenceState_state) begin // @[core.scala 869:28]
        if (!(_T_145)) begin // @[core.scala 876:54]
          if (decode_toExec_fired & _T_195 == 20'hf) begin // @[core.scala 880:119]
            fenceState_branchMask <= decode_toExec_branchMask; // @[core.scala 882:31]
          end
        end
      end else if (2'h2 == fenceState_state) begin // @[core.scala 869:28]
        if (!(branchEvals_valid & |_T_199 & _T)) begin // @[core.scala 886:110]
          fenceState_branchMask <= _GEN_231;
        end
      end
    end
    REG_1 <= _T_145 & (fetch_toDecode_instruction == 32'hff0000f & fetch_toDecode_fired); // @[core.scala 920:53]
    branchCounter <= _GEN_249[2:0]; // @[core.scala 1033:{30,30}]
    if (branchEvals_valid) begin // @[core.scala 1049:27]
      lastBranchExecRob <= branchEvals_robAddr; // @[core.scala 1050:23]
    end
    if (branchEvals_valid) begin // @[core.scala 1049:27]
      lastBranchExecPC <= lastBranchExecPC_REG; // @[core.scala 1051:22]
    end
    lastBranchExecPC_REG <= branchPCs_0_pc; // @[core.scala 1051:32]
    if (reset) begin // @[core.scala 1067:34]
      lastRetiredSystem <= 1'h0; // @[core.scala 1067:34]
    end else if (decode_fromFetch_fired) begin // @[core.scala 1068:32]
      lastRetiredSystem <= fetch_toDecode_instruction[6:0] == 7'h73; // @[core.scala 1068:52]
    end
    if (reset) begin // @[core.scala 1070:38]
      interruptInjectStatus <= 2'h0; // @[core.scala 1070:38]
    end else if (2'h0 == interruptInjectStatus) begin // @[core.scala 1071:33]
      if (decode_canTakeInterrupt & MTIP & ~lastRetiredSystem) begin // @[core.scala 1075:67]
        interruptInjectStatus <= 2'h1; // @[core.scala 1075:91]
      end
    end else if (2'h1 == interruptInjectStatus) begin // @[core.scala 1071:33]
      if (decode_canTakeInterrupt) begin // @[core.scala 1079:56]
        interruptInjectStatus <= _GEN_280;
      end
    end else if (2'h2 == interruptInjectStatus) begin // @[core.scala 1071:33]
      interruptInjectStatus <= 2'h3; // @[core.scala 1103:29]
    end else begin
      interruptInjectStatus <= _GEN_290;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  branchEvals_branchMask = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  branchEvals_passed = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  branchEvals_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  extnMResponse_prfDest = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  extnMResponse_valid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  extnResponseInstruction = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  mExtensionReady = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  addressGenerationInput_valid = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  addressGenerationInput_rs1 = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  addressGenerationInput_instruction = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  addressGenerationInput_prfDest = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  addressGenerationInput_robAddr = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  addressGenerationInput_branchMask = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  memoryRequest_valid = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  memoryRequest_address = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  memoryRequest_instruction = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  memoryRequest_branchMask = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  memoryRequest_robAddr = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  memoryRequest_prfDest = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  singleCycleArithmeticRequest_valid = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  singleCycleArithmeticRequest_rs1 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  singleCycleArithmeticRequest_rs2 = _RAND_21[63:0];
  _RAND_22 = {1{`RANDOM}};
  singleCycleArithmeticRequest_instruction = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  singleCycleArithmeticRequest_prfDest = _RAND_23[5:0];
  _RAND_24 = {1{`RANDOM}};
  singleCycleArithmeticRequest_robAddr = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  singleCycleArithmeticRequest_branchMask = _RAND_25[4:0];
  _RAND_26 = {1{`RANDOM}};
  singleCycleArithmeticResponse_valid = _RAND_26[0:0];
  _RAND_27 = {2{`RANDOM}};
  singleCycleArithmeticResponse_result = _RAND_27[63:0];
  _RAND_28 = {1{`RANDOM}};
  singleCycleArithmeticResponse_prfDest = _RAND_28[5:0];
  _RAND_29 = {1{`RANDOM}};
  singleCycleArithmeticResponse_robAddr = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  extnMRequest_valid = _RAND_30[0:0];
  _RAND_31 = {2{`RANDOM}};
  extnMRequest_rs1 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  extnMRequest_rs2 = _RAND_32[63:0];
  _RAND_33 = {1{`RANDOM}};
  extnMRequest_instruction = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  extnMRequest_prfDest = _RAND_34[5:0];
  _RAND_35 = {1{`RANDOM}};
  extnMRequest_robAddr = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  extnMRequest_branchMask = _RAND_36[4:0];
  _RAND_37 = {1{`RANDOM}};
  extnMServicing_valid = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  extnMServicing_instruction = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  extnMServicing_prfDest = _RAND_39[5:0];
  _RAND_40 = {1{`RANDOM}};
  extnMServicing_robAddr = _RAND_40[3:0];
  _RAND_41 = {1{`RANDOM}};
  extnMServicing_branchMask = _RAND_41[4:0];
  _RAND_42 = {1{`RANDOM}};
  extnMPartialServicing_valid = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  extnMPartialServicing_instruction = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  extnMPartialServicing_prfDest = _RAND_44[5:0];
  _RAND_45 = {1{`RANDOM}};
  extnMPartialServicing_robAddr = _RAND_45[3:0];
  _RAND_46 = {1{`RANDOM}};
  extnMPartialServicing_branchMask = _RAND_46[4:0];
  _RAND_47 = {3{`RANDOM}};
  muls_0 = _RAND_47[95:0];
  _RAND_48 = {3{`RANDOM}};
  muls_1 = _RAND_48[95:0];
  _RAND_49 = {3{`RANDOM}};
  muls_2 = _RAND_49[95:0];
  _RAND_50 = {3{`RANDOM}};
  muls_3 = _RAND_50[95:0];
  _RAND_51 = {3{`RANDOM}};
  muls_4 = _RAND_51[95:0];
  _RAND_52 = {3{`RANDOM}};
  muls_5 = _RAND_52[95:0];
  _RAND_53 = {2{`RANDOM}};
  extnMResponse_result = _RAND_53[63:0];
  _RAND_54 = {1{`RANDOM}};
  extnMResponse_robAddr = _RAND_54[3:0];
  _RAND_55 = {1{`RANDOM}};
  division_request_valid = _RAND_55[0:0];
  _RAND_56 = {2{`RANDOM}};
  division_request_rs1 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  division_request_rs2 = _RAND_57[63:0];
  _RAND_58 = {1{`RANDOM}};
  division_request_instruction = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  division_request_prfDest = _RAND_59[5:0];
  _RAND_60 = {1{`RANDOM}};
  division_request_robAddr = _RAND_60[3:0];
  _RAND_61 = {1{`RANDOM}};
  division_request_branchMask = _RAND_61[4:0];
  _RAND_62 = {3{`RANDOM}};
  division_quotient = _RAND_62[64:0];
  _RAND_63 = {3{`RANDOM}};
  division_remainder = _RAND_63[64:0];
  _RAND_64 = {3{`RANDOM}};
  division_divisor = _RAND_64[64:0];
  _RAND_65 = {1{`RANDOM}};
  division_counter = _RAND_65[6:0];
  _RAND_66 = {1{`RANDOM}};
  fwdBuffers_0_valid = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  fwdBuffers_0_prfDest = _RAND_67[5:0];
  _RAND_68 = {2{`RANDOM}};
  fwdBuffers_0_result = _RAND_68[63:0];
  _RAND_69 = {1{`RANDOM}};
  fwdBuffers_1_valid = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  fwdBuffers_1_prfDest = _RAND_70[5:0];
  _RAND_71 = {2{`RANDOM}};
  fwdBuffers_1_result = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  narrowMuls_0 = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  narrowMuls_1 = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  narrowMuls_2 = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  narrowMuls_3 = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  narrowMuls_4 = _RAND_76[63:0];
  _RAND_77 = {2{`RANDOM}};
  narrowMuls_5 = _RAND_77[63:0];
  _RAND_78 = {2{`RANDOM}};
  narrowMuls_6 = _RAND_78[63:0];
  _RAND_79 = {2{`RANDOM}};
  narrowMuls_7 = _RAND_79[63:0];
  _RAND_80 = {2{`RANDOM}};
  narrowMuls_8 = _RAND_80[63:0];
  _RAND_81 = {1{`RANDOM}};
  divBranchMask = _RAND_81[4:0];
  _RAND_82 = {1{`RANDOM}};
  branchPCs_0_valid = _RAND_82[0:0];
  _RAND_83 = {2{`RANDOM}};
  branchPCs_0_pc = _RAND_83[63:0];
  _RAND_84 = {1{`RANDOM}};
  branchPCs_0_branchMask = _RAND_84[4:0];
  _RAND_85 = {1{`RANDOM}};
  branchPCs_1_valid = _RAND_85[0:0];
  _RAND_86 = {2{`RANDOM}};
  branchPCs_1_pc = _RAND_86[63:0];
  _RAND_87 = {1{`RANDOM}};
  branchPCs_1_branchMask = _RAND_87[4:0];
  _RAND_88 = {1{`RANDOM}};
  branchPCs_2_valid = _RAND_88[0:0];
  _RAND_89 = {2{`RANDOM}};
  branchPCs_2_pc = _RAND_89[63:0];
  _RAND_90 = {1{`RANDOM}};
  branchPCs_2_branchMask = _RAND_90[4:0];
  _RAND_91 = {1{`RANDOM}};
  branchPCs_3_valid = _RAND_91[0:0];
  _RAND_92 = {2{`RANDOM}};
  branchPCs_3_pc = _RAND_92[63:0];
  _RAND_93 = {1{`RANDOM}};
  branchPCs_3_branchMask = _RAND_93[4:0];
  _RAND_94 = {1{`RANDOM}};
  predictedPCs_0_valid = _RAND_94[0:0];
  _RAND_95 = {2{`RANDOM}};
  predictedPCs_0_pc = _RAND_95[63:0];
  _RAND_96 = {1{`RANDOM}};
  predictedPCs_1_valid = _RAND_96[0:0];
  _RAND_97 = {2{`RANDOM}};
  predictedPCs_1_pc = _RAND_97[63:0];
  _RAND_98 = {1{`RANDOM}};
  predictedPCs_2_valid = _RAND_98[0:0];
  _RAND_99 = {2{`RANDOM}};
  predictedPCs_2_pc = _RAND_99[63:0];
  _RAND_100 = {1{`RANDOM}};
  predictedPCs_3_valid = _RAND_100[0:0];
  _RAND_101 = {2{`RANDOM}};
  predictedPCs_3_pc = _RAND_101[63:0];
  _RAND_102 = {1{`RANDOM}};
  branchInstruction_valid = _RAND_102[0:0];
  _RAND_103 = {2{`RANDOM}};
  branchInstruction_rs1 = _RAND_103[63:0];
  _RAND_104 = {2{`RANDOM}};
  branchInstruction_rs2 = _RAND_104[63:0];
  _RAND_105 = {1{`RANDOM}};
  branchInstruction_robAddr = _RAND_105[3:0];
  _RAND_106 = {1{`RANDOM}};
  branchInstruction_instruction = _RAND_106[31:0];
  _RAND_107 = {2{`RANDOM}};
  branchInstruction_immediate = _RAND_107[63:0];
  _RAND_108 = {1{`RANDOM}};
  branchEvals_robAddr = _RAND_108[3:0];
  _RAND_109 = {2{`RANDOM}};
  branchEvals_nextPC = _RAND_109[63:0];
  _RAND_110 = {1{`RANDOM}};
  coherentLoadInvalidReg = _RAND_110[0:0];
  _RAND_111 = {2{`RANDOM}};
  rob_execPorts_0_mtval_REG = _RAND_111[63:0];
  _RAND_112 = {1{`RANDOM}};
  REG = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  prf_fromStore_rs2Addr_REG = _RAND_113[5:0];
  _RAND_114 = {1{`RANDOM}};
  prf_fromStore_rs2Addr_REG_1 = _RAND_114[5:0];
  _RAND_115 = {1{`RANDOM}};
  prf_fromStore_valid_REG = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  prf_fromStore_valid_REG_1 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  fenceState_state = _RAND_117[1:0];
  _RAND_118 = {1{`RANDOM}};
  fenceState_branchMask = _RAND_118[4:0];
  _RAND_119 = {1{`RANDOM}};
  REG_1 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  branchCounter = _RAND_120[2:0];
  _RAND_121 = {1{`RANDOM}};
  lastBranchExecRob = _RAND_121[3:0];
  _RAND_122 = {2{`RANDOM}};
  lastBranchExecPC = _RAND_122[63:0];
  _RAND_123 = {2{`RANDOM}};
  lastBranchExecPC_REG = _RAND_123[63:0];
  _RAND_124 = {1{`RANDOM}};
  lastRetiredSystem = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  interruptInjectStatus = _RAND_125[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module arbiter_1(
  input        clock,
  input        reset,
  input        io_AWVALID_0,
  output       io_AWREADY_0,
  input        io_WVALID_0,
  input        io_WLAST_0,
  output       io_WREADY_0,
  input        io_ARVALID_0,
  output       io_ARREADY_0,
  input        io_ARVALID_1,
  output       io_ARREADY_1,
  output [2:0] io_select,
  output       io_enq_valid,
  input        io_enq_ready,
  input        io_nstall
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] stateReg; // @[arbitter.scala 66:31]
  reg  wlast; // @[arbitter.scala 71:28]
  wire [3:0] _GEN_0 = io_AWVALID_0 ? 4'h4 : stateReg; // @[arbitter.scala 66:31 79:37 80:42]
  wire [1:0] _GEN_3 = io_enq_ready ? 2'h2 : 2'h1; // @[arbitter.scala 85:31 86:26 88:42]
  wire [3:0] _GEN_4 = io_nstall ? 4'h8 : 4'h2; // @[arbitter.scala 96:28 97:26 99:26]
  wire [2:0] _GEN_5 = io_enq_ready ? 3'h5 : 3'h4; // @[arbitter.scala 103:31 104:26 106:42]
  wire [2:0] _GEN_8 = io_enq_ready & io_WVALID_0 ? 3'h7 : 3'h6; // @[arbitter.scala 127:46 128:26 130:42]
  wire [3:0] _GEN_9 = io_nstall ? 4'h8 : 4'h7; // @[arbitter.scala 139:48 140:30 142:30]
  wire [3:0] _GEN_10 = ~wlast ? 4'h6 : _GEN_9; // @[arbitter.scala 136:25 137:26]
  wire [3:0] _GEN_12 = io_ARVALID_1 ? 4'h9 : stateReg; // @[arbitter.scala 153:37 154:42]
  wire [3:0] _GEN_13 = ~io_ARVALID_1 ? 4'h0 : _GEN_12; // @[arbitter.scala 151:48 152:26]
  wire [3:0] _GEN_14 = io_enq_ready ? 4'ha : 4'h9; // @[arbitter.scala 161:31 162:26 164:42]
  wire [3:0] _GEN_15 = io_nstall ? 4'h0 : 4'ha; // @[arbitter.scala 172:28 173:26 175:26]
  wire [3:0] _GEN_16 = io_enq_ready ? 4'hd : 4'hc; // @[arbitter.scala 179:31 180:26 182:42]
  wire [3:0] _GEN_19 = 4'hf == stateReg ? 4'he : stateReg; // @[arbitter.scala 73:21 66:31]
  wire [2:0] _GEN_22 = 4'hf == stateReg ? 3'h6 : 3'h0; // @[arbitter.scala 73:21 208:35 64:19]
  wire [3:0] _GEN_23 = 4'he == stateReg ? 4'he : _GEN_19; // @[arbitter.scala 73:21]
  wire [2:0] _GEN_26 = 4'he == stateReg ? 3'h0 : _GEN_22; // @[arbitter.scala 64:19 73:21]
  wire [3:0] _GEN_27 = 4'hd == stateReg ? 4'he : _GEN_23; // @[arbitter.scala 73:21 187:22]
  wire [2:0] _GEN_30 = 4'hd == stateReg ? 3'h5 : _GEN_26; // @[arbitter.scala 73:21 190:23]
  wire [3:0] _GEN_32 = 4'hc == stateReg ? _GEN_16 : _GEN_27; // @[arbitter.scala 73:21]
  wire [2:0] _GEN_35 = 4'hc == stateReg ? 3'h0 : _GEN_30; // @[arbitter.scala 64:19 73:21]
  wire  _GEN_37 = 4'ha == stateReg & io_ARVALID_1; // @[arbitter.scala 73:21 169:26 61:22]
  wire [2:0] _GEN_39 = 4'ha == stateReg ? 3'h4 : _GEN_35; // @[arbitter.scala 73:21 171:23]
  wire [3:0] _GEN_40 = 4'ha == stateReg ? _GEN_15 : _GEN_32; // @[arbitter.scala 73:21]
  wire [3:0] _GEN_43 = 4'h9 == stateReg ? _GEN_14 : _GEN_40; // @[arbitter.scala 73:21]
  wire  _GEN_44 = 4'h9 == stateReg ? 1'h0 : _GEN_37; // @[arbitter.scala 73:21 166:26]
  wire [2:0] _GEN_46 = 4'h9 == stateReg ? 3'h0 : _GEN_39; // @[arbitter.scala 64:19 73:21]
  wire [3:0] _GEN_49 = 4'h8 == stateReg ? _GEN_13 : _GEN_43; // @[arbitter.scala 73:21]
  wire  _GEN_50 = 4'h8 == stateReg ? 1'h0 : _GEN_44; // @[arbitter.scala 73:21 158:26]
  wire [2:0] _GEN_52 = 4'h8 == stateReg ? 3'h0 : _GEN_46; // @[arbitter.scala 64:19 73:21]
  wire [3:0] _GEN_55 = 4'h7 == stateReg ? _GEN_10 : _GEN_49; // @[arbitter.scala 73:21]
  wire  _GEN_56 = 4'h7 == stateReg & io_WVALID_0; // @[arbitter.scala 73:21 145:37 56:21]
  wire  _GEN_57 = 4'h7 == stateReg ? io_WVALID_0 : _GEN_50; // @[arbitter.scala 73:21 146:38]
  wire [2:0] _GEN_58 = 4'h7 == stateReg ? 3'h2 : _GEN_52; // @[arbitter.scala 73:21 147:35]
  wire  _GEN_59 = 4'h7 == stateReg ? 1'h0 : _GEN_50; // @[arbitter.scala 73:21 61:22]
  wire [3:0] _GEN_62 = 4'h6 == stateReg ? {{1'd0}, _GEN_8} : _GEN_55; // @[arbitter.scala 73:21]
  wire  _GEN_63 = 4'h6 == stateReg ? 1'h0 : _GEN_57; // @[arbitter.scala 73:21 132:26]
  wire  _GEN_64 = 4'h6 == stateReg ? io_WLAST_0 : wlast; // @[arbitter.scala 133:19 73:21 71:28]
  wire  _GEN_65 = 4'h6 == stateReg ? 1'h0 : _GEN_56; // @[arbitter.scala 56:21 73:21]
  wire [2:0] _GEN_66 = 4'h6 == stateReg ? 3'h0 : _GEN_58; // @[arbitter.scala 64:19 73:21]
  wire  _GEN_67 = 4'h6 == stateReg ? 1'h0 : _GEN_59; // @[arbitter.scala 73:21 61:22]
  wire [3:0] _GEN_70 = 4'h5 == stateReg ? 4'h6 : _GEN_62; // @[arbitter.scala 73:21]
  wire  _GEN_71 = 4'h5 == stateReg & io_AWVALID_0; // @[arbitter.scala 73:21 122:26 55:22]
  wire  _GEN_72 = 4'h5 == stateReg ? io_AWVALID_0 : _GEN_63; // @[arbitter.scala 73:21 123:26]
  wire [2:0] _GEN_73 = 4'h5 == stateReg ? 3'h1 : _GEN_66; // @[arbitter.scala 73:21 124:23]
  wire  _GEN_74 = 4'h5 == stateReg ? wlast : _GEN_64; // @[arbitter.scala 73:21 71:28]
  wire  _GEN_75 = 4'h5 == stateReg ? 1'h0 : _GEN_65; // @[arbitter.scala 56:21 73:21]
  wire  _GEN_76 = 4'h5 == stateReg ? 1'h0 : _GEN_67; // @[arbitter.scala 73:21 61:22]
  wire [3:0] _GEN_79 = 4'h4 == stateReg ? {{1'd0}, _GEN_5} : _GEN_70; // @[arbitter.scala 73:21]
  wire  _GEN_80 = 4'h4 == stateReg ? 1'h0 : _GEN_72; // @[arbitter.scala 73:21 108:26]
  wire  _GEN_82 = 4'h4 == stateReg ? 1'h0 : _GEN_71; // @[arbitter.scala 73:21 55:22]
  wire [2:0] _GEN_83 = 4'h4 == stateReg ? 3'h0 : _GEN_73; // @[arbitter.scala 64:19 73:21]
  wire  _GEN_84 = 4'h4 == stateReg ? wlast : _GEN_74; // @[arbitter.scala 73:21 71:28]
  wire  _GEN_85 = 4'h4 == stateReg ? 1'h0 : _GEN_75; // @[arbitter.scala 56:21 73:21]
  wire  _GEN_86 = 4'h4 == stateReg ? 1'h0 : _GEN_76; // @[arbitter.scala 73:21 61:22]
  wire  _GEN_89 = 4'h2 == stateReg & io_ARVALID_0; // @[arbitter.scala 73:21 57:22 93:26]
  wire  _GEN_90 = 4'h2 == stateReg ? io_ARVALID_0 : _GEN_80; // @[arbitter.scala 73:21 94:26]
  wire [2:0] _GEN_91 = 4'h2 == stateReg ? 3'h0 : _GEN_83; // @[arbitter.scala 73:21 95:23]
  wire  _GEN_94 = 4'h2 == stateReg ? 1'h0 : _GEN_82; // @[arbitter.scala 73:21 55:22]
  wire  _GEN_96 = 4'h2 == stateReg ? 1'h0 : _GEN_85; // @[arbitter.scala 56:21 73:21]
  wire  _GEN_97 = 4'h2 == stateReg ? 1'h0 : _GEN_86; // @[arbitter.scala 73:21 61:22]
  wire  _GEN_101 = 4'h1 == stateReg ? 1'h0 : _GEN_90; // @[arbitter.scala 73:21 90:26]
  wire  _GEN_102 = 4'h1 == stateReg ? 1'h0 : _GEN_89; // @[arbitter.scala 73:21 57:22]
  wire [2:0] _GEN_103 = 4'h1 == stateReg ? 3'h0 : _GEN_91; // @[arbitter.scala 64:19 73:21]
  wire  _GEN_105 = 4'h1 == stateReg ? 1'h0 : _GEN_94; // @[arbitter.scala 73:21 55:22]
  wire  _GEN_107 = 4'h1 == stateReg ? 1'h0 : _GEN_96; // @[arbitter.scala 56:21 73:21]
  wire  _GEN_108 = 4'h1 == stateReg ? 1'h0 : _GEN_97; // @[arbitter.scala 73:21 61:22]
  assign io_AWREADY_0 = 4'h0 == stateReg ? 1'h0 : _GEN_105; // @[arbitter.scala 73:21 55:22]
  assign io_WREADY_0 = 4'h0 == stateReg ? 1'h0 : _GEN_107; // @[arbitter.scala 56:21 73:21]
  assign io_ARREADY_0 = 4'h0 == stateReg ? 1'h0 : _GEN_102; // @[arbitter.scala 73:21 57:22]
  assign io_ARREADY_1 = 4'h0 == stateReg ? 1'h0 : _GEN_108; // @[arbitter.scala 73:21 61:22]
  assign io_select = 4'h0 == stateReg ? 3'h0 : _GEN_103; // @[arbitter.scala 64:19 73:21]
  assign io_enq_valid = 4'h0 == stateReg ? 1'h0 : _GEN_101; // @[arbitter.scala 73:21 82:26]
  always @(posedge clock) begin
    if (reset) begin // @[arbitter.scala 66:31]
      stateReg <= 4'h0; // @[arbitter.scala 66:31]
    end else if (4'h0 == stateReg) begin // @[arbitter.scala 73:21]
      if (~io_AWVALID_0 & ~io_ARVALID_0) begin // @[arbitter.scala 75:48]
        stateReg <= 4'h8; // @[arbitter.scala 76:26]
      end else if (io_ARVALID_0) begin // @[arbitter.scala 77:37]
        stateReg <= 4'h1; // @[arbitter.scala 78:42]
      end else begin
        stateReg <= _GEN_0;
      end
    end else if (4'h1 == stateReg) begin // @[arbitter.scala 73:21]
      stateReg <= {{2'd0}, _GEN_3};
    end else if (4'h2 == stateReg) begin // @[arbitter.scala 73:21]
      stateReg <= _GEN_4;
    end else begin
      stateReg <= _GEN_79;
    end
    if (reset) begin // @[arbitter.scala 71:28]
      wlast <= 1'h0; // @[arbitter.scala 71:28]
    end else if (!(4'h0 == stateReg)) begin // @[arbitter.scala 73:21]
      if (!(4'h1 == stateReg)) begin // @[arbitter.scala 73:21]
        if (!(4'h2 == stateReg)) begin // @[arbitter.scala 73:21]
          wlast <= _GEN_84;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  wlast = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ringbuffer(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [69:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [69:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [95:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [69:0] memReg [0:31]; // @[ringbuffer.scala 19:20]
  wire  memReg_io_deq_bits_MPORT_en; // @[ringbuffer.scala 19:20]
  wire [4:0] memReg_io_deq_bits_MPORT_addr; // @[ringbuffer.scala 19:20]
  wire [69:0] memReg_io_deq_bits_MPORT_data; // @[ringbuffer.scala 19:20]
  wire [69:0] memReg_MPORT_data; // @[ringbuffer.scala 19:20]
  wire [4:0] memReg_MPORT_addr; // @[ringbuffer.scala 19:20]
  wire  memReg_MPORT_mask; // @[ringbuffer.scala 19:20]
  wire  memReg_MPORT_en; // @[ringbuffer.scala 19:20]
  wire [69:0] memReg_MPORT_1_data; // @[ringbuffer.scala 19:20]
  wire [4:0] memReg_MPORT_1_addr; // @[ringbuffer.scala 19:20]
  wire  memReg_MPORT_1_mask; // @[ringbuffer.scala 19:20]
  wire  memReg_MPORT_1_en; // @[ringbuffer.scala 19:20]
  reg [4:0] readPtr; // @[ringbuffer.scala 14:24]
  reg [4:0] writePtr; // @[ringbuffer.scala 15:25]
  wire [4:0] _nextRead_T_2 = readPtr + 5'h1; // @[ringbuffer.scala 16:55]
  wire [4:0] nextRead = readPtr == 5'h1f ? 5'h0 : _nextRead_T_2; // @[ringbuffer.scala 16:21]
  wire [4:0] _nextWrite_T_2 = writePtr + 5'h1; // @[ringbuffer.scala 17:58]
  wire [4:0] nextWrite = writePtr == 5'h1f ? 5'h0 : _nextWrite_T_2; // @[ringbuffer.scala 17:22]
  reg  fullReg; // @[ringbuffer.scala 22:24]
  reg  emptyReg; // @[ringbuffer.scala 23:25]
  wire  _T = io_enq_valid & io_enq_ready; // @[ringbuffer.scala 39:23]
  wire  _T_1 = io_enq_valid & io_enq_ready & io_deq_valid; // @[ringbuffer.scala 39:39]
  wire  _T_2 = io_enq_valid & io_enq_ready & io_deq_valid & io_deq_ready; // @[ringbuffer.scala 39:55]
  wire  _T_4 = io_deq_valid & io_deq_ready; // @[ringbuffer.scala 48:29]
  wire  _GEN_12 = _T ? 1'h0 : _T_4; // @[ringbuffer.scala 43:45]
  wire  incrRead = io_enq_valid & io_enq_ready & io_deq_valid & io_deq_ready | _GEN_12; // @[ringbuffer.scala 39:70 40:15]
  wire  incrWrite = io_enq_valid & io_enq_ready & io_deq_valid & io_deq_ready | io_enq_valid & io_enq_ready; // @[ringbuffer.scala 39:70 41:16]
  wire  _GEN_4 = io_deq_valid & io_deq_ready ? nextRead == writePtr : emptyReg; // @[ringbuffer.scala 48:45 51:15 23:25]
  wire  _GEN_6 = _T ? 1'h0 : _GEN_4; // @[ringbuffer.scala 43:45 45:15]
  wire  _GEN_20 = io_enq_valid & io_enq_ready & io_deq_valid & io_deq_ready ? emptyReg : _GEN_6; // @[ringbuffer.scala 23:25 39:70]
  assign memReg_io_deq_bits_MPORT_en = 1'h1;
  assign memReg_io_deq_bits_MPORT_addr = readPtr;
  assign memReg_io_deq_bits_MPORT_data = memReg[memReg_io_deq_bits_MPORT_addr]; // @[ringbuffer.scala 19:20]
  assign memReg_MPORT_data = io_enq_bits;
  assign memReg_MPORT_addr = writePtr;
  assign memReg_MPORT_mask = 1'h1;
  assign memReg_MPORT_en = _T_1 & io_deq_ready;
  assign memReg_MPORT_1_data = io_enq_bits;
  assign memReg_MPORT_1_addr = writePtr;
  assign memReg_MPORT_1_mask = 1'h1;
  assign memReg_MPORT_1_en = _T_2 ? 1'h0 : _T;
  assign io_enq_ready = ~fullReg | io_deq_ready & io_deq_valid; // @[ringbuffer.scala 56:29]
  assign io_deq_valid = ~emptyReg; // @[ringbuffer.scala 57:20]
  assign io_deq_bits = memReg_io_deq_bits_MPORT_data; // @[ringbuffer.scala 54:16]
  always @(posedge clock) begin
    if (memReg_MPORT_en & memReg_MPORT_mask) begin
      memReg[memReg_MPORT_addr] <= memReg_MPORT_data; // @[ringbuffer.scala 19:20]
    end
    if (memReg_MPORT_1_en & memReg_MPORT_1_mask) begin
      memReg[memReg_MPORT_1_addr] <= memReg_MPORT_1_data; // @[ringbuffer.scala 19:20]
    end
    if (reset) begin // @[ringbuffer.scala 14:24]
      readPtr <= 5'h0; // @[ringbuffer.scala 14:24]
    end else if (incrRead) begin // @[ringbuffer.scala 31:19]
      if (readPtr == 5'h1f) begin // @[ringbuffer.scala 16:21]
        readPtr <= 5'h0;
      end else begin
        readPtr <= _nextRead_T_2;
      end
    end
    if (reset) begin // @[ringbuffer.scala 15:25]
      writePtr <= 5'h0; // @[ringbuffer.scala 15:25]
    end else if (incrWrite) begin // @[ringbuffer.scala 35:20]
      if (writePtr == 5'h1f) begin // @[ringbuffer.scala 17:22]
        writePtr <= 5'h0;
      end else begin
        writePtr <= _nextWrite_T_2;
      end
    end
    if (reset) begin // @[ringbuffer.scala 22:24]
      fullReg <= 1'h0; // @[ringbuffer.scala 22:24]
    end else if (!(io_enq_valid & io_enq_ready & io_deq_valid & io_deq_ready)) begin // @[ringbuffer.scala 39:70]
      if (_T) begin // @[ringbuffer.scala 43:45]
        fullReg <= nextWrite == readPtr; // @[ringbuffer.scala 46:14]
      end else if (io_deq_valid & io_deq_ready) begin // @[ringbuffer.scala 48:45]
        fullReg <= 1'h0; // @[ringbuffer.scala 50:14]
      end
    end
    emptyReg <= reset | _GEN_20; // @[ringbuffer.scala 23:{25,25}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {3{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    memReg[initvar] = _RAND_0[69:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  readPtr = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  writePtr = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  fullReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  emptyReg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ccu(
  input         clock,
  input         reset,
  output        deq_ready,
  input         deq_valid,
  input  [69:0] deq_data,
  output        L2_AWVALID,
  input         L2_AWREADY,
  output [1:0]  L2_AWID,
  output [63:0] L2_AWADDR,
  output        L2_ARVALID,
  input         L2_ARREADY,
  output [1:0]  L2_ARID,
  output [63:0] L2_ARADDR,
  output        L2_WVALID,
  input         L2_WREADY,
  output [63:0] L2_WDATA,
  output        L2_WLAST,
  input         L2_RVALID,
  output        L2_RREADY,
  input  [63:0] L2_RDATA,
  input  [1:0]  L2_RRESP,
  input         L2_RLAST,
  input         L2_BVALID,
  output        L2_BREADY,
  input  [1:0]  L2_BID,
  input  [1:0]  L2_BRESP,
  output        core0_ACVALID,
  input         core0_ACREADY,
  output [63:0] core0_ACADDR,
  output [3:0]  core0_ACSNOOP,
  input         core0_CRVALID,
  output        core0_CRREADY,
  input  [4:0]  core0_CRRESP,
  input         core0_CDVALID,
  output        core0_CDREADY,
  input  [63:0] core0_CDDATA,
  input         core0_CDLAST,
  output        core0_RVALID,
  input         core0_RREADY,
  output [63:0] core0_RDATA,
  output [3:0]  core0_RRESP,
  output        core0_RLAST,
  output        core0_BVALID,
  input         core0_BREADY,
  output [1:0]  core0_BRESP,
  output        core1_RVALID,
  input         core1_RREADY,
  output [63:0] core1_RDATA,
  output        core1_RLAST,
  output        core1_BVALID,
  input         core1_BREADY
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] stateReg_1; // @[ccu.scala 236:33]
  reg [2:0] stateReg_2; // @[ccu.scala 237:33]
  reg [1:0] coreid_reg; // @[ccu.scala 239:33]
  wire [2:0] _GEN_0 = deq_valid & deq_data[3:0] == 4'h8 ? 3'h7 : 3'h0; // @[ccu.scala 247:92 248:52 250:52]
  wire [1:0] _GEN_3 = L2_AWREADY ? 2'h2 : 2'h1; // @[ccu.scala 258:41 259:44 261:44]
  wire [2:0] _GEN_4 = deq_valid ? 3'h4 : 3'h3; // @[ccu.scala 270:40 271:44 273:44]
  wire [2:0] _GEN_5 = L2_WREADY ? 3'h5 : 3'h4; // @[ccu.scala 277:40 278:44 280:44]
  wire [2:0] _GEN_6 = deq_data[0] ? 3'h6 : 3'h3; // @[ccu.scala 285:42 286:44 288:44]
  wire [2:0] _GEN_7 = stateReg_2 == 3'h7 ? 3'h0 : 3'h7; // @[ccu.scala 296:59 297:44 299:44]
  wire [2:0] _GEN_8 = 3'h7 == stateReg_1 ? _GEN_7 : stateReg_1; // @[ccu.scala 242:27 236:33]
  wire [1:0] _GEN_10 = 3'h7 == stateReg_1 ? deq_data[69:68] : coreid_reg; // @[ccu.scala 242:27 239:33 302:36]
  wire [2:0] _GEN_11 = 3'h6 == stateReg_1 ? 3'h0 : _GEN_8; // @[ccu.scala 242:27 293:36]
  wire  _GEN_12 = 3'h6 == stateReg_1 ? 1'h0 : 3'h7 == stateReg_1; // @[ccu.scala 234:15 242:27]
  wire [1:0] _GEN_13 = 3'h6 == stateReg_1 ? coreid_reg : _GEN_10; // @[ccu.scala 242:27 239:33]
  wire [2:0] _GEN_14 = 3'h5 == stateReg_1 ? _GEN_6 : _GEN_11; // @[ccu.scala 242:27]
  wire  _GEN_15 = 3'h5 == stateReg_1 | _GEN_12; // @[ccu.scala 242:27 290:31]
  wire [1:0] _GEN_16 = 3'h5 == stateReg_1 ? coreid_reg : _GEN_13; // @[ccu.scala 242:27 239:33]
  wire [2:0] _GEN_17 = 3'h4 == stateReg_1 ? _GEN_5 : _GEN_14; // @[ccu.scala 242:27]
  wire  _GEN_19 = 3'h4 == stateReg_1 ? 1'h0 : _GEN_15; // @[ccu.scala 234:15 242:27]
  wire [1:0] _GEN_20 = 3'h4 == stateReg_1 ? coreid_reg : _GEN_16; // @[ccu.scala 242:27 239:33]
  wire [2:0] _GEN_21 = 3'h3 == stateReg_1 ? _GEN_4 : _GEN_17; // @[ccu.scala 242:27]
  wire  _GEN_22 = 3'h3 == stateReg_1 ? 1'h0 : 3'h4 == stateReg_1; // @[ccu.scala 193:19 242:27]
  wire  _GEN_23 = 3'h3 == stateReg_1 ? 1'h0 : _GEN_19; // @[ccu.scala 234:15 242:27]
  wire [1:0] _GEN_24 = 3'h3 == stateReg_1 ? coreid_reg : _GEN_20; // @[ccu.scala 242:27 239:33]
  wire  _GEN_26 = 3'h2 == stateReg_1 | _GEN_23; // @[ccu.scala 242:27 267:31]
  wire  _GEN_27 = 3'h2 == stateReg_1 ? 1'h0 : _GEN_22; // @[ccu.scala 193:19 242:27]
  wire  _GEN_31 = 3'h1 == stateReg_1 ? 1'h0 : _GEN_26; // @[ccu.scala 234:15 242:27]
  wire  _GEN_32 = 3'h1 == stateReg_1 ? 1'h0 : _GEN_27; // @[ccu.scala 193:19 242:27]
  wire  deq_1 = 3'h0 == stateReg_1 ? 1'h0 : _GEN_31; // @[ccu.scala 234:15 242:27]
  wire [1:0] _GEN_41 = L2_BID == 2'h0 ? 2'h2 : 2'h3; // @[ccu.scala 320:60 321:44 323:44]
  wire [1:0] _GEN_42 = ~L2_BVALID ? 2'h1 : _GEN_41; // @[ccu.scala 318:41 319:44]
  wire [1:0] _GEN_43 = core0_BREADY ? 2'h0 : 2'h2; // @[ccu.scala 328:43 329:44 331:44]
  wire  _T_26 = coreid_reg == 2'h0; // @[ccu.scala 344:41]
  wire [2:0] _GEN_46 = coreid_reg == 2'h0 & core0_BREADY ? 3'h7 : 3'h6; // @[ccu.scala 344:74 345:44]
  wire  _GEN_48 = _T_26 ? 1'h0 : 1'h1; // @[ccu.scala 218:22 352:58 355:46]
  wire [2:0] _GEN_49 = 3'h7 == stateReg_2 ? 3'h0 : stateReg_2; // @[ccu.scala 307:23 237:33 359:36]
  wire [2:0] _GEN_50 = 3'h6 == stateReg_2 ? _GEN_46 : _GEN_49; // @[ccu.scala 307:23]
  wire  _GEN_52 = 3'h6 == stateReg_2 & _GEN_48; // @[ccu.scala 218:22 307:23]
  wire [2:0] _GEN_53 = 3'h3 == stateReg_2 ? 3'h3 : _GEN_50; // @[ccu.scala 307:23]
  wire  _GEN_54 = 3'h3 == stateReg_2 | _GEN_52; // @[ccu.scala 307:23 341:38]
  wire  _GEN_55 = 3'h3 == stateReg_2 ? 1'h0 : 3'h6 == stateReg_2 & _T_26; // @[ccu.scala 211:22 307:23]
  wire  _GEN_57 = 3'h2 == stateReg_2 | _GEN_55; // @[ccu.scala 307:23 333:38]
  wire  _GEN_58 = 3'h2 == stateReg_2 ? 1'h0 : _GEN_54; // @[ccu.scala 218:22 307:23]
  wire  _GEN_61 = 3'h1 == stateReg_2 ? 1'h0 : _GEN_57; // @[ccu.scala 211:22 307:23]
  wire  _GEN_62 = 3'h1 == stateReg_2 ? 1'h0 : _GEN_58; // @[ccu.scala 218:22 307:23]
  reg [1:0] core_id_pbuf_1; // @[ccu.scala 370:33]
  reg [3:0] tran_pbuf_1; // @[ccu.scala 371:30]
  reg [63:0] addr_pbuf_1; // @[ccu.scala 372:30]
  reg [1:0] core_id_pbuf_2; // @[ccu.scala 375:33]
  reg [3:0] tran_pbuf_2; // @[ccu.scala 376:30]
  reg [63:0] addr_pbuf_2; // @[ccu.scala 377:30]
  reg [4:0] crpbuf_2_0; // @[ccu.scala 378:25]
  reg [1:0] core_id_pbuf_3; // @[ccu.scala 383:33]
  reg [3:0] tran_pbuf_3; // @[ccu.scala 384:30]
  reg [4:0] crpbuf_3_0; // @[ccu.scala 385:25]
  reg [2:0] stateReg_3; // @[ccu.scala 390:33]
  reg [2:0] stateReg_4; // @[ccu.scala 391:29]
  reg [2:0] stateReg_5; // @[ccu.scala 392:29]
  reg [2:0] stateReg_8; // @[ccu.scala 395:29]
  wire [1:0] _GEN_67 = deq_valid & (deq_data[3:0] == 4'h4 | deq_data[3:0] == 4'hb) ? 2'h2 : 2'h0; // @[ccu.scala 404:132 405:52 407:52]
  wire [1:0] _GEN_68 = deq_valid & (deq_data[3:0] == 4'h1 | deq_data[3:0] == 4'h7 | deq_data[3:0] == 4'h0) ? 2'h1 :
    _GEN_67; // @[ccu.scala 402:164 403:52]
  wire [1:0] _GEN_69 = stateReg_1 == 3'h0 ? _GEN_68 : 2'h0; // @[ccu.scala 401:59 410:44]
  wire [1:0] _GEN_70 = ~L2_ARREADY ? 2'h1 : 2'h2; // @[ccu.scala 415:42 416:44 418:44]
  wire [2:0] _GEN_71 = stateReg_4 == 3'h0 & stateReg_5 == 3'h0 ? 3'h5 : 3'h4; // @[ccu.scala 433:91 434:44 436:44]
  wire  _T_59 = stateReg_8 == 3'h7; // @[ccu.scala 446:41]
  wire [2:0] _GEN_72 = stateReg_8 == 3'h7 ? 3'h0 : 3'h6; // @[ccu.scala 446:59 447:44 449:44]
  wire [2:0] _GEN_73 = 3'h6 == stateReg_3 ? _GEN_72 : stateReg_3; // @[ccu.scala 399:23 390:33]
  wire [1:0] _GEN_74 = 3'h5 == stateReg_3 ? core_id_pbuf_1 : core_id_pbuf_2; // @[ccu.scala 399:23 375:33 440:40]
  wire [3:0] _GEN_75 = 3'h5 == stateReg_3 ? tran_pbuf_1 : tran_pbuf_2; // @[ccu.scala 399:23 376:30 441:37]
  wire [63:0] _GEN_76 = 3'h5 == stateReg_3 ? addr_pbuf_1 : addr_pbuf_2; // @[ccu.scala 399:23 377:30 442:37]
  wire [2:0] _GEN_77 = 3'h5 == stateReg_3 ? 3'h6 : _GEN_73; // @[ccu.scala 399:23 443:36]
  wire [2:0] _GEN_78 = 3'h4 == stateReg_3 ? _GEN_71 : _GEN_77; // @[ccu.scala 399:23]
  wire [1:0] _GEN_79 = 3'h4 == stateReg_3 ? core_id_pbuf_2 : _GEN_74; // @[ccu.scala 399:23 375:33]
  wire [3:0] _GEN_80 = 3'h4 == stateReg_3 ? tran_pbuf_2 : _GEN_75; // @[ccu.scala 399:23 376:30]
  wire [63:0] _GEN_81 = 3'h4 == stateReg_3 ? addr_pbuf_2 : _GEN_76; // @[ccu.scala 399:23 377:30]
  wire [2:0] _GEN_83 = 3'h3 == stateReg_3 ? 3'h4 : _GEN_78; // @[ccu.scala 399:23 430:36]
  wire [1:0] _GEN_84 = 3'h3 == stateReg_3 ? core_id_pbuf_2 : _GEN_79; // @[ccu.scala 399:23 375:33]
  wire [3:0] _GEN_85 = 3'h3 == stateReg_3 ? tran_pbuf_2 : _GEN_80; // @[ccu.scala 399:23 376:30]
  wire [63:0] _GEN_86 = 3'h3 == stateReg_3 ? addr_pbuf_2 : _GEN_81; // @[ccu.scala 399:23 377:30]
  wire  _GEN_91 = 3'h2 == stateReg_3 ? 1'h0 : 3'h3 == stateReg_3; // @[ccu.scala 367:15 399:23]
  wire  _GEN_100 = 3'h1 == stateReg_3 ? 1'h0 : _GEN_91; // @[ccu.scala 367:15 399:23]
  wire  deq_3 = 3'h0 == stateReg_3 ? 1'h0 : _GEN_100; // @[ccu.scala 367:15 399:23]
  wire  _T_61 = stateReg_3 == 3'h6; // @[ccu.scala 465:42]
  wire  _T_65 = stateReg_3 == 3'h6 & (tran_pbuf_2 == 4'h4 | tran_pbuf_2 == 4'h0); // @[ccu.scala 465:61]
  wire  _T_67 = core_id_pbuf_2 == 2'h0; // @[ccu.scala 467:86]
  wire  _T_72 = _T_61 & ~_T_67; // @[ccu.scala 469:67]
  wire [1:0] _GEN_116 = ~core0_ACREADY ? 2'h1 : 2'h2; // @[ccu.scala 477:45 478:44 480:44]
  wire [3:0] _GEN_117 = tran_pbuf_2 == 4'hb ? 4'h9 : 4'h0; // @[ccu.scala 488:67 489:47 491:47]
  wire [3:0] _GEN_118 = tran_pbuf_2 == 4'h7 ? 4'h7 : _GEN_117; // @[ccu.scala 486:67 487:47]
  wire [3:0] _GEN_119 = tran_pbuf_2 == 4'h1 ? 4'h1 : _GEN_118; // @[ccu.scala 484:61 485:47]
  wire [1:0] _GEN_120 = ~core0_CRVALID ? 2'h2 : 2'h3; // @[ccu.scala 496:45 497:44 499:44]
  wire [2:0] _GEN_121 = stateReg_4 == 3'h4 & stateReg_5 == 3'h4 ? 3'h5 : 3'h4; // @[ccu.scala 508:95 509:44 511:44]
  wire [2:0] _GEN_122 = stateReg_8 == 3'h0 ? 3'h6 : 3'h5; // @[ccu.scala 515:59 516:44 518:44]
  wire [2:0] _GEN_123 = _T_59 ? 3'h0 : 3'h7; // @[ccu.scala 528:59 529:44 531:44]
  wire [2:0] _GEN_124 = 3'h7 == stateReg_4 ? _GEN_123 : stateReg_4; // @[ccu.scala 463:27 391:29]
  wire [1:0] _GEN_125 = 3'h6 == stateReg_4 ? core_id_pbuf_2 : core_id_pbuf_3; // @[ccu.scala 463:27 383:33 522:40]
  wire [3:0] _GEN_126 = 3'h6 == stateReg_4 ? tran_pbuf_2 : tran_pbuf_3; // @[ccu.scala 463:27 384:30 523:37]
  wire [4:0] _GEN_127 = 3'h6 == stateReg_4 ? crpbuf_2_0 : crpbuf_3_0; // @[ccu.scala 385:25 463:27 524:36]
  wire [2:0] _GEN_128 = 3'h6 == stateReg_4 ? 3'h7 : _GEN_124; // @[ccu.scala 463:27 525:36]
  wire [2:0] _GEN_129 = 3'h5 == stateReg_4 ? _GEN_122 : _GEN_128; // @[ccu.scala 463:27]
  wire [1:0] _GEN_130 = 3'h5 == stateReg_4 ? core_id_pbuf_3 : _GEN_125; // @[ccu.scala 463:27 383:33]
  wire [3:0] _GEN_131 = 3'h5 == stateReg_4 ? tran_pbuf_3 : _GEN_126; // @[ccu.scala 463:27 384:30]
  wire [4:0] _GEN_132 = 3'h5 == stateReg_4 ? crpbuf_3_0 : _GEN_127; // @[ccu.scala 385:25 463:27]
  wire [2:0] _GEN_133 = 3'h4 == stateReg_4 ? _GEN_121 : _GEN_129; // @[ccu.scala 463:27]
  wire [1:0] _GEN_134 = 3'h4 == stateReg_4 ? core_id_pbuf_3 : _GEN_130; // @[ccu.scala 463:27 383:33]
  wire [3:0] _GEN_135 = 3'h4 == stateReg_4 ? tran_pbuf_3 : _GEN_131; // @[ccu.scala 463:27 384:30]
  wire [4:0] _GEN_136 = 3'h4 == stateReg_4 ? crpbuf_3_0 : _GEN_132; // @[ccu.scala 385:25 463:27]
  wire [2:0] _GEN_138 = 3'h3 == stateReg_4 ? 3'h4 : _GEN_133; // @[ccu.scala 463:27 505:36]
  wire [1:0] _GEN_139 = 3'h3 == stateReg_4 ? core_id_pbuf_3 : _GEN_134; // @[ccu.scala 463:27 383:33]
  wire [3:0] _GEN_140 = 3'h3 == stateReg_4 ? tran_pbuf_3 : _GEN_135; // @[ccu.scala 463:27 384:30]
  wire  _GEN_144 = 3'h2 == stateReg_4 ? 1'h0 : 3'h3 == stateReg_4; // @[ccu.scala 461:23 463:27]
  wire [3:0] _GEN_150 = 3'h1 == stateReg_4 ? _GEN_119 : 4'h0; // @[ccu.scala 459:23 463:27]
  wire  _GEN_152 = 3'h1 == stateReg_4 ? 1'h0 : _GEN_144; // @[ccu.scala 461:23 463:27]
  wire  _T_97 = core_id_pbuf_2 == 2'h1; // @[ccu.scala 548:86]
  wire  _T_102 = _T_61 & ~_T_97; // @[ccu.scala 550:67]
  wire [2:0] _GEN_175 = 3'h7 == stateReg_5 ? _GEN_123 : stateReg_5; // @[ccu.scala 544:27 392:29]
  wire [2:0] _GEN_177 = 3'h6 == stateReg_5 ? 3'h7 : _GEN_175; // @[ccu.scala 544:27 605:36]
  wire [2:0] _GEN_178 = 3'h5 == stateReg_5 ? _GEN_122 : _GEN_177; // @[ccu.scala 544:27]
  wire [2:0] _GEN_180 = 3'h4 == stateReg_5 ? _GEN_121 : _GEN_178; // @[ccu.scala 544:27]
  wire [2:0] _GEN_183 = 3'h3 == stateReg_5 ? 3'h4 : _GEN_180; // @[ccu.scala 544:27 587:36]
  reg [2:0] select_buff; // @[ccu.scala 618:38]
  reg [63:0] beat_buff; // @[ccu.scala 619:36]
  reg  last_buff; // @[ccu.scala 620:36]
  reg [3:0] rsp_buff; // @[ccu.scala 621:31]
  wire  _T_121 = stateReg_4 == 3'h7; // @[ccu.scala 636:41]
  wire [1:0] _GEN_205 = (~crpbuf_3_0[0] | core0_CDVALID) & L2_RVALID ? 2'h3 : 2'h2; // @[ccu.scala 655:114 656:44 658:44]
  wire [3:0] _rsp_buff_T_2 = {crpbuf_3_0[3],crpbuf_3_0[2],2'h0}; // @[Cat.scala 33:92]
  wire [3:0] _rsp_buff_T_6 = {2'h0,L2_RRESP}; // @[Cat.scala 33:92]
  wire [63:0] _GEN_206 = select_buff == 3'h1 ? 64'h0 : L2_RDATA; // @[ccu.scala 668:66 669:43 673:43]
  wire  _GEN_207 = select_buff == 3'h1 ? 1'h0 : L2_RLAST; // @[ccu.scala 668:66 670:43 674:43]
  wire [3:0] _GEN_208 = select_buff == 3'h1 ? 4'h0 : _rsp_buff_T_6; // @[ccu.scala 668:66 671:42 675:42]
  wire [63:0] _GEN_209 = select_buff == 3'h0 ? core0_CDDATA : _GEN_206; // @[ccu.scala 664:60 665:43]
  wire  _GEN_210 = select_buff == 3'h0 ? core0_CDLAST : _GEN_207; // @[ccu.scala 664:60 666:43]
  wire [3:0] _GEN_211 = select_buff == 3'h0 ? _rsp_buff_T_2 : _GEN_208; // @[ccu.scala 664:60 667:42]
  wire  _T_152 = core_id_pbuf_3 == 2'h0; // @[ccu.scala 695:49]
  wire  _T_156 = core_id_pbuf_3 == 2'h0 & core0_RREADY | core_id_pbuf_3 == 2'h1 & core1_RREADY; // @[ccu.scala 695:84]
  wire [2:0] _GEN_214 = last_buff ? 3'h7 : 3'h2; // @[ccu.scala 697:46 698:44 700:44]
  wire [2:0] _GEN_215 = ~(core_id_pbuf_3 == 2'h0 & core0_RREADY | core_id_pbuf_3 == 2'h1 & core1_RREADY) ? 3'h5 :
    _GEN_214; // @[ccu.scala 695:140 696:44]
  wire  _GEN_217 = _T_152 ? 1'h0 : 1'h1; // @[ccu.scala 628:22 704:62 707:46]
  wire [2:0] _GEN_218 = _T_156 ? 3'h7 : 3'h6; // @[ccu.scala 711:137 712:44 714:44]
  wire [2:0] _GEN_221 = 3'h7 == stateReg_8 ? 3'h0 : stateReg_8; // @[ccu.scala 634:27 395:29 729:36]
  wire [2:0] _GEN_222 = 3'h6 == stateReg_8 ? _GEN_218 : _GEN_221; // @[ccu.scala 634:27]
  wire  _GEN_223 = 3'h6 == stateReg_8 & _T_152; // @[ccu.scala 622:22 634:27]
  wire  _GEN_224 = 3'h6 == stateReg_8 & _GEN_217; // @[ccu.scala 628:22 634:27]
  wire [3:0] _GEN_225 = 3'h6 == stateReg_8 ? 4'h0 : rsp_buff; // @[ccu.scala 626:21 634:27 725:37]
  wire [2:0] _GEN_226 = 3'h5 == stateReg_8 ? _GEN_215 : _GEN_222; // @[ccu.scala 634:27]
  wire  _GEN_227 = 3'h5 == stateReg_8 ? _T_152 : _GEN_223; // @[ccu.scala 634:27]
  wire  _GEN_228 = 3'h5 == stateReg_8 ? _GEN_217 : _GEN_224; // @[ccu.scala 634:27]
  wire [3:0] _GEN_229 = 3'h5 == stateReg_8 ? rsp_buff : _GEN_225; // @[ccu.scala 626:21 634:27]
  wire [2:0] _GEN_230 = 3'h4 == stateReg_8 ? 3'h5 : _GEN_226; // @[ccu.scala 634:27 680:36]
  wire  _GEN_234 = 3'h4 == stateReg_8 ? 1'h0 : _GEN_227; // @[ccu.scala 622:22 634:27]
  wire  _GEN_235 = 3'h4 == stateReg_8 ? 1'h0 : _GEN_228; // @[ccu.scala 628:22 634:27]
  wire [3:0] _GEN_236 = 3'h4 == stateReg_8 ? rsp_buff : _GEN_229; // @[ccu.scala 626:21 634:27]
  wire [2:0] _GEN_237 = 3'h3 == stateReg_8 ? 3'h4 : _GEN_230; // @[ccu.scala 634:27 663:36]
  wire [63:0] _GEN_238 = 3'h3 == stateReg_8 ? _GEN_209 : beat_buff; // @[ccu.scala 634:27 619:36]
  wire  _GEN_239 = 3'h3 == stateReg_8 ? _GEN_210 : last_buff; // @[ccu.scala 634:27 620:36]
  wire [3:0] _GEN_240 = 3'h3 == stateReg_8 ? _GEN_211 : rsp_buff; // @[ccu.scala 634:27 621:31]
  wire  _GEN_241 = 3'h3 == stateReg_8 ? 1'h0 : 3'h4 == stateReg_8 & crpbuf_3_0[0]; // @[ccu.scala 215:23 634:27]
  wire  _GEN_243 = 3'h3 == stateReg_8 ? 1'h0 : 3'h4 == stateReg_8; // @[ccu.scala 203:19 634:27]
  wire  _GEN_244 = 3'h3 == stateReg_8 ? 1'h0 : _GEN_234; // @[ccu.scala 622:22 634:27]
  wire  _GEN_245 = 3'h3 == stateReg_8 ? 1'h0 : _GEN_235; // @[ccu.scala 628:22 634:27]
  wire [3:0] _GEN_246 = 3'h3 == stateReg_8 ? rsp_buff : _GEN_236; // @[ccu.scala 626:21 634:27]
  wire  _GEN_251 = 3'h2 == stateReg_8 ? 1'h0 : _GEN_241; // @[ccu.scala 215:23 634:27]
  wire  _GEN_253 = 3'h2 == stateReg_8 ? 1'h0 : _GEN_243; // @[ccu.scala 203:19 634:27]
  wire  _GEN_254 = 3'h2 == stateReg_8 ? 1'h0 : _GEN_244; // @[ccu.scala 622:22 634:27]
  wire  _GEN_255 = 3'h2 == stateReg_8 ? 1'h0 : _GEN_245; // @[ccu.scala 628:22 634:27]
  wire [3:0] _GEN_256 = 3'h2 == stateReg_8 ? rsp_buff : _GEN_246; // @[ccu.scala 626:21 634:27]
  wire  _GEN_262 = 3'h1 == stateReg_8 ? 1'h0 : _GEN_251; // @[ccu.scala 215:23 634:27]
  wire  _GEN_264 = 3'h1 == stateReg_8 ? 1'h0 : _GEN_253; // @[ccu.scala 203:19 634:27]
  wire  _GEN_265 = 3'h1 == stateReg_8 ? 1'h0 : _GEN_254; // @[ccu.scala 622:22 634:27]
  wire  _GEN_266 = 3'h1 == stateReg_8 ? 1'h0 : _GEN_255; // @[ccu.scala 628:22 634:27]
  wire [3:0] _GEN_267 = 3'h1 == stateReg_8 ? rsp_buff : _GEN_256; // @[ccu.scala 626:21 634:27]
  assign deq_ready = deq_1 | deq_3; // @[ccu.scala 454:28]
  assign L2_AWVALID = 3'h0 == stateReg_1 ? 1'h0 : 3'h1 == stateReg_1; // @[ccu.scala 190:20 242:27]
  assign L2_AWID = deq_data[69:68]; // @[ccu.scala 191:28]
  assign L2_AWADDR = deq_data[67:4]; // @[ccu.scala 192:30]
  assign L2_ARVALID = 3'h0 == stateReg_3 ? 1'h0 : 3'h1 == stateReg_3; // @[ccu.scala 198:20 399:23]
  assign L2_ARID = deq_data[69:68]; // @[ccu.scala 200:28]
  assign L2_ARADDR = deq_data[67:4]; // @[ccu.scala 199:30]
  assign L2_WVALID = 3'h0 == stateReg_1 ? 1'h0 : _GEN_32; // @[ccu.scala 193:19 242:27]
  assign L2_WDATA = deq_data[67:4]; // @[ccu.scala 194:29]
  assign L2_WLAST = deq_data[0]; // @[ccu.scala 195:29]
  assign L2_RREADY = 3'h0 == stateReg_8 ? 1'h0 : _GEN_264; // @[ccu.scala 203:19 634:27]
  assign L2_BREADY = 3'h0 == stateReg_2 ? 1'h0 : 3'h1 == stateReg_2; // @[ccu.scala 206:19 307:23]
  assign core0_ACVALID = 3'h0 == stateReg_4 ? 1'h0 : 3'h1 == stateReg_4; // @[ccu.scala 457:23 463:27]
  assign core0_ACADDR = addr_pbuf_2; // @[ccu.scala 458:22]
  assign core0_ACSNOOP = 3'h0 == stateReg_4 ? 4'h0 : _GEN_150; // @[ccu.scala 459:23 463:27]
  assign core0_CRREADY = 3'h0 == stateReg_4 ? 1'h0 : _GEN_152; // @[ccu.scala 461:23 463:27]
  assign core0_CDREADY = 3'h0 == stateReg_8 ? 1'h0 : _GEN_262; // @[ccu.scala 215:23 634:27]
  assign core0_RVALID = 3'h0 == stateReg_8 ? 1'h0 : _GEN_265; // @[ccu.scala 622:22 634:27]
  assign core0_RDATA = beat_buff; // @[ccu.scala 624:21]
  assign core0_RRESP = 3'h0 == stateReg_8 ? rsp_buff : _GEN_267; // @[ccu.scala 626:21 634:27]
  assign core0_RLAST = last_buff; // @[ccu.scala 625:21]
  assign core0_BVALID = 3'h0 == stateReg_2 ? 1'h0 : _GEN_61; // @[ccu.scala 211:22 307:23]
  assign core0_BRESP = L2_BRESP; // @[ccu.scala 212:21]
  assign core1_RVALID = 3'h0 == stateReg_8 ? 1'h0 : _GEN_266; // @[ccu.scala 628:22 634:27]
  assign core1_RDATA = beat_buff; // @[ccu.scala 630:21]
  assign core1_RLAST = last_buff; // @[ccu.scala 631:21]
  assign core1_BVALID = 3'h0 == stateReg_2 ? 1'h0 : _GEN_62; // @[ccu.scala 218:22 307:23]
  always @(posedge clock) begin
    if (reset) begin // @[ccu.scala 236:33]
      stateReg_1 <= 3'h0; // @[ccu.scala 236:33]
    end else if (3'h0 == stateReg_1) begin // @[ccu.scala 242:27]
      if (stateReg_2 == 3'h0) begin // @[ccu.scala 244:59]
        if (deq_valid & deq_data[3:0] == 4'h3) begin // @[ccu.scala 245:86]
          stateReg_1 <= 3'h1; // @[ccu.scala 246:52]
        end else begin
          stateReg_1 <= _GEN_0;
        end
      end else begin
        stateReg_1 <= 3'h0; // @[ccu.scala 253:44]
      end
    end else if (3'h1 == stateReg_1) begin // @[ccu.scala 242:27]
      stateReg_1 <= {{1'd0}, _GEN_3};
    end else if (3'h2 == stateReg_1) begin // @[ccu.scala 242:27]
      stateReg_1 <= 3'h3; // @[ccu.scala 266:36]
    end else begin
      stateReg_1 <= _GEN_21;
    end
    if (reset) begin // @[ccu.scala 237:33]
      stateReg_2 <= 3'h0; // @[ccu.scala 237:33]
    end else if (3'h0 == stateReg_2) begin // @[ccu.scala 307:23]
      if (stateReg_1 == 3'h6) begin // @[ccu.scala 309:59]
        stateReg_2 <= 3'h1; // @[ccu.scala 310:44]
      end else if (stateReg_1 == 3'h7) begin // @[ccu.scala 311:65]
        stateReg_2 <= 3'h6; // @[ccu.scala 312:44]
      end else begin
        stateReg_2 <= 3'h0; // @[ccu.scala 314:44]
      end
    end else if (3'h1 == stateReg_2) begin // @[ccu.scala 307:23]
      stateReg_2 <= {{1'd0}, _GEN_42};
    end else if (3'h2 == stateReg_2) begin // @[ccu.scala 307:23]
      stateReg_2 <= {{1'd0}, _GEN_43};
    end else begin
      stateReg_2 <= _GEN_53;
    end
    if (reset) begin // @[ccu.scala 239:33]
      coreid_reg <= 2'h0; // @[ccu.scala 239:33]
    end else if (!(3'h0 == stateReg_1)) begin // @[ccu.scala 242:27]
      if (!(3'h1 == stateReg_1)) begin // @[ccu.scala 242:27]
        if (!(3'h2 == stateReg_1)) begin // @[ccu.scala 242:27]
          coreid_reg <= _GEN_24;
        end
      end
    end
    if (reset) begin // @[ccu.scala 370:33]
      core_id_pbuf_1 <= 2'h0; // @[ccu.scala 370:33]
    end else if (!(3'h0 == stateReg_3)) begin // @[ccu.scala 399:23]
      if (!(3'h1 == stateReg_3)) begin // @[ccu.scala 399:23]
        if (3'h2 == stateReg_3) begin // @[ccu.scala 399:23]
          core_id_pbuf_1 <= deq_data[69:68]; // @[ccu.scala 423:40]
        end
      end
    end
    if (reset) begin // @[ccu.scala 371:30]
      tran_pbuf_1 <= 4'h0; // @[ccu.scala 371:30]
    end else if (!(3'h0 == stateReg_3)) begin // @[ccu.scala 399:23]
      if (!(3'h1 == stateReg_3)) begin // @[ccu.scala 399:23]
        if (3'h2 == stateReg_3) begin // @[ccu.scala 399:23]
          tran_pbuf_1 <= deq_data[3:0]; // @[ccu.scala 424:37]
        end
      end
    end
    if (reset) begin // @[ccu.scala 372:30]
      addr_pbuf_1 <= 64'h0; // @[ccu.scala 372:30]
    end else if (!(3'h0 == stateReg_3)) begin // @[ccu.scala 399:23]
      if (!(3'h1 == stateReg_3)) begin // @[ccu.scala 399:23]
        if (3'h2 == stateReg_3) begin // @[ccu.scala 399:23]
          addr_pbuf_1 <= deq_data[67:4]; // @[ccu.scala 425:37]
        end
      end
    end
    if (reset) begin // @[ccu.scala 375:33]
      core_id_pbuf_2 <= 2'h0; // @[ccu.scala 375:33]
    end else if (!(3'h0 == stateReg_3)) begin // @[ccu.scala 399:23]
      if (!(3'h1 == stateReg_3)) begin // @[ccu.scala 399:23]
        if (!(3'h2 == stateReg_3)) begin // @[ccu.scala 399:23]
          core_id_pbuf_2 <= _GEN_84;
        end
      end
    end
    if (reset) begin // @[ccu.scala 376:30]
      tran_pbuf_2 <= 4'h0; // @[ccu.scala 376:30]
    end else if (!(3'h0 == stateReg_3)) begin // @[ccu.scala 399:23]
      if (!(3'h1 == stateReg_3)) begin // @[ccu.scala 399:23]
        if (!(3'h2 == stateReg_3)) begin // @[ccu.scala 399:23]
          tran_pbuf_2 <= _GEN_85;
        end
      end
    end
    if (reset) begin // @[ccu.scala 377:30]
      addr_pbuf_2 <= 64'h0; // @[ccu.scala 377:30]
    end else if (!(3'h0 == stateReg_3)) begin // @[ccu.scala 399:23]
      if (!(3'h1 == stateReg_3)) begin // @[ccu.scala 399:23]
        if (!(3'h2 == stateReg_3)) begin // @[ccu.scala 399:23]
          addr_pbuf_2 <= _GEN_86;
        end
      end
    end
    if (3'h0 == stateReg_4) begin // @[ccu.scala 463:27]
      crpbuf_2_0 <= 5'h0; // @[ccu.scala 474:36]
    end else if (!(3'h1 == stateReg_4)) begin // @[ccu.scala 463:27]
      if (3'h2 == stateReg_4) begin // @[ccu.scala 463:27]
        crpbuf_2_0 <= core0_CRRESP; // @[ccu.scala 501:36]
      end
    end
    if (reset) begin // @[ccu.scala 383:33]
      core_id_pbuf_3 <= 2'h0; // @[ccu.scala 383:33]
    end else if (!(3'h0 == stateReg_4)) begin // @[ccu.scala 463:27]
      if (!(3'h1 == stateReg_4)) begin // @[ccu.scala 463:27]
        if (!(3'h2 == stateReg_4)) begin // @[ccu.scala 463:27]
          core_id_pbuf_3 <= _GEN_139;
        end
      end
    end
    if (reset) begin // @[ccu.scala 384:30]
      tran_pbuf_3 <= 4'h0; // @[ccu.scala 384:30]
    end else if (!(3'h0 == stateReg_4)) begin // @[ccu.scala 463:27]
      if (!(3'h1 == stateReg_4)) begin // @[ccu.scala 463:27]
        if (!(3'h2 == stateReg_4)) begin // @[ccu.scala 463:27]
          tran_pbuf_3 <= _GEN_140;
        end
      end
    end
    if (!(3'h0 == stateReg_4)) begin // @[ccu.scala 463:27]
      if (!(3'h1 == stateReg_4)) begin // @[ccu.scala 463:27]
        if (!(3'h2 == stateReg_4)) begin // @[ccu.scala 463:27]
          if (!(3'h3 == stateReg_4)) begin // @[ccu.scala 463:27]
            crpbuf_3_0 <= _GEN_136;
          end
        end
      end
    end
    if (reset) begin // @[ccu.scala 390:33]
      stateReg_3 <= 3'h0; // @[ccu.scala 390:33]
    end else if (3'h0 == stateReg_3) begin // @[ccu.scala 399:23]
      stateReg_3 <= {{1'd0}, _GEN_69};
    end else if (3'h1 == stateReg_3) begin // @[ccu.scala 399:23]
      stateReg_3 <= {{1'd0}, _GEN_70};
    end else if (3'h2 == stateReg_3) begin // @[ccu.scala 399:23]
      stateReg_3 <= 3'h3; // @[ccu.scala 426:36]
    end else begin
      stateReg_3 <= _GEN_83;
    end
    if (reset) begin // @[ccu.scala 391:29]
      stateReg_4 <= 3'h0; // @[ccu.scala 391:29]
    end else if (3'h0 == stateReg_4) begin // @[ccu.scala 463:27]
      if (stateReg_3 == 3'h6 & (tran_pbuf_2 == 4'h4 | tran_pbuf_2 == 4'h0)) begin // @[ccu.scala 465:135]
        stateReg_4 <= 3'h4; // @[ccu.scala 466:44]
      end else if (_T_61 & core_id_pbuf_2 == 2'h0) begin // @[ccu.scala 467:104]
        stateReg_4 <= 3'h4; // @[ccu.scala 468:44]
      end else begin
        stateReg_4 <= {{2'd0}, _T_72};
      end
    end else if (3'h1 == stateReg_4) begin // @[ccu.scala 463:27]
      stateReg_4 <= {{1'd0}, _GEN_116};
    end else if (3'h2 == stateReg_4) begin // @[ccu.scala 463:27]
      stateReg_4 <= {{1'd0}, _GEN_120};
    end else begin
      stateReg_4 <= _GEN_138;
    end
    if (reset) begin // @[ccu.scala 392:29]
      stateReg_5 <= 3'h0; // @[ccu.scala 392:29]
    end else if (3'h0 == stateReg_5) begin // @[ccu.scala 544:27]
      if (_T_65) begin // @[ccu.scala 546:135]
        stateReg_5 <= 3'h4; // @[ccu.scala 547:44]
      end else if (_T_61 & core_id_pbuf_2 == 2'h1) begin // @[ccu.scala 548:104]
        stateReg_5 <= 3'h4; // @[ccu.scala 549:44]
      end else begin
        stateReg_5 <= {{2'd0}, _T_102};
      end
    end else if (3'h1 == stateReg_5) begin // @[ccu.scala 544:27]
      stateReg_5 <= 3'h2;
    end else if (3'h2 == stateReg_5) begin // @[ccu.scala 544:27]
      stateReg_5 <= 3'h3;
    end else begin
      stateReg_5 <= _GEN_183;
    end
    if (reset) begin // @[ccu.scala 395:29]
      stateReg_8 <= 3'h0; // @[ccu.scala 395:29]
    end else if (3'h0 == stateReg_8) begin // @[ccu.scala 634:27]
      if (stateReg_4 == 3'h7 & (tran_pbuf_3 == 4'h1 | tran_pbuf_3 == 4'h7 | tran_pbuf_3 == 4'h0)) begin // @[ccu.scala 636:169]
        stateReg_8 <= 3'h1; // @[ccu.scala 637:44]
      end else if (_T_121 & (tran_pbuf_3 == 4'h4 | tran_pbuf_3 == 4'hb)) begin // @[ccu.scala 638:139]
        stateReg_8 <= 3'h6; // @[ccu.scala 639:44]
      end else begin
        stateReg_8 <= 3'h0; // @[ccu.scala 641:44]
      end
    end else if (3'h1 == stateReg_8) begin // @[ccu.scala 634:27]
      stateReg_8 <= 3'h2; // @[ccu.scala 645:36]
    end else if (3'h2 == stateReg_8) begin // @[ccu.scala 634:27]
      stateReg_8 <= {{1'd0}, _GEN_205};
    end else begin
      stateReg_8 <= _GEN_237;
    end
    if (reset) begin // @[ccu.scala 618:38]
      select_buff <= 3'h0; // @[ccu.scala 618:38]
    end else if (!(3'h0 == stateReg_8)) begin // @[ccu.scala 634:27]
      if (3'h1 == stateReg_8) begin // @[ccu.scala 634:27]
        if (crpbuf_3_0[3]) begin // @[ccu.scala 646:44]
          select_buff <= 3'h0; // @[ccu.scala 647:45]
        end else begin
          select_buff <= 3'h4;
        end
      end
    end
    if (reset) begin // @[ccu.scala 619:36]
      beat_buff <= 64'h0; // @[ccu.scala 619:36]
    end else if (!(3'h0 == stateReg_8)) begin // @[ccu.scala 634:27]
      if (!(3'h1 == stateReg_8)) begin // @[ccu.scala 634:27]
        if (!(3'h2 == stateReg_8)) begin // @[ccu.scala 634:27]
          beat_buff <= _GEN_238;
        end
      end
    end
    if (reset) begin // @[ccu.scala 620:36]
      last_buff <= 1'h0; // @[ccu.scala 620:36]
    end else if (!(3'h0 == stateReg_8)) begin // @[ccu.scala 634:27]
      if (!(3'h1 == stateReg_8)) begin // @[ccu.scala 634:27]
        if (!(3'h2 == stateReg_8)) begin // @[ccu.scala 634:27]
          last_buff <= _GEN_239;
        end
      end
    end
    if (reset) begin // @[ccu.scala 621:31]
      rsp_buff <= 4'h0; // @[ccu.scala 621:31]
    end else if (!(3'h0 == stateReg_8)) begin // @[ccu.scala 634:27]
      if (!(3'h1 == stateReg_8)) begin // @[ccu.scala 634:27]
        if (!(3'h2 == stateReg_8)) begin // @[ccu.scala 634:27]
          rsp_buff <= _GEN_240;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stateReg_1 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  stateReg_2 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  coreid_reg = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  core_id_pbuf_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  tran_pbuf_1 = _RAND_4[3:0];
  _RAND_5 = {2{`RANDOM}};
  addr_pbuf_1 = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  core_id_pbuf_2 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  tran_pbuf_2 = _RAND_7[3:0];
  _RAND_8 = {2{`RANDOM}};
  addr_pbuf_2 = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  crpbuf_2_0 = _RAND_9[4:0];
  _RAND_10 = {1{`RANDOM}};
  core_id_pbuf_3 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  tran_pbuf_3 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  crpbuf_3_0 = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  stateReg_3 = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  stateReg_4 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  stateReg_5 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  stateReg_8 = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  select_buff = _RAND_17[2:0];
  _RAND_18 = {2{`RANDOM}};
  beat_buff = _RAND_18[63:0];
  _RAND_19 = {1{`RANDOM}};
  last_buff = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  rsp_buff = _RAND_20[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Interconnect(
  input         clock,
  input         reset,
  input         io_acePort0_AWVALID,
  output        io_acePort0_AWREADY,
  input  [63:0] io_acePort0_AWADDR,
  input  [2:0]  io_acePort0_AWSNOOP,
  input         io_acePort0_WVALID,
  output        io_acePort0_WREADY,
  input  [63:0] io_acePort0_WDATA,
  input         io_acePort0_WLAST,
  output        io_acePort0_BVALID,
  input         io_acePort0_BREADY,
  output [1:0]  io_acePort0_BRESP,
  input         io_acePort0_ARVALID,
  output        io_acePort0_ARREADY,
  input  [63:0] io_acePort0_ARADDR,
  input  [3:0]  io_acePort0_ARSNOOP,
  output        io_acePort0_RVALID,
  input         io_acePort0_RREADY,
  output [63:0] io_acePort0_RDATA,
  output [3:0]  io_acePort0_RRESP,
  output        io_acePort0_RLAST,
  output        io_acePort0_ACVALID,
  input         io_acePort0_ACREADY,
  output [63:0] io_acePort0_ACADDR,
  output [3:0]  io_acePort0_ACSNOOP,
  input         io_acePort0_CRVALID,
  output        io_acePort0_CRREADY,
  input  [4:0]  io_acePort0_CRRESP,
  input         io_acePort0_CDVALID,
  output        io_acePort0_CDREADY,
  input  [63:0] io_acePort0_CDDATA,
  input         io_acePort0_CDLAST,
  input         io_acePort1_ARVALID,
  output        io_acePort1_ARREADY,
  input  [63:0] io_acePort1_ARADDR,
  output        io_acePort1_RVALID,
  input         io_acePort1_RREADY,
  output [63:0] io_acePort1_RDATA,
  output        io_acePort1_RLAST,
  output        io_L2_AWVALID,
  input         io_L2_AWREADY,
  output [1:0]  io_L2_AWID,
  output [63:0] io_L2_AWADDR,
  output        io_L2_ARVALID,
  input         io_L2_ARREADY,
  output [1:0]  io_L2_ARID,
  output [63:0] io_L2_ARADDR,
  output        io_L2_WVALID,
  input         io_L2_WREADY,
  output [63:0] io_L2_WDATA,
  output        io_L2_WLAST,
  input         io_L2_RVALID,
  output        io_L2_RREADY,
  input  [63:0] io_L2_RDATA,
  input  [1:0]  io_L2_RRESP,
  input         io_L2_RLAST,
  input         io_L2_BVALID,
  output        io_L2_BREADY,
  input  [1:0]  io_L2_BID,
  input  [1:0]  io_L2_BRESP
);
  wire  Arbiter_clock; // @[Interconnect.scala 88:23]
  wire  Arbiter_reset; // @[Interconnect.scala 88:23]
  wire  Arbiter_io_AWVALID_0; // @[Interconnect.scala 88:23]
  wire  Arbiter_io_AWREADY_0; // @[Interconnect.scala 88:23]
  wire  Arbiter_io_WVALID_0; // @[Interconnect.scala 88:23]
  wire  Arbiter_io_WLAST_0; // @[Interconnect.scala 88:23]
  wire  Arbiter_io_WREADY_0; // @[Interconnect.scala 88:23]
  wire  Arbiter_io_ARVALID_0; // @[Interconnect.scala 88:23]
  wire  Arbiter_io_ARREADY_0; // @[Interconnect.scala 88:23]
  wire  Arbiter_io_ARVALID_1; // @[Interconnect.scala 88:23]
  wire  Arbiter_io_ARREADY_1; // @[Interconnect.scala 88:23]
  wire [2:0] Arbiter_io_select; // @[Interconnect.scala 88:23]
  wire  Arbiter_io_enq_valid; // @[Interconnect.scala 88:23]
  wire  Arbiter_io_enq_ready; // @[Interconnect.scala 88:23]
  wire  Arbiter_io_nstall; // @[Interconnect.scala 88:23]
  wire  FIFO_clock; // @[Interconnect.scala 112:20]
  wire  FIFO_reset; // @[Interconnect.scala 112:20]
  wire  FIFO_io_enq_ready; // @[Interconnect.scala 112:20]
  wire  FIFO_io_enq_valid; // @[Interconnect.scala 112:20]
  wire [69:0] FIFO_io_enq_bits; // @[Interconnect.scala 112:20]
  wire  FIFO_io_deq_ready; // @[Interconnect.scala 112:20]
  wire  FIFO_io_deq_valid; // @[Interconnect.scala 112:20]
  wire [69:0] FIFO_io_deq_bits; // @[Interconnect.scala 112:20]
  wire  CCU_clock; // @[Interconnect.scala 146:19]
  wire  CCU_reset; // @[Interconnect.scala 146:19]
  wire  CCU_deq_ready; // @[Interconnect.scala 146:19]
  wire  CCU_deq_valid; // @[Interconnect.scala 146:19]
  wire [69:0] CCU_deq_data; // @[Interconnect.scala 146:19]
  wire  CCU_L2_AWVALID; // @[Interconnect.scala 146:19]
  wire  CCU_L2_AWREADY; // @[Interconnect.scala 146:19]
  wire [1:0] CCU_L2_AWID; // @[Interconnect.scala 146:19]
  wire [63:0] CCU_L2_AWADDR; // @[Interconnect.scala 146:19]
  wire  CCU_L2_ARVALID; // @[Interconnect.scala 146:19]
  wire  CCU_L2_ARREADY; // @[Interconnect.scala 146:19]
  wire [1:0] CCU_L2_ARID; // @[Interconnect.scala 146:19]
  wire [63:0] CCU_L2_ARADDR; // @[Interconnect.scala 146:19]
  wire  CCU_L2_WVALID; // @[Interconnect.scala 146:19]
  wire  CCU_L2_WREADY; // @[Interconnect.scala 146:19]
  wire [63:0] CCU_L2_WDATA; // @[Interconnect.scala 146:19]
  wire  CCU_L2_WLAST; // @[Interconnect.scala 146:19]
  wire  CCU_L2_RVALID; // @[Interconnect.scala 146:19]
  wire  CCU_L2_RREADY; // @[Interconnect.scala 146:19]
  wire [63:0] CCU_L2_RDATA; // @[Interconnect.scala 146:19]
  wire [1:0] CCU_L2_RRESP; // @[Interconnect.scala 146:19]
  wire  CCU_L2_RLAST; // @[Interconnect.scala 146:19]
  wire  CCU_L2_BVALID; // @[Interconnect.scala 146:19]
  wire  CCU_L2_BREADY; // @[Interconnect.scala 146:19]
  wire [1:0] CCU_L2_BID; // @[Interconnect.scala 146:19]
  wire [1:0] CCU_L2_BRESP; // @[Interconnect.scala 146:19]
  wire  CCU_core0_ACVALID; // @[Interconnect.scala 146:19]
  wire  CCU_core0_ACREADY; // @[Interconnect.scala 146:19]
  wire [63:0] CCU_core0_ACADDR; // @[Interconnect.scala 146:19]
  wire [3:0] CCU_core0_ACSNOOP; // @[Interconnect.scala 146:19]
  wire  CCU_core0_CRVALID; // @[Interconnect.scala 146:19]
  wire  CCU_core0_CRREADY; // @[Interconnect.scala 146:19]
  wire [4:0] CCU_core0_CRRESP; // @[Interconnect.scala 146:19]
  wire  CCU_core0_CDVALID; // @[Interconnect.scala 146:19]
  wire  CCU_core0_CDREADY; // @[Interconnect.scala 146:19]
  wire [63:0] CCU_core0_CDDATA; // @[Interconnect.scala 146:19]
  wire  CCU_core0_CDLAST; // @[Interconnect.scala 146:19]
  wire  CCU_core0_RVALID; // @[Interconnect.scala 146:19]
  wire  CCU_core0_RREADY; // @[Interconnect.scala 146:19]
  wire [63:0] CCU_core0_RDATA; // @[Interconnect.scala 146:19]
  wire [3:0] CCU_core0_RRESP; // @[Interconnect.scala 146:19]
  wire  CCU_core0_RLAST; // @[Interconnect.scala 146:19]
  wire  CCU_core0_BVALID; // @[Interconnect.scala 146:19]
  wire  CCU_core0_BREADY; // @[Interconnect.scala 146:19]
  wire [1:0] CCU_core0_BRESP; // @[Interconnect.scala 146:19]
  wire  CCU_core1_RVALID; // @[Interconnect.scala 146:19]
  wire  CCU_core1_RREADY; // @[Interconnect.scala 146:19]
  wire [63:0] CCU_core1_RDATA; // @[Interconnect.scala 146:19]
  wire  CCU_core1_RLAST; // @[Interconnect.scala 146:19]
  wire  CCU_core1_BVALID; // @[Interconnect.scala 146:19]
  wire  CCU_core1_BREADY; // @[Interconnect.scala 146:19]
  wire [69:0] _FIFO_io_enq_bits_T_2 = {2'h0,io_acePort0_ARADDR,io_acePort0_ARSNOOP}; // @[Cat.scala 33:92]
  wire [69:0] _FIFO_io_enq_bits_T_4 = {2'h0,io_acePort0_AWADDR,1'h0,io_acePort0_AWSNOOP}; // @[Cat.scala 33:92]
  wire [69:0] _FIFO_io_enq_bits_T_5 = {2'h0,io_acePort0_WDATA,3'h0,io_acePort0_WLAST}; // @[Cat.scala 33:92]
  wire [69:0] _FIFO_io_enq_bits_T_8 = {2'h1,io_acePort1_ARADDR,4'h1}; // @[Cat.scala 33:92]
  wire [69:0] _GEN_1 = Arbiter_io_select == 3'h5 ? 70'h100000000000000000 : 70'h0; // @[Interconnect.scala 137:45 138:22]
  wire [69:0] _GEN_2 = Arbiter_io_select == 3'h4 ? _FIFO_io_enq_bits_T_8 : _GEN_1; // @[Interconnect.scala 135:45 136:22]
  wire [69:0] _GEN_3 = Arbiter_io_select == 3'h2 ? _FIFO_io_enq_bits_T_5 : _GEN_2; // @[Interconnect.scala 133:45 134:22]
  wire [69:0] _GEN_4 = Arbiter_io_select == 3'h1 ? _FIFO_io_enq_bits_T_4 : _GEN_3; // @[Interconnect.scala 131:45 132:22]
  arbiter_1 Arbiter ( // @[Interconnect.scala 88:23]
    .clock(Arbiter_clock),
    .reset(Arbiter_reset),
    .io_AWVALID_0(Arbiter_io_AWVALID_0),
    .io_AWREADY_0(Arbiter_io_AWREADY_0),
    .io_WVALID_0(Arbiter_io_WVALID_0),
    .io_WLAST_0(Arbiter_io_WLAST_0),
    .io_WREADY_0(Arbiter_io_WREADY_0),
    .io_ARVALID_0(Arbiter_io_ARVALID_0),
    .io_ARREADY_0(Arbiter_io_ARREADY_0),
    .io_ARVALID_1(Arbiter_io_ARVALID_1),
    .io_ARREADY_1(Arbiter_io_ARREADY_1),
    .io_select(Arbiter_io_select),
    .io_enq_valid(Arbiter_io_enq_valid),
    .io_enq_ready(Arbiter_io_enq_ready),
    .io_nstall(Arbiter_io_nstall)
  );
  ringbuffer FIFO ( // @[Interconnect.scala 112:20]
    .clock(FIFO_clock),
    .reset(FIFO_reset),
    .io_enq_ready(FIFO_io_enq_ready),
    .io_enq_valid(FIFO_io_enq_valid),
    .io_enq_bits(FIFO_io_enq_bits),
    .io_deq_ready(FIFO_io_deq_ready),
    .io_deq_valid(FIFO_io_deq_valid),
    .io_deq_bits(FIFO_io_deq_bits)
  );
  ccu CCU ( // @[Interconnect.scala 146:19]
    .clock(CCU_clock),
    .reset(CCU_reset),
    .deq_ready(CCU_deq_ready),
    .deq_valid(CCU_deq_valid),
    .deq_data(CCU_deq_data),
    .L2_AWVALID(CCU_L2_AWVALID),
    .L2_AWREADY(CCU_L2_AWREADY),
    .L2_AWID(CCU_L2_AWID),
    .L2_AWADDR(CCU_L2_AWADDR),
    .L2_ARVALID(CCU_L2_ARVALID),
    .L2_ARREADY(CCU_L2_ARREADY),
    .L2_ARID(CCU_L2_ARID),
    .L2_ARADDR(CCU_L2_ARADDR),
    .L2_WVALID(CCU_L2_WVALID),
    .L2_WREADY(CCU_L2_WREADY),
    .L2_WDATA(CCU_L2_WDATA),
    .L2_WLAST(CCU_L2_WLAST),
    .L2_RVALID(CCU_L2_RVALID),
    .L2_RREADY(CCU_L2_RREADY),
    .L2_RDATA(CCU_L2_RDATA),
    .L2_RRESP(CCU_L2_RRESP),
    .L2_RLAST(CCU_L2_RLAST),
    .L2_BVALID(CCU_L2_BVALID),
    .L2_BREADY(CCU_L2_BREADY),
    .L2_BID(CCU_L2_BID),
    .L2_BRESP(CCU_L2_BRESP),
    .core0_ACVALID(CCU_core0_ACVALID),
    .core0_ACREADY(CCU_core0_ACREADY),
    .core0_ACADDR(CCU_core0_ACADDR),
    .core0_ACSNOOP(CCU_core0_ACSNOOP),
    .core0_CRVALID(CCU_core0_CRVALID),
    .core0_CRREADY(CCU_core0_CRREADY),
    .core0_CRRESP(CCU_core0_CRRESP),
    .core0_CDVALID(CCU_core0_CDVALID),
    .core0_CDREADY(CCU_core0_CDREADY),
    .core0_CDDATA(CCU_core0_CDDATA),
    .core0_CDLAST(CCU_core0_CDLAST),
    .core0_RVALID(CCU_core0_RVALID),
    .core0_RREADY(CCU_core0_RREADY),
    .core0_RDATA(CCU_core0_RDATA),
    .core0_RRESP(CCU_core0_RRESP),
    .core0_RLAST(CCU_core0_RLAST),
    .core0_BVALID(CCU_core0_BVALID),
    .core0_BREADY(CCU_core0_BREADY),
    .core0_BRESP(CCU_core0_BRESP),
    .core1_RVALID(CCU_core1_RVALID),
    .core1_RREADY(CCU_core1_RREADY),
    .core1_RDATA(CCU_core1_RDATA),
    .core1_RLAST(CCU_core1_RLAST),
    .core1_BVALID(CCU_core1_BVALID),
    .core1_BREADY(CCU_core1_BREADY)
  );
  assign io_acePort0_AWREADY = Arbiter_io_AWREADY_0; // @[Interconnect.scala 93:23]
  assign io_acePort0_WREADY = Arbiter_io_WREADY_0; // @[Interconnect.scala 96:22]
  assign io_acePort0_BVALID = CCU_core0_BVALID; // @[Interconnect.scala 213:22]
  assign io_acePort0_BRESP = CCU_core0_BRESP; // @[Interconnect.scala 216:21]
  assign io_acePort0_ARREADY = Arbiter_io_ARREADY_0; // @[Interconnect.scala 98:23]
  assign io_acePort0_RVALID = CCU_core0_RVALID; // @[Interconnect.scala 205:22]
  assign io_acePort0_RDATA = CCU_core0_RDATA; // @[Interconnect.scala 209:21]
  assign io_acePort0_RRESP = CCU_core0_RRESP; // @[Interconnect.scala 208:21]
  assign io_acePort0_RLAST = CCU_core0_RLAST; // @[Interconnect.scala 210:21]
  assign io_acePort0_ACVALID = CCU_core0_ACVALID; // @[Interconnect.scala 188:23]
  assign io_acePort0_ACADDR = CCU_core0_ACADDR; // @[Interconnect.scala 190:22]
  assign io_acePort0_ACSNOOP = CCU_core0_ACSNOOP; // @[Interconnect.scala 191:23]
  assign io_acePort0_CRREADY = CCU_core0_CRREADY; // @[Interconnect.scala 195:23]
  assign io_acePort0_CDREADY = CCU_core0_CDREADY; // @[Interconnect.scala 200:23]
  assign io_acePort1_ARREADY = Arbiter_io_ARREADY_1; // @[Interconnect.scala 106:23]
  assign io_acePort1_RVALID = CCU_core1_RVALID; // @[Interconnect.scala 237:22]
  assign io_acePort1_RDATA = CCU_core1_RDATA; // @[Interconnect.scala 241:21]
  assign io_acePort1_RLAST = CCU_core1_RLAST; // @[Interconnect.scala 242:21]
  assign io_L2_AWVALID = CCU_L2_AWVALID; // @[Interconnect.scala 155:17]
  assign io_L2_AWID = CCU_L2_AWID; // @[Interconnect.scala 157:14]
  assign io_L2_AWADDR = CCU_L2_AWADDR; // @[Interconnect.scala 158:16]
  assign io_L2_ARVALID = CCU_L2_ARVALID; // @[Interconnect.scala 173:17]
  assign io_L2_ARID = CCU_L2_ARID; // @[Interconnect.scala 175:14]
  assign io_L2_ARADDR = CCU_L2_ARADDR; // @[Interconnect.scala 176:16]
  assign io_L2_WVALID = CCU_L2_WVALID; // @[Interconnect.scala 161:16]
  assign io_L2_WDATA = CCU_L2_WDATA; // @[Interconnect.scala 163:15]
  assign io_L2_WLAST = CCU_L2_WLAST; // @[Interconnect.scala 164:15]
  assign io_L2_RREADY = CCU_L2_RREADY; // @[Interconnect.scala 180:16]
  assign io_L2_BREADY = CCU_L2_BREADY; // @[Interconnect.scala 168:16]
  assign Arbiter_clock = clock;
  assign Arbiter_reset = reset;
  assign Arbiter_io_AWVALID_0 = io_acePort0_AWVALID; // @[Interconnect.scala 91:24]
  assign Arbiter_io_WVALID_0 = io_acePort0_WVALID; // @[Interconnect.scala 94:23]
  assign Arbiter_io_WLAST_0 = io_acePort0_WLAST; // @[Interconnect.scala 95:22]
  assign Arbiter_io_ARVALID_0 = io_acePort0_ARVALID; // @[Interconnect.scala 97:24]
  assign Arbiter_io_ARVALID_1 = io_acePort1_ARVALID; // @[Interconnect.scala 105:24]
  assign Arbiter_io_enq_ready = FIFO_io_enq_ready; // @[Interconnect.scala 116:24]
  assign Arbiter_io_nstall = CCU_core0_BVALID & CCU_core0_BREADY | CCU_core1_BVALID & CCU_core1_BREADY |
    CCU_core0_RVALID & CCU_core0_RREADY & CCU_core0_RLAST | CCU_core1_RVALID & CCU_core1_RREADY & CCU_core1_RLAST; // @[Interconnect.scala 250:166]
  assign FIFO_clock = clock;
  assign FIFO_reset = reset;
  assign FIFO_io_enq_valid = Arbiter_io_enq_valid; // @[Interconnect.scala 115:21]
  assign FIFO_io_enq_bits = Arbiter_io_select == 3'h0 ? _FIFO_io_enq_bits_T_2 : _GEN_4; // @[Interconnect.scala 129:39 130:22]
  assign FIFO_io_deq_ready = CCU_deq_ready; // @[Interconnect.scala 151:21]
  assign CCU_clock = clock;
  assign CCU_reset = reset;
  assign CCU_deq_valid = FIFO_io_deq_valid; // @[Interconnect.scala 149:17]
  assign CCU_deq_data = FIFO_io_deq_bits; // @[Interconnect.scala 150:16]
  assign CCU_L2_AWREADY = io_L2_AWREADY; // @[Interconnect.scala 156:18]
  assign CCU_L2_ARREADY = io_L2_ARREADY; // @[Interconnect.scala 174:18]
  assign CCU_L2_WREADY = io_L2_WREADY; // @[Interconnect.scala 162:17]
  assign CCU_L2_RVALID = io_L2_RVALID; // @[Interconnect.scala 179:17]
  assign CCU_L2_RDATA = io_L2_RDATA; // @[Interconnect.scala 183:16]
  assign CCU_L2_RRESP = io_L2_RRESP; // @[Interconnect.scala 182:16]
  assign CCU_L2_RLAST = io_L2_RLAST; // @[Interconnect.scala 184:16]
  assign CCU_L2_BVALID = io_L2_BVALID; // @[Interconnect.scala 167:17]
  assign CCU_L2_BID = io_L2_BID; // @[Interconnect.scala 169:14]
  assign CCU_L2_BRESP = io_L2_BRESP; // @[Interconnect.scala 170:16]
  assign CCU_core0_ACREADY = io_acePort0_ACREADY; // @[Interconnect.scala 189:21]
  assign CCU_core0_CRVALID = io_acePort0_CRVALID; // @[Interconnect.scala 194:21]
  assign CCU_core0_CRRESP = io_acePort0_CRRESP; // @[Interconnect.scala 196:20]
  assign CCU_core0_CDVALID = io_acePort0_CDVALID; // @[Interconnect.scala 199:21]
  assign CCU_core0_CDDATA = io_acePort0_CDDATA; // @[Interconnect.scala 201:20]
  assign CCU_core0_CDLAST = io_acePort0_CDLAST; // @[Interconnect.scala 202:20]
  assign CCU_core0_RREADY = io_acePort0_RREADY; // @[Interconnect.scala 206:20]
  assign CCU_core0_BREADY = io_acePort0_BREADY; // @[Interconnect.scala 214:20]
  assign CCU_core1_RREADY = io_acePort1_RREADY; // @[Interconnect.scala 238:20]
  assign CCU_core1_BREADY = 1'h0; // @[Interconnect.scala 246:20]
endmodule
module soc1(
  input         clock,
  input         reset,
  output        L2_AWVALID,
  input         L2_AWREADY,
  output [1:0]  L2_AWID,
  output [63:0] L2_AWADDR,
  output [7:0]  L2_AWLEN,
  output [2:0]  L2_AWSIZE,
  output [1:0]  L2_AWBURST,
  output        L2_AWLOCK,
  output [3:0]  L2_AWCACHE,
  output [2:0]  L2_AWPROT,
  output [3:0]  L2_AWQOS,
  output        L2_ARVALID,
  input         L2_ARREADY,
  output [1:0]  L2_ARID,
  output [63:0] L2_ARADDR,
  output [7:0]  L2_ARLEN,
  output [2:0]  L2_ARSIZE,
  output [1:0]  L2_ARBURST,
  output        L2_ARLOCK,
  output [3:0]  L2_ARCACHE,
  output [2:0]  L2_ARPROT,
  output [3:0]  L2_ARQOS,
  output        L2_WVALID,
  input         L2_WREADY,
  output [63:0] L2_WDATA,
  output [7:0]  L2_WSTRB,
  output        L2_WLAST,
  input         L2_RVALID,
  output        L2_RREADY,
  input  [1:0]  L2_RID,
  input  [63:0] L2_RDATA,
  input  [1:0]  L2_RRESP,
  input         L2_RLAST,
  input         L2_BVALID,
  output        L2_BREADY,
  input  [1:0]  L2_BID,
  input  [1:0]  L2_BRESP,
  input         MTIP,
  output        core_sample0,
  output        core_sample1,
  output        peripheral_AWID,
  output [31:0] peripheral_AWADDR,
  output [7:0]  peripheral_AWLEN,
  output [2:0]  peripheral_AWSIZE,
  output [1:0]  peripheral_AWBURST,
  output        peripheral_AWLOCK,
  output [3:0]  peripheral_AWCACHE,
  output [2:0]  peripheral_AWPROT,
  output [3:0]  peripheral_AWQOS,
  output        peripheral_AWVALID,
  input         peripheral_AWREADY,
  output [31:0] peripheral_WDATA,
  output [3:0]  peripheral_WSTRB,
  output        peripheral_WLAST,
  output        peripheral_WVALID,
  input         peripheral_WREADY,
  input         peripheral_BID,
  input  [1:0]  peripheral_BRESP,
  input         peripheral_BVALID,
  output        peripheral_BREADY,
  output        peripheral_ARID,
  output [31:0] peripheral_ARADDR,
  output [7:0]  peripheral_ARLEN,
  output [2:0]  peripheral_ARSIZE,
  output [1:0]  peripheral_ARBURST,
  output        peripheral_ARLOCK,
  output [3:0]  peripheral_ARCACHE,
  output [2:0]  peripheral_ARPROT,
  output [3:0]  peripheral_ARQOS,
  output        peripheral_ARVALID,
  input         peripheral_ARREADY,
  input         peripheral_RID,
  input  [31:0] peripheral_RDATA,
  input  [1:0]  peripheral_RRESP,
  input         peripheral_RLAST,
  input         peripheral_RVALID,
  output        peripheral_RREADY,
  output        debug_probe_arvalid_internal,
  output        debug_probe_cacheMissed,
  output        debug_probe_rready_signal,
  output        debug_probe_cacheFill_valid,
  output        debug_probe_axi_arvalid,
  output        debug_probe_axi_arready,
  output        debug_probe_req_valid,
  output [63:0] debug_probe_req_pc,
  output        fdbg_probe_redirect_bit,
  output        fdbg_probe_fifo_enq_ready,
  output        fdbg_probe_is_fence,
  output        fdbg_probe_handle_fence
);
  wire  core0_clock; // @[soc.scala 89:21]
  wire  core0_reset; // @[soc.scala 89:21]
  wire [31:0] core0_iPort_ARADDR; // @[soc.scala 89:21]
  wire  core0_iPort_ARVALID; // @[soc.scala 89:21]
  wire  core0_iPort_ARREADY; // @[soc.scala 89:21]
  wire [63:0] core0_iPort_RDATA; // @[soc.scala 89:21]
  wire  core0_iPort_RLAST; // @[soc.scala 89:21]
  wire  core0_iPort_RVALID; // @[soc.scala 89:21]
  wire  core0_iPort_RREADY; // @[soc.scala 89:21]
  wire  core0_debug_probe_arvalid_internal; // @[soc.scala 89:21]
  wire  core0_debug_probe_cacheMissed; // @[soc.scala 89:21]
  wire  core0_debug_probe_rready_signal; // @[soc.scala 89:21]
  wire  core0_debug_probe_cacheFill_valid; // @[soc.scala 89:21]
  wire  core0_debug_probe_axi_arvalid; // @[soc.scala 89:21]
  wire  core0_debug_probe_axi_arready; // @[soc.scala 89:21]
  wire  core0_debug_probe_req_valid; // @[soc.scala 89:21]
  wire [63:0] core0_debug_probe_req_pc; // @[soc.scala 89:21]
  wire  core0_fdbg_probe_redirect_bit; // @[soc.scala 89:21]
  wire  core0_fdbg_probe_fifo_enq_ready; // @[soc.scala 89:21]
  wire  core0_fdbg_probe_is_fence; // @[soc.scala 89:21]
  wire  core0_fdbg_probe_handle_fence; // @[soc.scala 89:21]
  wire [31:0] core0_dPort_AWADDR; // @[soc.scala 89:21]
  wire  core0_dPort_AWVALID; // @[soc.scala 89:21]
  wire  core0_dPort_AWREADY; // @[soc.scala 89:21]
  wire [63:0] core0_dPort_WDATA; // @[soc.scala 89:21]
  wire  core0_dPort_WLAST; // @[soc.scala 89:21]
  wire  core0_dPort_WVALID; // @[soc.scala 89:21]
  wire  core0_dPort_WREADY; // @[soc.scala 89:21]
  wire [1:0] core0_dPort_BRESP; // @[soc.scala 89:21]
  wire  core0_dPort_BVALID; // @[soc.scala 89:21]
  wire  core0_dPort_BREADY; // @[soc.scala 89:21]
  wire [31:0] core0_dPort_ARADDR; // @[soc.scala 89:21]
  wire  core0_dPort_ARVALID; // @[soc.scala 89:21]
  wire  core0_dPort_ARREADY; // @[soc.scala 89:21]
  wire [63:0] core0_dPort_RDATA; // @[soc.scala 89:21]
  wire  core0_dPort_RLAST; // @[soc.scala 89:21]
  wire  core0_dPort_RVALID; // @[soc.scala 89:21]
  wire  core0_dPort_RREADY; // @[soc.scala 89:21]
  wire [2:0] core0_dPort_AWSNOOP; // @[soc.scala 89:21]
  wire [3:0] core0_dPort_ARSNOOP; // @[soc.scala 89:21]
  wire [3:0] core0_dPort_RRESP; // @[soc.scala 89:21]
  wire  core0_dPort_ACVALID; // @[soc.scala 89:21]
  wire  core0_dPort_ACREADY; // @[soc.scala 89:21]
  wire [31:0] core0_dPort_ACADDR; // @[soc.scala 89:21]
  wire [3:0] core0_dPort_ACSNOOP; // @[soc.scala 89:21]
  wire  core0_dPort_CRVALID; // @[soc.scala 89:21]
  wire  core0_dPort_CRREADY; // @[soc.scala 89:21]
  wire [4:0] core0_dPort_CRRESP; // @[soc.scala 89:21]
  wire  core0_dPort_CDVALID; // @[soc.scala 89:21]
  wire  core0_dPort_CDREADY; // @[soc.scala 89:21]
  wire [63:0] core0_dPort_CDDATA; // @[soc.scala 89:21]
  wire  core0_dPort_CDLAST; // @[soc.scala 89:21]
  wire [31:0] core0_peripheral_AWADDR; // @[soc.scala 89:21]
  wire [7:0] core0_peripheral_AWLEN; // @[soc.scala 89:21]
  wire [2:0] core0_peripheral_AWSIZE; // @[soc.scala 89:21]
  wire [1:0] core0_peripheral_AWBURST; // @[soc.scala 89:21]
  wire [2:0] core0_peripheral_AWPROT; // @[soc.scala 89:21]
  wire  core0_peripheral_AWVALID; // @[soc.scala 89:21]
  wire  core0_peripheral_AWREADY; // @[soc.scala 89:21]
  wire [31:0] core0_peripheral_WDATA; // @[soc.scala 89:21]
  wire [3:0] core0_peripheral_WSTRB; // @[soc.scala 89:21]
  wire  core0_peripheral_WLAST; // @[soc.scala 89:21]
  wire  core0_peripheral_WVALID; // @[soc.scala 89:21]
  wire  core0_peripheral_WREADY; // @[soc.scala 89:21]
  wire  core0_peripheral_BID; // @[soc.scala 89:21]
  wire [1:0] core0_peripheral_BRESP; // @[soc.scala 89:21]
  wire  core0_peripheral_BVALID; // @[soc.scala 89:21]
  wire  core0_peripheral_BREADY; // @[soc.scala 89:21]
  wire [31:0] core0_peripheral_ARADDR; // @[soc.scala 89:21]
  wire [7:0] core0_peripheral_ARLEN; // @[soc.scala 89:21]
  wire [2:0] core0_peripheral_ARSIZE; // @[soc.scala 89:21]
  wire [1:0] core0_peripheral_ARBURST; // @[soc.scala 89:21]
  wire [2:0] core0_peripheral_ARPROT; // @[soc.scala 89:21]
  wire  core0_peripheral_ARVALID; // @[soc.scala 89:21]
  wire  core0_peripheral_ARREADY; // @[soc.scala 89:21]
  wire  core0_peripheral_RID; // @[soc.scala 89:21]
  wire [31:0] core0_peripheral_RDATA; // @[soc.scala 89:21]
  wire [1:0] core0_peripheral_RRESP; // @[soc.scala 89:21]
  wire  core0_peripheral_RLAST; // @[soc.scala 89:21]
  wire  core0_peripheral_RVALID; // @[soc.scala 89:21]
  wire  core0_peripheral_RREADY; // @[soc.scala 89:21]
  wire  core0_core_sample0; // @[soc.scala 89:21]
  wire  core0_core_sample1; // @[soc.scala 89:21]
  wire  core0_MTIP; // @[soc.scala 89:21]
  wire  interconnect__clock; // @[soc.scala 115:28]
  wire  interconnect__reset; // @[soc.scala 115:28]
  wire  interconnect__io_acePort0_AWVALID; // @[soc.scala 115:28]
  wire  interconnect__io_acePort0_AWREADY; // @[soc.scala 115:28]
  wire [63:0] interconnect__io_acePort0_AWADDR; // @[soc.scala 115:28]
  wire [2:0] interconnect__io_acePort0_AWSNOOP; // @[soc.scala 115:28]
  wire  interconnect__io_acePort0_WVALID; // @[soc.scala 115:28]
  wire  interconnect__io_acePort0_WREADY; // @[soc.scala 115:28]
  wire [63:0] interconnect__io_acePort0_WDATA; // @[soc.scala 115:28]
  wire  interconnect__io_acePort0_WLAST; // @[soc.scala 115:28]
  wire  interconnect__io_acePort0_BVALID; // @[soc.scala 115:28]
  wire  interconnect__io_acePort0_BREADY; // @[soc.scala 115:28]
  wire [1:0] interconnect__io_acePort0_BRESP; // @[soc.scala 115:28]
  wire  interconnect__io_acePort0_ARVALID; // @[soc.scala 115:28]
  wire  interconnect__io_acePort0_ARREADY; // @[soc.scala 115:28]
  wire [63:0] interconnect__io_acePort0_ARADDR; // @[soc.scala 115:28]
  wire [3:0] interconnect__io_acePort0_ARSNOOP; // @[soc.scala 115:28]
  wire  interconnect__io_acePort0_RVALID; // @[soc.scala 115:28]
  wire  interconnect__io_acePort0_RREADY; // @[soc.scala 115:28]
  wire [63:0] interconnect__io_acePort0_RDATA; // @[soc.scala 115:28]
  wire [3:0] interconnect__io_acePort0_RRESP; // @[soc.scala 115:28]
  wire  interconnect__io_acePort0_RLAST; // @[soc.scala 115:28]
  wire  interconnect__io_acePort0_ACVALID; // @[soc.scala 115:28]
  wire  interconnect__io_acePort0_ACREADY; // @[soc.scala 115:28]
  wire [63:0] interconnect__io_acePort0_ACADDR; // @[soc.scala 115:28]
  wire [3:0] interconnect__io_acePort0_ACSNOOP; // @[soc.scala 115:28]
  wire  interconnect__io_acePort0_CRVALID; // @[soc.scala 115:28]
  wire  interconnect__io_acePort0_CRREADY; // @[soc.scala 115:28]
  wire [4:0] interconnect__io_acePort0_CRRESP; // @[soc.scala 115:28]
  wire  interconnect__io_acePort0_CDVALID; // @[soc.scala 115:28]
  wire  interconnect__io_acePort0_CDREADY; // @[soc.scala 115:28]
  wire [63:0] interconnect__io_acePort0_CDDATA; // @[soc.scala 115:28]
  wire  interconnect__io_acePort0_CDLAST; // @[soc.scala 115:28]
  wire  interconnect__io_acePort1_ARVALID; // @[soc.scala 115:28]
  wire  interconnect__io_acePort1_ARREADY; // @[soc.scala 115:28]
  wire [63:0] interconnect__io_acePort1_ARADDR; // @[soc.scala 115:28]
  wire  interconnect__io_acePort1_RVALID; // @[soc.scala 115:28]
  wire  interconnect__io_acePort1_RREADY; // @[soc.scala 115:28]
  wire [63:0] interconnect__io_acePort1_RDATA; // @[soc.scala 115:28]
  wire  interconnect__io_acePort1_RLAST; // @[soc.scala 115:28]
  wire  interconnect__io_L2_AWVALID; // @[soc.scala 115:28]
  wire  interconnect__io_L2_AWREADY; // @[soc.scala 115:28]
  wire [1:0] interconnect__io_L2_AWID; // @[soc.scala 115:28]
  wire [63:0] interconnect__io_L2_AWADDR; // @[soc.scala 115:28]
  wire  interconnect__io_L2_ARVALID; // @[soc.scala 115:28]
  wire  interconnect__io_L2_ARREADY; // @[soc.scala 115:28]
  wire [1:0] interconnect__io_L2_ARID; // @[soc.scala 115:28]
  wire [63:0] interconnect__io_L2_ARADDR; // @[soc.scala 115:28]
  wire  interconnect__io_L2_WVALID; // @[soc.scala 115:28]
  wire  interconnect__io_L2_WREADY; // @[soc.scala 115:28]
  wire [63:0] interconnect__io_L2_WDATA; // @[soc.scala 115:28]
  wire  interconnect__io_L2_WLAST; // @[soc.scala 115:28]
  wire  interconnect__io_L2_RVALID; // @[soc.scala 115:28]
  wire  interconnect__io_L2_RREADY; // @[soc.scala 115:28]
  wire [63:0] interconnect__io_L2_RDATA; // @[soc.scala 115:28]
  wire [1:0] interconnect__io_L2_RRESP; // @[soc.scala 115:28]
  wire  interconnect__io_L2_RLAST; // @[soc.scala 115:28]
  wire  interconnect__io_L2_BVALID; // @[soc.scala 115:28]
  wire  interconnect__io_L2_BREADY; // @[soc.scala 115:28]
  wire [1:0] interconnect__io_L2_BID; // @[soc.scala 115:28]
  wire [1:0] interconnect__io_L2_BRESP; // @[soc.scala 115:28]
  soc1_Anon core0 ( // @[soc.scala 89:21]
    .clock(core0_clock),
    .reset(core0_reset),
    .iPort_ARADDR(core0_iPort_ARADDR),
    .iPort_ARVALID(core0_iPort_ARVALID),
    .iPort_ARREADY(core0_iPort_ARREADY),
    .iPort_RDATA(core0_iPort_RDATA),
    .iPort_RLAST(core0_iPort_RLAST),
    .iPort_RVALID(core0_iPort_RVALID),
    .iPort_RREADY(core0_iPort_RREADY),
    .debug_probe_arvalid_internal(core0_debug_probe_arvalid_internal),
    .debug_probe_cacheMissed(core0_debug_probe_cacheMissed),
    .debug_probe_rready_signal(core0_debug_probe_rready_signal),
    .debug_probe_cacheFill_valid(core0_debug_probe_cacheFill_valid),
    .debug_probe_axi_arvalid(core0_debug_probe_axi_arvalid),
    .debug_probe_axi_arready(core0_debug_probe_axi_arready),
    .debug_probe_req_valid(core0_debug_probe_req_valid),
    .debug_probe_req_pc(core0_debug_probe_req_pc),
    .fdbg_probe_redirect_bit(core0_fdbg_probe_redirect_bit),
    .fdbg_probe_fifo_enq_ready(core0_fdbg_probe_fifo_enq_ready),
    .fdbg_probe_is_fence(core0_fdbg_probe_is_fence),
    .fdbg_probe_handle_fence(core0_fdbg_probe_handle_fence),
    .dPort_AWADDR(core0_dPort_AWADDR),
    .dPort_AWVALID(core0_dPort_AWVALID),
    .dPort_AWREADY(core0_dPort_AWREADY),
    .dPort_WDATA(core0_dPort_WDATA),
    .dPort_WLAST(core0_dPort_WLAST),
    .dPort_WVALID(core0_dPort_WVALID),
    .dPort_WREADY(core0_dPort_WREADY),
    .dPort_BRESP(core0_dPort_BRESP),
    .dPort_BVALID(core0_dPort_BVALID),
    .dPort_BREADY(core0_dPort_BREADY),
    .dPort_ARADDR(core0_dPort_ARADDR),
    .dPort_ARVALID(core0_dPort_ARVALID),
    .dPort_ARREADY(core0_dPort_ARREADY),
    .dPort_RDATA(core0_dPort_RDATA),
    .dPort_RLAST(core0_dPort_RLAST),
    .dPort_RVALID(core0_dPort_RVALID),
    .dPort_RREADY(core0_dPort_RREADY),
    .dPort_AWSNOOP(core0_dPort_AWSNOOP),
    .dPort_ARSNOOP(core0_dPort_ARSNOOP),
    .dPort_RRESP(core0_dPort_RRESP),
    .dPort_ACVALID(core0_dPort_ACVALID),
    .dPort_ACREADY(core0_dPort_ACREADY),
    .dPort_ACADDR(core0_dPort_ACADDR),
    .dPort_ACSNOOP(core0_dPort_ACSNOOP),
    .dPort_CRVALID(core0_dPort_CRVALID),
    .dPort_CRREADY(core0_dPort_CRREADY),
    .dPort_CRRESP(core0_dPort_CRRESP),
    .dPort_CDVALID(core0_dPort_CDVALID),
    .dPort_CDREADY(core0_dPort_CDREADY),
    .dPort_CDDATA(core0_dPort_CDDATA),
    .dPort_CDLAST(core0_dPort_CDLAST),
    .peripheral_AWADDR(core0_peripheral_AWADDR),
    .peripheral_AWLEN(core0_peripheral_AWLEN),
    .peripheral_AWSIZE(core0_peripheral_AWSIZE),
    .peripheral_AWBURST(core0_peripheral_AWBURST),
    .peripheral_AWPROT(core0_peripheral_AWPROT),
    .peripheral_AWVALID(core0_peripheral_AWVALID),
    .peripheral_AWREADY(core0_peripheral_AWREADY),
    .peripheral_WDATA(core0_peripheral_WDATA),
    .peripheral_WSTRB(core0_peripheral_WSTRB),
    .peripheral_WLAST(core0_peripheral_WLAST),
    .peripheral_WVALID(core0_peripheral_WVALID),
    .peripheral_WREADY(core0_peripheral_WREADY),
    .peripheral_BID(core0_peripheral_BID),
    .peripheral_BRESP(core0_peripheral_BRESP),
    .peripheral_BVALID(core0_peripheral_BVALID),
    .peripheral_BREADY(core0_peripheral_BREADY),
    .peripheral_ARADDR(core0_peripheral_ARADDR),
    .peripheral_ARLEN(core0_peripheral_ARLEN),
    .peripheral_ARSIZE(core0_peripheral_ARSIZE),
    .peripheral_ARBURST(core0_peripheral_ARBURST),
    .peripheral_ARPROT(core0_peripheral_ARPROT),
    .peripheral_ARVALID(core0_peripheral_ARVALID),
    .peripheral_ARREADY(core0_peripheral_ARREADY),
    .peripheral_RID(core0_peripheral_RID),
    .peripheral_RDATA(core0_peripheral_RDATA),
    .peripheral_RRESP(core0_peripheral_RRESP),
    .peripheral_RLAST(core0_peripheral_RLAST),
    .peripheral_RVALID(core0_peripheral_RVALID),
    .peripheral_RREADY(core0_peripheral_RREADY),
    .core_sample0(core0_core_sample0),
    .core_sample1(core0_core_sample1),
    .MTIP(core0_MTIP)
  );
  Interconnect interconnect_ ( // @[soc.scala 115:28]
    .clock(interconnect__clock),
    .reset(interconnect__reset),
    .io_acePort0_AWVALID(interconnect__io_acePort0_AWVALID),
    .io_acePort0_AWREADY(interconnect__io_acePort0_AWREADY),
    .io_acePort0_AWADDR(interconnect__io_acePort0_AWADDR),
    .io_acePort0_AWSNOOP(interconnect__io_acePort0_AWSNOOP),
    .io_acePort0_WVALID(interconnect__io_acePort0_WVALID),
    .io_acePort0_WREADY(interconnect__io_acePort0_WREADY),
    .io_acePort0_WDATA(interconnect__io_acePort0_WDATA),
    .io_acePort0_WLAST(interconnect__io_acePort0_WLAST),
    .io_acePort0_BVALID(interconnect__io_acePort0_BVALID),
    .io_acePort0_BREADY(interconnect__io_acePort0_BREADY),
    .io_acePort0_BRESP(interconnect__io_acePort0_BRESP),
    .io_acePort0_ARVALID(interconnect__io_acePort0_ARVALID),
    .io_acePort0_ARREADY(interconnect__io_acePort0_ARREADY),
    .io_acePort0_ARADDR(interconnect__io_acePort0_ARADDR),
    .io_acePort0_ARSNOOP(interconnect__io_acePort0_ARSNOOP),
    .io_acePort0_RVALID(interconnect__io_acePort0_RVALID),
    .io_acePort0_RREADY(interconnect__io_acePort0_RREADY),
    .io_acePort0_RDATA(interconnect__io_acePort0_RDATA),
    .io_acePort0_RRESP(interconnect__io_acePort0_RRESP),
    .io_acePort0_RLAST(interconnect__io_acePort0_RLAST),
    .io_acePort0_ACVALID(interconnect__io_acePort0_ACVALID),
    .io_acePort0_ACREADY(interconnect__io_acePort0_ACREADY),
    .io_acePort0_ACADDR(interconnect__io_acePort0_ACADDR),
    .io_acePort0_ACSNOOP(interconnect__io_acePort0_ACSNOOP),
    .io_acePort0_CRVALID(interconnect__io_acePort0_CRVALID),
    .io_acePort0_CRREADY(interconnect__io_acePort0_CRREADY),
    .io_acePort0_CRRESP(interconnect__io_acePort0_CRRESP),
    .io_acePort0_CDVALID(interconnect__io_acePort0_CDVALID),
    .io_acePort0_CDREADY(interconnect__io_acePort0_CDREADY),
    .io_acePort0_CDDATA(interconnect__io_acePort0_CDDATA),
    .io_acePort0_CDLAST(interconnect__io_acePort0_CDLAST),
    .io_acePort1_ARVALID(interconnect__io_acePort1_ARVALID),
    .io_acePort1_ARREADY(interconnect__io_acePort1_ARREADY),
    .io_acePort1_ARADDR(interconnect__io_acePort1_ARADDR),
    .io_acePort1_RVALID(interconnect__io_acePort1_RVALID),
    .io_acePort1_RREADY(interconnect__io_acePort1_RREADY),
    .io_acePort1_RDATA(interconnect__io_acePort1_RDATA),
    .io_acePort1_RLAST(interconnect__io_acePort1_RLAST),
    .io_L2_AWVALID(interconnect__io_L2_AWVALID),
    .io_L2_AWREADY(interconnect__io_L2_AWREADY),
    .io_L2_AWID(interconnect__io_L2_AWID),
    .io_L2_AWADDR(interconnect__io_L2_AWADDR),
    .io_L2_ARVALID(interconnect__io_L2_ARVALID),
    .io_L2_ARREADY(interconnect__io_L2_ARREADY),
    .io_L2_ARID(interconnect__io_L2_ARID),
    .io_L2_ARADDR(interconnect__io_L2_ARADDR),
    .io_L2_WVALID(interconnect__io_L2_WVALID),
    .io_L2_WREADY(interconnect__io_L2_WREADY),
    .io_L2_WDATA(interconnect__io_L2_WDATA),
    .io_L2_WLAST(interconnect__io_L2_WLAST),
    .io_L2_RVALID(interconnect__io_L2_RVALID),
    .io_L2_RREADY(interconnect__io_L2_RREADY),
    .io_L2_RDATA(interconnect__io_L2_RDATA),
    .io_L2_RRESP(interconnect__io_L2_RRESP),
    .io_L2_RLAST(interconnect__io_L2_RLAST),
    .io_L2_BVALID(interconnect__io_L2_BVALID),
    .io_L2_BREADY(interconnect__io_L2_BREADY),
    .io_L2_BID(interconnect__io_L2_BID),
    .io_L2_BRESP(interconnect__io_L2_BRESP)
  );
  assign L2_AWVALID = interconnect__io_L2_AWVALID; // @[soc.scala 278:14]
  assign L2_AWID = interconnect__io_L2_AWID; // @[soc.scala 280:11]
  assign L2_AWADDR = interconnect__io_L2_AWADDR; // @[soc.scala 281:13]
  assign L2_AWLEN = 8'h7; // @[soc.scala 282:12]
  assign L2_AWSIZE = 3'h3; // @[soc.scala 283:13]
  assign L2_AWBURST = 2'h1; // @[soc.scala 284:14]
  assign L2_AWLOCK = 1'h0; // @[soc.scala 285:13]
  assign L2_AWCACHE = 4'h2; // @[soc.scala 286:14]
  assign L2_AWPROT = 3'h0; // @[soc.scala 287:13]
  assign L2_AWQOS = 4'h0; // @[soc.scala 288:12]
  assign L2_ARVALID = interconnect__io_L2_ARVALID; // @[soc.scala 291:14]
  assign L2_ARID = interconnect__io_L2_ARID; // @[soc.scala 293:11]
  assign L2_ARADDR = interconnect__io_L2_ARADDR; // @[soc.scala 294:13]
  assign L2_ARLEN = 8'h7; // @[soc.scala 295:12]
  assign L2_ARSIZE = 3'h3; // @[soc.scala 296:13]
  assign L2_ARBURST = 2'h1; // @[soc.scala 297:14]
  assign L2_ARLOCK = 1'h0; // @[soc.scala 298:13]
  assign L2_ARCACHE = 4'h2; // @[soc.scala 299:14]
  assign L2_ARPROT = 3'h0; // @[soc.scala 300:13]
  assign L2_ARQOS = 4'h0; // @[soc.scala 301:12]
  assign L2_WVALID = interconnect__io_L2_WVALID; // @[soc.scala 305:13]
  assign L2_WDATA = interconnect__io_L2_WDATA; // @[soc.scala 307:12]
  assign L2_WSTRB = 8'hff; // @[soc.scala 309:12]
  assign L2_WLAST = interconnect__io_L2_WLAST; // @[soc.scala 308:12]
  assign L2_RREADY = interconnect__io_L2_RREADY; // @[soc.scala 313:13]
  assign L2_BREADY = interconnect__io_L2_BREADY; // @[soc.scala 322:13]
  assign core_sample0 = core0_core_sample0; // @[soc.scala 118:16]
  assign core_sample1 = core0_core_sample1; // @[soc.scala 119:16]
  assign peripheral_AWID = 1'h0; // @[soc.scala 120:20]
  assign peripheral_AWADDR = core0_peripheral_AWADDR; // @[soc.scala 120:20]
  assign peripheral_AWLEN = core0_peripheral_AWLEN; // @[soc.scala 120:20]
  assign peripheral_AWSIZE = core0_peripheral_AWSIZE; // @[soc.scala 120:20]
  assign peripheral_AWBURST = core0_peripheral_AWBURST; // @[soc.scala 120:20]
  assign peripheral_AWLOCK = 1'h0; // @[soc.scala 120:20]
  assign peripheral_AWCACHE = 4'h0; // @[soc.scala 120:20]
  assign peripheral_AWPROT = core0_peripheral_AWPROT; // @[soc.scala 120:20]
  assign peripheral_AWQOS = 4'h0; // @[soc.scala 120:20]
  assign peripheral_AWVALID = core0_peripheral_AWVALID; // @[soc.scala 120:20]
  assign peripheral_WDATA = core0_peripheral_WDATA; // @[soc.scala 120:20]
  assign peripheral_WSTRB = core0_peripheral_WSTRB; // @[soc.scala 120:20]
  assign peripheral_WLAST = core0_peripheral_WLAST; // @[soc.scala 120:20]
  assign peripheral_WVALID = core0_peripheral_WVALID; // @[soc.scala 120:20]
  assign peripheral_BREADY = core0_peripheral_BREADY; // @[soc.scala 120:20]
  assign peripheral_ARID = 1'h0; // @[soc.scala 120:20]
  assign peripheral_ARADDR = core0_peripheral_ARADDR; // @[soc.scala 120:20]
  assign peripheral_ARLEN = core0_peripheral_ARLEN; // @[soc.scala 120:20]
  assign peripheral_ARSIZE = core0_peripheral_ARSIZE; // @[soc.scala 120:20]
  assign peripheral_ARBURST = core0_peripheral_ARBURST; // @[soc.scala 120:20]
  assign peripheral_ARLOCK = 1'h0; // @[soc.scala 120:20]
  assign peripheral_ARCACHE = 4'h0; // @[soc.scala 120:20]
  assign peripheral_ARPROT = core0_peripheral_ARPROT; // @[soc.scala 120:20]
  assign peripheral_ARQOS = 4'h0; // @[soc.scala 120:20]
  assign peripheral_ARVALID = core0_peripheral_ARVALID; // @[soc.scala 120:20]
  assign peripheral_RREADY = core0_peripheral_RREADY; // @[soc.scala 120:20]
  assign debug_probe_arvalid_internal = core0_debug_probe_arvalid_internal; // @[soc.scala 124:9]
  assign debug_probe_cacheMissed = core0_debug_probe_cacheMissed; // @[soc.scala 124:9]
  assign debug_probe_rready_signal = core0_debug_probe_rready_signal; // @[soc.scala 124:9]
  assign debug_probe_cacheFill_valid = core0_debug_probe_cacheFill_valid; // @[soc.scala 124:9]
  assign debug_probe_axi_arvalid = core0_debug_probe_axi_arvalid; // @[soc.scala 124:9]
  assign debug_probe_axi_arready = core0_debug_probe_axi_arready; // @[soc.scala 124:9]
  assign debug_probe_req_valid = core0_debug_probe_req_valid; // @[soc.scala 124:9]
  assign debug_probe_req_pc = core0_debug_probe_req_pc; // @[soc.scala 124:9]
  assign fdbg_probe_redirect_bit = core0_fdbg_probe_redirect_bit; // @[soc.scala 126:8]
  assign fdbg_probe_fifo_enq_ready = core0_fdbg_probe_fifo_enq_ready; // @[soc.scala 126:8]
  assign fdbg_probe_is_fence = core0_fdbg_probe_is_fence; // @[soc.scala 126:8]
  assign fdbg_probe_handle_fence = core0_fdbg_probe_handle_fence; // @[soc.scala 126:8]
  assign core0_clock = clock;
  assign core0_reset = reset;
  assign core0_iPort_ARREADY = interconnect__io_acePort1_ARREADY; // @[soc.scala 211:23]
  assign core0_iPort_RDATA = interconnect__io_acePort1_RDATA; // @[soc.scala 221:21]
  assign core0_iPort_RLAST = interconnect__io_acePort1_RLAST; // @[soc.scala 223:21]
  assign core0_iPort_RVALID = interconnect__io_acePort1_RVALID; // @[soc.scala 218:22]
  assign core0_dPort_AWREADY = interconnect__io_acePort0_AWREADY; // @[soc.scala 136:23]
  assign core0_dPort_WREADY = interconnect__io_acePort0_WREADY; // @[soc.scala 146:22]
  assign core0_dPort_BRESP = interconnect__io_acePort0_BRESP; // @[soc.scala 151:21]
  assign core0_dPort_BVALID = interconnect__io_acePort0_BVALID; // @[soc.scala 149:22]
  assign core0_dPort_ARREADY = interconnect__io_acePort0_ARREADY; // @[soc.scala 156:23]
  assign core0_dPort_RDATA = interconnect__io_acePort0_RDATA; // @[soc.scala 166:21]
  assign core0_dPort_RLAST = interconnect__io_acePort0_RLAST; // @[soc.scala 168:21]
  assign core0_dPort_RVALID = interconnect__io_acePort0_RVALID; // @[soc.scala 163:22]
  assign core0_dPort_RRESP = interconnect__io_acePort0_RRESP; // @[soc.scala 167:21]
  assign core0_dPort_ACVALID = interconnect__io_acePort0_ACVALID; // @[soc.scala 171:23]
  assign core0_dPort_ACADDR = interconnect__io_acePort0_ACADDR[31:0]; // @[soc.scala 172:22]
  assign core0_dPort_ACSNOOP = interconnect__io_acePort0_ACSNOOP; // @[soc.scala 173:23]
  assign core0_dPort_CRREADY = interconnect__io_acePort0_CRREADY; // @[soc.scala 180:23]
  assign core0_dPort_CDREADY = interconnect__io_acePort0_CDREADY; // @[soc.scala 184:23]
  assign core0_peripheral_AWREADY = peripheral_AWREADY; // @[soc.scala 120:20]
  assign core0_peripheral_WREADY = peripheral_WREADY; // @[soc.scala 120:20]
  assign core0_peripheral_BID = peripheral_BID; // @[soc.scala 120:20]
  assign core0_peripheral_BRESP = peripheral_BRESP; // @[soc.scala 120:20]
  assign core0_peripheral_BVALID = peripheral_BVALID; // @[soc.scala 120:20]
  assign core0_peripheral_ARREADY = peripheral_ARREADY; // @[soc.scala 120:20]
  assign core0_peripheral_RID = peripheral_RID; // @[soc.scala 120:20]
  assign core0_peripheral_RDATA = peripheral_RDATA; // @[soc.scala 120:20]
  assign core0_peripheral_RRESP = peripheral_RRESP; // @[soc.scala 120:20]
  assign core0_peripheral_RLAST = peripheral_RLAST; // @[soc.scala 120:20]
  assign core0_peripheral_RVALID = peripheral_RVALID; // @[soc.scala 120:20]
  assign core0_MTIP = MTIP; // @[soc.scala 117:14]
  assign interconnect__clock = clock;
  assign interconnect__reset = reset;
  assign interconnect__io_acePort0_AWVALID = core0_dPort_AWVALID; // @[soc.scala 135:36]
  assign interconnect__io_acePort0_AWADDR = {{32'd0}, core0_dPort_AWADDR}; // @[soc.scala 138:35]
  assign interconnect__io_acePort0_AWSNOOP = core0_dPort_AWSNOOP; // @[soc.scala 139:36]
  assign interconnect__io_acePort0_WVALID = core0_dPort_WVALID; // @[soc.scala 143:35]
  assign interconnect__io_acePort0_WDATA = core0_dPort_WDATA; // @[soc.scala 144:34]
  assign interconnect__io_acePort0_WLAST = core0_dPort_WLAST; // @[soc.scala 145:34]
  assign interconnect__io_acePort0_BREADY = core0_dPort_BREADY; // @[soc.scala 152:35]
  assign interconnect__io_acePort0_ARVALID = core0_dPort_ARVALID; // @[soc.scala 155:36]
  assign interconnect__io_acePort0_ARADDR = {{32'd0}, core0_dPort_ARADDR}; // @[soc.scala 158:35]
  assign interconnect__io_acePort0_ARSNOOP = core0_dPort_ARSNOOP; // @[soc.scala 159:36]
  assign interconnect__io_acePort0_RREADY = core0_dPort_RREADY; // @[soc.scala 164:35]
  assign interconnect__io_acePort0_ACREADY = core0_dPort_ACREADY; // @[soc.scala 175:36]
  assign interconnect__io_acePort0_CRVALID = core0_dPort_CRVALID; // @[soc.scala 178:36]
  assign interconnect__io_acePort0_CRRESP = core0_dPort_CRRESP; // @[soc.scala 179:35]
  assign interconnect__io_acePort0_CDVALID = core0_dPort_CDVALID; // @[soc.scala 183:36]
  assign interconnect__io_acePort0_CDDATA = core0_dPort_CDDATA; // @[soc.scala 185:35]
  assign interconnect__io_acePort0_CDLAST = core0_dPort_CDLAST; // @[soc.scala 186:35]
  assign interconnect__io_acePort1_ARVALID = core0_iPort_ARVALID; // @[soc.scala 210:36]
  assign interconnect__io_acePort1_ARADDR = {{32'd0}, core0_iPort_ARADDR}; // @[soc.scala 213:35]
  assign interconnect__io_acePort1_RREADY = core0_iPort_RREADY; // @[soc.scala 219:35]
  assign interconnect__io_L2_AWREADY = L2_AWREADY; // @[soc.scala 279:30]
  assign interconnect__io_L2_ARREADY = L2_ARREADY; // @[soc.scala 292:30]
  assign interconnect__io_L2_WREADY = L2_WREADY; // @[soc.scala 306:29]
  assign interconnect__io_L2_RVALID = L2_RVALID; // @[soc.scala 312:29]
  assign interconnect__io_L2_RDATA = L2_RDATA; // @[soc.scala 315:28]
  assign interconnect__io_L2_RRESP = L2_RRESP; // @[soc.scala 317:39]
  assign interconnect__io_L2_RLAST = L2_RLAST; // @[soc.scala 316:28]
  assign interconnect__io_L2_BVALID = L2_BVALID; // @[soc.scala 321:29]
  assign interconnect__io_L2_BID = L2_BID; // @[soc.scala 323:26]
  assign interconnect__io_L2_BRESP = L2_BRESP; // @[soc.scala 324:28]
endmodule
