module iCache(
  input         clock,
  input         reset,
  output        fromFetch_req_ready,
  input         fromFetch_req_valid,
  input  [63:0] fromFetch_req_bits,
  input         fromFetch_resp_ready,
  output        fromFetch_resp_valid,
  output [31:0] fromFetch_resp_bits,
  output        updateAllCachelines_ready,
  input         updateAllCachelines_fired,
  output        cachelinesUpdatesResp_ready,
  input         cachelinesUpdatesResp_fired,
  output [31:0] lowLevelMem_ARADDR,
  output        lowLevelMem_ARVALID,
  input         lowLevelMem_ARREADY,
  input  [31:0] lowLevelMem_RDATA,
  input         lowLevelMem_RLAST,
  input         lowLevelMem_RVALID,
  output        lowLevelMem_RREADY
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [127:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] cache_address; // @[ICache.scala 78:21]
  wire [31:0] cache_instruction; // @[ICache.scala 78:21]
  wire [21:0] cache_tag; // @[ICache.scala 78:21]
  wire  cache_tag_valid; // @[ICache.scala 78:21]
  wire [5:0] cache_write_line_index; // @[ICache.scala 78:21]
  wire [127:0] cache_write_block; // @[ICache.scala 78:21]
  wire [21:0] cache_write_tag; // @[ICache.scala 78:21]
  wire  cache_write_in; // @[ICache.scala 78:21]
  wire  cache_invalidate_all; // @[ICache.scala 78:21]
  wire  cache_clock; // @[ICache.scala 78:21]
  wire  cache_reset; // @[ICache.scala 78:21]
  reg  commitFence; // @[ICache.scala 63:28]
  reg  requests_0_valid; // @[ICache.scala 70:25]
  reg [63:0] requests_0_address; // @[ICache.scala 70:25]
  reg  requests_1_valid; // @[ICache.scala 70:25]
  reg [63:0] requests_1_address; // @[ICache.scala 70:25]
  reg  requests_2_valid; // @[ICache.scala 70:25]
  reg [63:0] requests_2_address; // @[ICache.scala 70:25]
  reg  results_0_valid; // @[ICache.scala 80:24]
  reg [63:0] results_0_address; // @[ICache.scala 80:24]
  reg [31:0] results_0_instruction; // @[ICache.scala 80:24]
  reg [21:0] results_0_tag; // @[ICache.scala 80:24]
  reg  results_0_tagValid; // @[ICache.scala 80:24]
  reg  results_1_valid; // @[ICache.scala 80:24]
  reg [63:0] results_1_address; // @[ICache.scala 80:24]
  reg [31:0] results_1_instruction; // @[ICache.scala 80:24]
  reg [21:0] results_1_tag; // @[ICache.scala 80:24]
  reg  results_1_tagValid; // @[ICache.scala 80:24]
  reg  cacheFill_valid; // @[ICache.scala 94:26]
  reg [127:0] cacheFill_block; // @[ICache.scala 94:26]
  wire [53:0] _GEN_44 = {{32'd0}, results_0_tag}; // @[ICache.scala 101:96]
  wire  cacheMissed = ~(results_0_tagValid & results_0_address[63:10] == _GEN_44) & results_0_valid; // @[ICache.scala 101:119]
  reg  arvalid; // @[ICache.scala 102:33]
  reg  rready; // @[ICache.scala 102:33]
  wire [127:0] _cacheFill_block_T_1 = {lowLevelMem_RDATA,cacheFill_block[127:32]}; // @[Cat.scala 33:92]
  wire  _arvalid_T = ~rready; // @[ICache.scala 106:46]
  wire  _arvalid_T_2 = ~cacheFill_valid; // @[ICache.scala 106:57]
  wire  _arvalid_T_4 = lowLevelMem_ARVALID & lowLevelMem_ARREADY; // @[ICache.scala 107:49]
  wire  _rready_T_2 = lowLevelMem_RLAST & lowLevelMem_RREADY & lowLevelMem_RVALID; // @[ICache.scala 110:68]
  wire  _GEN_3 = _arvalid_T_2 & _rready_T_2; // @[ICache.scala 112:{26,44} 113:32]
  wire  _cacheStalled_T = ~fromFetch_resp_ready; // @[ICache.scala 122:62]
  wire  cacheStalled = cacheMissed | fromFetch_resp_valid & ~fromFetch_resp_ready; // @[ICache.scala 122:34]
  wire  _T_4 = ~cacheMissed; // @[ICache.scala 123:9]
  wire [21:0] _GEN_7 = results_1_valid ? results_1_tag : cache_tag; // @[ICache.scala 124:{35,51} 129:25]
  wire  _T_9 = cacheMissed & cacheFill_valid; // @[ICache.scala 132:26]
  wire [31:0] _GEN_10 = 2'h1 == results_0_address[3:2] ? cacheFill_block[63:32] : cacheFill_block[31:0]; // @[ICache.scala 133:{31,31}]
  wire [31:0] _GEN_11 = 2'h2 == results_0_address[3:2] ? cacheFill_block[95:64] : _GEN_10; // @[ICache.scala 133:{31,31}]
  wire [22:0] _GEN_14 = cacheMissed & cacheFill_valid ? results_0_address[32:10] : {{1'd0}, results_0_tag}; // @[ICache.scala 132:46 134:23 80:24]
  wire  _GEN_15 = cacheMissed & cacheFill_valid | results_0_tagValid; // @[ICache.scala 132:46 135:28 80:24]
  wire [22:0] _GEN_19 = ~cacheMissed & (fromFetch_resp_ready | commitFence) | ~results_0_valid ? {{1'd0}, _GEN_7} :
    _GEN_14; // @[ICache.scala 123:89]
  wire  _T_10 = ~results_1_valid; // @[ICache.scala 138:8]
  wire [31:0] _GEN_22 = 2'h1 == results_1_address[3:2] ? cacheFill_block[63:32] : cacheFill_block[31:0]; // @[ICache.scala 145:{35,35}]
  wire [31:0] _GEN_23 = 2'h2 == results_1_address[3:2] ? cacheFill_block[95:64] : _GEN_22; // @[ICache.scala 145:{35,35}]
  wire  _T_16 = ~cacheStalled; // @[ICache.scala 148:14]
  wire [22:0] _GEN_27 = _T_9 & results_0_address[31:4] == results_1_address[31:4] ? results_0_address[32:10] : {{1'd0},
    results_1_tag}; // @[ICache.scala 144:157 146:27 80:24]
  wire  _GEN_28 = _T_9 & results_0_address[31:4] == results_1_address[31:4] | results_1_tagValid; // @[ICache.scala 144:157 147:32 80:24]
  wire [22:0] _GEN_33 = ~results_1_valid ? {{1'd0}, cache_tag} : _GEN_27; // @[ICache.scala 138:34 142:27]
  wire  _GEN_35 = _T_10 & (_T_16 & requests_0_valid); // @[ICache.scala 152:34 154:31 156:31]
  wire  _requests_0_valid_T = fromFetch_req_ready & fromFetch_req_valid; // @[ICache.scala 162:52]
  wire  _T_23 = ~requests_1_valid; // @[ICache.scala 167:8]
  wire  _fromFetch_req_ready_T_1 = ~commitFence; // @[ICache.scala 176:55]
  wire  _commitFence_T_3 = requests_0_valid | requests_1_valid | requests_2_valid | results_0_valid | results_1_valid; // @[ICache.scala 182:74]
  wire [22:0] _GEN_45 = reset ? 23'h0 : _GEN_19; // @[ICache.scala 80:{24,24}]
  wire [22:0] _GEN_46 = reset ? 23'h0 : _GEN_33; // @[ICache.scala 80:{24,24}]
  iCacheRegisters #(.offset_width (2), .line_width(6)) cache ( // @[ICache.scala 78:21]
    .address(cache_address),
    .instruction(cache_instruction),
    .tag(cache_tag),
    .tag_valid(cache_tag_valid),
    .write_line_index(cache_write_line_index),
    .write_block(cache_write_block),
    .write_tag(cache_write_tag),
    .write_in(cache_write_in),
    .invalidate_all(cache_invalidate_all),
    .clock(cache_clock),
    .reset(cache_reset)
  );
  assign fromFetch_req_ready = _T_23 & ~commitFence; // @[ICache.scala 176:52]
  assign fromFetch_resp_valid = _T_4 & results_0_valid; // @[ICache.scala 174:40]
  assign fromFetch_resp_bits = results_0_instruction; // @[ICache.scala 175:23]
  assign updateAllCachelines_ready = ~commitFence; // @[ICache.scala 184:32]
  assign cachelinesUpdatesResp_ready = ~_commitFence_T_3 & commitFence; // @[ICache.scala 185:96]
  assign lowLevelMem_ARADDR = {results_0_address[31:4],4'h0}; // @[Cat.scala 33:92]
  assign lowLevelMem_ARVALID = arvalid; // @[ICache.scala 198:23]
  assign lowLevelMem_RREADY = rready; // @[ICache.scala 200:22]
  assign cache_address = requests_0_address[31:0]; // @[ICache.scala 178:20]
  assign cache_write_line_index = results_0_address[9:4]; // @[ICache.scala 117:29]
  assign cache_write_block = cacheFill_block; // @[ICache.scala 115:24]
  assign cache_write_tag = results_0_address[31:10]; // @[ICache.scala 118:22]
  assign cache_write_in = cacheFill_valid; // @[ICache.scala 116:21]
  assign cache_invalidate_all = cachelinesUpdatesResp_fired; // @[ICache.scala 186:27]
  assign cache_clock = clock; // @[ICache.scala 119:18]
  assign cache_reset = reset; // @[ICache.scala 120:18]
  always @(posedge clock) begin
    if (reset) begin // @[ICache.scala 63:28]
      commitFence <= 1'h0; // @[ICache.scala 63:28]
    end else if (_fromFetch_req_ready_T_1) begin // @[ICache.scala 179:22]
      commitFence <= updateAllCachelines_fired; // @[ICache.scala 180:17]
    end else begin
      commitFence <= requests_0_valid | requests_1_valid | requests_2_valid | results_0_valid | results_1_valid | ~
        cachelinesUpdatesResp_fired; // @[ICache.scala 182:17]
    end
    if (reset) begin // @[ICache.scala 70:25]
      requests_0_valid <= 1'h0; // @[ICache.scala 70:25]
    end else if (_T_16 & _T_10 | ~requests_0_valid) begin // @[ICache.scala 159:78]
      if (requests_1_valid) begin // @[ICache.scala 160:36]
        requests_0_valid <= requests_1_valid; // @[ICache.scala 160:53]
      end else begin
        requests_0_valid <= fromFetch_req_ready & fromFetch_req_valid; // @[ICache.scala 162:28]
      end
    end
    if (reset) begin // @[ICache.scala 70:25]
      requests_0_address <= 64'h0; // @[ICache.scala 70:25]
    end else if (_T_16 & _T_10 | ~requests_0_valid) begin // @[ICache.scala 159:78]
      if (requests_1_valid) begin // @[ICache.scala 160:36]
        requests_0_address <= requests_1_address; // @[ICache.scala 160:53]
      end else begin
        requests_0_address <= fromFetch_req_bits; // @[ICache.scala 163:30]
      end
    end
    if (reset) begin // @[ICache.scala 70:25]
      requests_1_valid <= 1'h0; // @[ICache.scala 70:25]
    end else if (~requests_1_valid) begin // @[ICache.scala 167:35]
      requests_1_valid <= (cacheStalled | results_1_valid) & _requests_0_valid_T & requests_0_valid; // @[ICache.scala 168:30]
    end else begin
      requests_1_valid <= cacheStalled | results_1_valid; // @[ICache.scala 171:30]
    end
    if (reset) begin // @[ICache.scala 70:25]
      requests_1_address <= 64'h0; // @[ICache.scala 70:25]
    end else if (~requests_1_valid) begin // @[ICache.scala 167:35]
      requests_1_address <= fromFetch_req_bits; // @[ICache.scala 169:32]
    end
    if (reset) begin // @[ICache.scala 70:25]
      requests_2_valid <= 1'h0; // @[ICache.scala 70:25]
    end else begin
      requests_2_valid <= _GEN_35;
    end
    if (reset) begin // @[ICache.scala 70:25]
      requests_2_address <= 64'h0; // @[ICache.scala 70:25]
    end else if (_T_10) begin // @[ICache.scala 152:34]
      requests_2_address <= requests_0_address; // @[ICache.scala 153:25]
    end
    if (reset) begin // @[ICache.scala 80:24]
      results_0_valid <= 1'h0; // @[ICache.scala 80:24]
    end else if (~cacheMissed & (fromFetch_resp_ready | commitFence) | ~results_0_valid) begin // @[ICache.scala 123:89]
      if (results_1_valid) begin // @[ICache.scala 124:35]
        results_0_valid <= results_1_valid; // @[ICache.scala 124:51]
      end else begin
        results_0_valid <= requests_2_valid; // @[ICache.scala 126:27]
      end
    end
    if (reset) begin // @[ICache.scala 80:24]
      results_0_address <= 64'h0; // @[ICache.scala 80:24]
    end else if (~cacheMissed & (fromFetch_resp_ready | commitFence) | ~results_0_valid) begin // @[ICache.scala 123:89]
      if (results_1_valid) begin // @[ICache.scala 124:35]
        results_0_address <= results_1_address; // @[ICache.scala 124:51]
      end else begin
        results_0_address <= requests_2_address; // @[ICache.scala 127:29]
      end
    end
    if (reset) begin // @[ICache.scala 80:24]
      results_0_instruction <= 32'h0; // @[ICache.scala 80:24]
    end else if (~cacheMissed & (fromFetch_resp_ready | commitFence) | ~results_0_valid) begin // @[ICache.scala 123:89]
      if (results_1_valid) begin // @[ICache.scala 124:35]
        results_0_instruction <= results_1_instruction; // @[ICache.scala 124:51]
      end else begin
        results_0_instruction <= cache_instruction; // @[ICache.scala 128:33]
      end
    end else if (cacheMissed & cacheFill_valid) begin // @[ICache.scala 132:46]
      if (2'h3 == results_0_address[3:2]) begin // @[ICache.scala 133:31]
        results_0_instruction <= cacheFill_block[127:96]; // @[ICache.scala 133:31]
      end else begin
        results_0_instruction <= _GEN_11;
      end
    end
    results_0_tag <= _GEN_45[21:0]; // @[ICache.scala 80:{24,24}]
    if (reset) begin // @[ICache.scala 80:24]
      results_0_tagValid <= 1'h0; // @[ICache.scala 80:24]
    end else if (~cacheMissed & (fromFetch_resp_ready | commitFence) | ~results_0_valid) begin // @[ICache.scala 123:89]
      if (results_1_valid) begin // @[ICache.scala 124:35]
        results_0_tagValid <= results_1_tagValid; // @[ICache.scala 124:51]
      end else begin
        results_0_tagValid <= cache_tag_valid; // @[ICache.scala 130:30]
      end
    end else begin
      results_0_tagValid <= _GEN_15;
    end
    if (reset) begin // @[ICache.scala 80:24]
      results_1_valid <= 1'h0; // @[ICache.scala 80:24]
    end else if (~results_1_valid) begin // @[ICache.scala 138:34]
      results_1_valid <= requests_2_valid & results_0_valid & (cacheMissed | _cacheStalled_T); // @[ICache.scala 139:29]
    end else if (!(_T_9 & results_0_address[31:4] == results_1_address[31:4])) begin // @[ICache.scala 144:157]
      if (~cacheStalled) begin // @[ICache.scala 148:29]
        results_1_valid <= 1'h0; // @[ICache.scala 149:29]
      end
    end
    if (reset) begin // @[ICache.scala 80:24]
      results_1_address <= 64'h0; // @[ICache.scala 80:24]
    end else if (~results_1_valid) begin // @[ICache.scala 138:34]
      results_1_address <= requests_2_address; // @[ICache.scala 140:31]
    end
    if (reset) begin // @[ICache.scala 80:24]
      results_1_instruction <= 32'h0; // @[ICache.scala 80:24]
    end else if (~results_1_valid) begin // @[ICache.scala 138:34]
      results_1_instruction <= cache_instruction; // @[ICache.scala 141:35]
    end else if (_T_9 & results_0_address[31:4] == results_1_address[31:4]) begin // @[ICache.scala 144:157]
      if (2'h3 == results_1_address[3:2]) begin // @[ICache.scala 145:35]
        results_1_instruction <= cacheFill_block[127:96]; // @[ICache.scala 145:35]
      end else begin
        results_1_instruction <= _GEN_23;
      end
    end
    results_1_tag <= _GEN_46[21:0]; // @[ICache.scala 80:{24,24}]
    if (reset) begin // @[ICache.scala 80:24]
      results_1_tagValid <= 1'h0; // @[ICache.scala 80:24]
    end else if (~results_1_valid) begin // @[ICache.scala 138:34]
      results_1_tagValid <= cache_tag_valid; // @[ICache.scala 143:32]
    end else begin
      results_1_tagValid <= _GEN_28;
    end
    if (reset) begin // @[ICache.scala 94:26]
      cacheFill_valid <= 1'h0; // @[ICache.scala 94:26]
    end else begin
      cacheFill_valid <= _GEN_3;
    end
    if (reset) begin // @[ICache.scala 94:26]
      cacheFill_block <= 128'h0; // @[ICache.scala 94:26]
    end else if (lowLevelMem_RREADY & lowLevelMem_RVALID) begin // @[ICache.scala 104:50]
      cacheFill_block <= _cacheFill_block_T_1; // @[ICache.scala 104:68]
    end
    if (reset) begin // @[ICache.scala 102:33]
      arvalid <= 1'h0; // @[ICache.scala 102:33]
    end else if (~arvalid) begin // @[ICache.scala 106:18]
      arvalid <= cacheMissed & ~rready & ~cacheFill_valid; // @[ICache.scala 106:28]
    end else begin
      arvalid <= ~(lowLevelMem_ARVALID & lowLevelMem_ARREADY); // @[ICache.scala 107:24]
    end
    if (reset) begin // @[ICache.scala 102:33]
      rready <= 1'h0; // @[ICache.scala 102:33]
    end else if (_arvalid_T) begin // @[ICache.scala 109:17]
      rready <= _arvalid_T_4; // @[ICache.scala 109:26]
    end else begin
      rready <= ~(lowLevelMem_RLAST & lowLevelMem_RREADY & lowLevelMem_RVALID); // @[ICache.scala 110:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  commitFence = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  requests_0_valid = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  requests_0_address = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  requests_1_valid = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  requests_1_address = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  requests_2_valid = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  requests_2_address = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  results_0_valid = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  results_0_address = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  results_0_instruction = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  results_0_tag = _RAND_10[21:0];
  _RAND_11 = {1{`RANDOM}};
  results_0_tagValid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  results_1_valid = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  results_1_address = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  results_1_instruction = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  results_1_tag = _RAND_15[21:0];
  _RAND_16 = {1{`RANDOM}};
  results_1_tagValid = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  cacheFill_valid = _RAND_17[0:0];
  _RAND_18 = {4{`RANDOM}};
  cacheFill_block = _RAND_18[127:0];
  _RAND_19 = {1{`RANDOM}};
  arvalid = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  rready = _RAND_20[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module shiftReg(
  input   clock,
  input   reset,
  input   in,
  input   en,
  output  output_0,
  output  output_1,
  output  output_2,
  output  output_3,
  output  output_4
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  shiftregs_0; // @[fetch.scala 89:56]
  reg  shiftregs_1; // @[fetch.scala 89:56]
  reg  shiftregs_2; // @[fetch.scala 89:56]
  reg  shiftregs_3; // @[fetch.scala 89:56]
  reg  shiftregs_4; // @[fetch.scala 89:56]
  assign output_0 = shiftregs_0; // @[fetch.scala 98:54]
  assign output_1 = shiftregs_1; // @[fetch.scala 98:54]
  assign output_2 = shiftregs_2; // @[fetch.scala 98:54]
  assign output_3 = shiftregs_3; // @[fetch.scala 98:54]
  assign output_4 = shiftregs_4; // @[fetch.scala 98:54]
  always @(posedge clock) begin
    if (reset) begin // @[fetch.scala 89:56]
      shiftregs_0 <= 1'h0; // @[fetch.scala 89:56]
    end else if (en) begin // @[fetch.scala 91:14]
      shiftregs_0 <= in; // @[fetch.scala 92:20]
    end
    if (reset) begin // @[fetch.scala 89:56]
      shiftregs_1 <= 1'h0; // @[fetch.scala 89:56]
    end else if (en) begin // @[fetch.scala 91:14]
      shiftregs_1 <= shiftregs_0; // @[fetch.scala 94:22]
    end
    if (reset) begin // @[fetch.scala 89:56]
      shiftregs_2 <= 1'h0; // @[fetch.scala 89:56]
    end else if (en) begin // @[fetch.scala 91:14]
      shiftregs_2 <= shiftregs_1; // @[fetch.scala 94:22]
    end
    if (reset) begin // @[fetch.scala 89:56]
      shiftregs_3 <= 1'h0; // @[fetch.scala 89:56]
    end else if (en) begin // @[fetch.scala 91:14]
      shiftregs_3 <= shiftregs_2; // @[fetch.scala 94:22]
    end
    if (reset) begin // @[fetch.scala 89:56]
      shiftregs_4 <= 1'h0; // @[fetch.scala 89:56]
    end else if (en) begin // @[fetch.scala 91:14]
      shiftregs_4 <= shiftregs_3; // @[fetch.scala 94:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shiftregs_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  shiftregs_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  shiftregs_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  shiftregs_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  shiftregs_4 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module updateShiftReg(
  input   clock,
  input   reset,
  input   in,
  input   en,
  output  output_0,
  output  output_1,
  output  output_2,
  output  output_3,
  output  output_4,
  input   updateVals_0,
  input   updateVals_1,
  input   updateVals_2,
  input   updateVals_3,
  input   updateVals_4,
  input   update
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  shiftregs_0; // @[fetch.scala 89:56]
  reg  shiftregs_1; // @[fetch.scala 89:56]
  reg  shiftregs_2; // @[fetch.scala 89:56]
  reg  shiftregs_3; // @[fetch.scala 89:56]
  reg  shiftregs_4; // @[fetch.scala 89:56]
  assign output_0 = shiftregs_0; // @[fetch.scala 98:54]
  assign output_1 = shiftregs_1; // @[fetch.scala 98:54]
  assign output_2 = shiftregs_2; // @[fetch.scala 98:54]
  assign output_3 = shiftregs_3; // @[fetch.scala 98:54]
  assign output_4 = shiftregs_4; // @[fetch.scala 98:54]
  always @(posedge clock) begin
    if (reset) begin // @[fetch.scala 89:56]
      shiftregs_0 <= 1'h0; // @[fetch.scala 89:56]
    end else if (update) begin // @[fetch.scala 105:17]
      shiftregs_0 <= updateVals_0; // @[fetch.scala 106:48]
    end else if (en) begin // @[fetch.scala 91:14]
      shiftregs_0 <= in; // @[fetch.scala 92:20]
    end
    if (reset) begin // @[fetch.scala 89:56]
      shiftregs_1 <= 1'h0; // @[fetch.scala 89:56]
    end else if (update) begin // @[fetch.scala 105:17]
      shiftregs_1 <= updateVals_1; // @[fetch.scala 106:48]
    end else if (en) begin // @[fetch.scala 91:14]
      shiftregs_1 <= shiftregs_0; // @[fetch.scala 94:22]
    end
    if (reset) begin // @[fetch.scala 89:56]
      shiftregs_2 <= 1'h0; // @[fetch.scala 89:56]
    end else if (update) begin // @[fetch.scala 105:17]
      shiftregs_2 <= updateVals_2; // @[fetch.scala 106:48]
    end else if (en) begin // @[fetch.scala 91:14]
      shiftregs_2 <= shiftregs_1; // @[fetch.scala 94:22]
    end
    if (reset) begin // @[fetch.scala 89:56]
      shiftregs_3 <= 1'h0; // @[fetch.scala 89:56]
    end else if (update) begin // @[fetch.scala 105:17]
      shiftregs_3 <= updateVals_3; // @[fetch.scala 106:48]
    end else if (en) begin // @[fetch.scala 91:14]
      shiftregs_3 <= shiftregs_2; // @[fetch.scala 94:22]
    end
    if (reset) begin // @[fetch.scala 89:56]
      shiftregs_4 <= 1'h0; // @[fetch.scala 89:56]
    end else if (update) begin // @[fetch.scala 105:17]
      shiftregs_4 <= updateVals_4; // @[fetch.scala 106:48]
    end else if (en) begin // @[fetch.scala 91:14]
      shiftregs_4 <= shiftregs_3; // @[fetch.scala 94:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shiftregs_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  shiftregs_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  shiftregs_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  shiftregs_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  shiftregs_4 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module gshare_predictor(
  input         clock,
  input         reset,
  input         io_branchres_fired,
  input         io_branchres_branchTaken,
  input  [63:0] io_branchres_pc,
  input  [63:0] io_branchres_pcAfterBrnach,
  input  [63:0] io_curr_pc,
  output [63:0] io_next_pc,
  input         requestSent,
  input         mispredicted
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
`endif // RANDOMIZE_REG_INIT
  wire  correct_history_clock; // @[fetch.scala 120:31]
  wire  correct_history_reset; // @[fetch.scala 120:31]
  wire  correct_history_in; // @[fetch.scala 120:31]
  wire  correct_history_en; // @[fetch.scala 120:31]
  wire  correct_history_output_0; // @[fetch.scala 120:31]
  wire  correct_history_output_1; // @[fetch.scala 120:31]
  wire  correct_history_output_2; // @[fetch.scala 120:31]
  wire  correct_history_output_3; // @[fetch.scala 120:31]
  wire  correct_history_output_4; // @[fetch.scala 120:31]
  wire  predicted_history_clock; // @[fetch.scala 121:33]
  wire  predicted_history_reset; // @[fetch.scala 121:33]
  wire  predicted_history_in; // @[fetch.scala 121:33]
  wire  predicted_history_en; // @[fetch.scala 121:33]
  wire  predicted_history_output_0; // @[fetch.scala 121:33]
  wire  predicted_history_output_1; // @[fetch.scala 121:33]
  wire  predicted_history_output_2; // @[fetch.scala 121:33]
  wire  predicted_history_output_3; // @[fetch.scala 121:33]
  wire  predicted_history_output_4; // @[fetch.scala 121:33]
  wire  predicted_history_updateVals_0; // @[fetch.scala 121:33]
  wire  predicted_history_updateVals_1; // @[fetch.scala 121:33]
  wire  predicted_history_updateVals_2; // @[fetch.scala 121:33]
  wire  predicted_history_updateVals_3; // @[fetch.scala 121:33]
  wire  predicted_history_updateVals_4; // @[fetch.scala 121:33]
  wire  predicted_history_update; // @[fetch.scala 121:33]
  reg [63:0] btb [0:255]; // @[fetch.scala 145:16]
  wire  btb_io_next_pc_MPORT_en; // @[fetch.scala 145:16]
  wire [7:0] btb_io_next_pc_MPORT_addr; // @[fetch.scala 145:16]
  wire [63:0] btb_io_next_pc_MPORT_data; // @[fetch.scala 145:16]
  wire [63:0] btb_MPORT_1_data; // @[fetch.scala 145:16]
  wire [7:0] btb_MPORT_1_addr; // @[fetch.scala 145:16]
  wire  btb_MPORT_1_mask; // @[fetch.scala 145:16]
  wire  btb_MPORT_1_en; // @[fetch.scala 145:16]
  reg [1:0] counters [0:2047]; // @[fetch.scala 146:21]
  wire  counters_MPORT_2_en; // @[fetch.scala 146:21]
  wire [10:0] counters_MPORT_2_addr; // @[fetch.scala 146:21]
  wire [1:0] counters_MPORT_2_data; // @[fetch.scala 146:21]
  wire  counters_MPORT_4_en; // @[fetch.scala 146:21]
  wire [10:0] counters_MPORT_4_addr; // @[fetch.scala 146:21]
  wire [1:0] counters_MPORT_4_data; // @[fetch.scala 146:21]
  wire  counters_MPORT_5_en; // @[fetch.scala 146:21]
  wire [10:0] counters_MPORT_5_addr; // @[fetch.scala 146:21]
  wire [1:0] counters_MPORT_5_data; // @[fetch.scala 146:21]
  wire  counters_MPORT_7_en; // @[fetch.scala 146:21]
  wire [10:0] counters_MPORT_7_addr; // @[fetch.scala 146:21]
  wire [1:0] counters_MPORT_7_data; // @[fetch.scala 146:21]
  wire  counters_prediction_MPORT_en; // @[fetch.scala 146:21]
  wire [10:0] counters_prediction_MPORT_addr; // @[fetch.scala 146:21]
  wire [1:0] counters_prediction_MPORT_data; // @[fetch.scala 146:21]
  wire [1:0] counters_MPORT_3_data; // @[fetch.scala 146:21]
  wire [10:0] counters_MPORT_3_addr; // @[fetch.scala 146:21]
  wire  counters_MPORT_3_mask; // @[fetch.scala 146:21]
  wire  counters_MPORT_3_en; // @[fetch.scala 146:21]
  wire [1:0] counters_MPORT_6_data; // @[fetch.scala 146:21]
  wire [10:0] counters_MPORT_6_addr; // @[fetch.scala 146:21]
  wire  counters_MPORT_6_mask; // @[fetch.scala 146:21]
  wire  counters_MPORT_6_en; // @[fetch.scala 146:21]
  reg [53:0] tag_store [0:255]; // @[fetch.scala 148:22]
  wire  tag_store_btb_hit_MPORT_en; // @[fetch.scala 148:22]
  wire [7:0] tag_store_btb_hit_MPORT_addr; // @[fetch.scala 148:22]
  wire [53:0] tag_store_btb_hit_MPORT_data; // @[fetch.scala 148:22]
  wire [53:0] tag_store_MPORT_data; // @[fetch.scala 148:22]
  wire [7:0] tag_store_MPORT_addr; // @[fetch.scala 148:22]
  wire  tag_store_MPORT_mask; // @[fetch.scala 148:22]
  wire  tag_store_MPORT_en; // @[fetch.scala 148:22]
  wire [4:0] _counterIndex_pred_T_2 = {predicted_history_output_4,predicted_history_output_3,predicted_history_output_2,
    predicted_history_output_1,predicted_history_output_0}; // @[fetch.scala 130:178]
  wire [4:0] _counterIndex_pred_T_14 = {_counterIndex_pred_T_2[0],_counterIndex_pred_T_2[1],_counterIndex_pred_T_2[2],
    _counterIndex_pred_T_2[3],_counterIndex_pred_T_2[4]}; // @[Cat.scala 33:92]
  wire [4:0] _counterIndex_pred_T_15 = io_curr_pc[6:2] ^ _counterIndex_pred_T_14; // @[fetch.scala 130:143]
  wire [4:0] _counterIndex_train_T_2 = {correct_history_output_4,correct_history_output_3,correct_history_output_2,
    correct_history_output_1,correct_history_output_0}; // @[fetch.scala 131:187]
  wire [4:0] _counterIndex_train_T_14 = {_counterIndex_train_T_2[0],_counterIndex_train_T_2[1],_counterIndex_train_T_2[2
    ],_counterIndex_train_T_2[3],_counterIndex_train_T_2[4]}; // @[Cat.scala 33:92]
  wire [4:0] _counterIndex_train_T_15 = io_branchres_pc[6:2] ^ _counterIndex_train_T_14; // @[fetch.scala 131:154]
  wire [7:0] btb_addr = io_curr_pc[9:2]; // @[fetch.scala 139:28]
  wire [53:0] tag = io_curr_pc[63:10]; // @[fetch.scala 140:23]
  wire [7:0] result_addr = io_branchres_pc[9:2]; // @[fetch.scala 141:36]
  reg  valid_bits_0; // @[fetch.scala 147:27]
  reg  valid_bits_1; // @[fetch.scala 147:27]
  reg  valid_bits_2; // @[fetch.scala 147:27]
  reg  valid_bits_3; // @[fetch.scala 147:27]
  reg  valid_bits_4; // @[fetch.scala 147:27]
  reg  valid_bits_5; // @[fetch.scala 147:27]
  reg  valid_bits_6; // @[fetch.scala 147:27]
  reg  valid_bits_7; // @[fetch.scala 147:27]
  reg  valid_bits_8; // @[fetch.scala 147:27]
  reg  valid_bits_9; // @[fetch.scala 147:27]
  reg  valid_bits_10; // @[fetch.scala 147:27]
  reg  valid_bits_11; // @[fetch.scala 147:27]
  reg  valid_bits_12; // @[fetch.scala 147:27]
  reg  valid_bits_13; // @[fetch.scala 147:27]
  reg  valid_bits_14; // @[fetch.scala 147:27]
  reg  valid_bits_15; // @[fetch.scala 147:27]
  reg  valid_bits_16; // @[fetch.scala 147:27]
  reg  valid_bits_17; // @[fetch.scala 147:27]
  reg  valid_bits_18; // @[fetch.scala 147:27]
  reg  valid_bits_19; // @[fetch.scala 147:27]
  reg  valid_bits_20; // @[fetch.scala 147:27]
  reg  valid_bits_21; // @[fetch.scala 147:27]
  reg  valid_bits_22; // @[fetch.scala 147:27]
  reg  valid_bits_23; // @[fetch.scala 147:27]
  reg  valid_bits_24; // @[fetch.scala 147:27]
  reg  valid_bits_25; // @[fetch.scala 147:27]
  reg  valid_bits_26; // @[fetch.scala 147:27]
  reg  valid_bits_27; // @[fetch.scala 147:27]
  reg  valid_bits_28; // @[fetch.scala 147:27]
  reg  valid_bits_29; // @[fetch.scala 147:27]
  reg  valid_bits_30; // @[fetch.scala 147:27]
  reg  valid_bits_31; // @[fetch.scala 147:27]
  reg  valid_bits_32; // @[fetch.scala 147:27]
  reg  valid_bits_33; // @[fetch.scala 147:27]
  reg  valid_bits_34; // @[fetch.scala 147:27]
  reg  valid_bits_35; // @[fetch.scala 147:27]
  reg  valid_bits_36; // @[fetch.scala 147:27]
  reg  valid_bits_37; // @[fetch.scala 147:27]
  reg  valid_bits_38; // @[fetch.scala 147:27]
  reg  valid_bits_39; // @[fetch.scala 147:27]
  reg  valid_bits_40; // @[fetch.scala 147:27]
  reg  valid_bits_41; // @[fetch.scala 147:27]
  reg  valid_bits_42; // @[fetch.scala 147:27]
  reg  valid_bits_43; // @[fetch.scala 147:27]
  reg  valid_bits_44; // @[fetch.scala 147:27]
  reg  valid_bits_45; // @[fetch.scala 147:27]
  reg  valid_bits_46; // @[fetch.scala 147:27]
  reg  valid_bits_47; // @[fetch.scala 147:27]
  reg  valid_bits_48; // @[fetch.scala 147:27]
  reg  valid_bits_49; // @[fetch.scala 147:27]
  reg  valid_bits_50; // @[fetch.scala 147:27]
  reg  valid_bits_51; // @[fetch.scala 147:27]
  reg  valid_bits_52; // @[fetch.scala 147:27]
  reg  valid_bits_53; // @[fetch.scala 147:27]
  reg  valid_bits_54; // @[fetch.scala 147:27]
  reg  valid_bits_55; // @[fetch.scala 147:27]
  reg  valid_bits_56; // @[fetch.scala 147:27]
  reg  valid_bits_57; // @[fetch.scala 147:27]
  reg  valid_bits_58; // @[fetch.scala 147:27]
  reg  valid_bits_59; // @[fetch.scala 147:27]
  reg  valid_bits_60; // @[fetch.scala 147:27]
  reg  valid_bits_61; // @[fetch.scala 147:27]
  reg  valid_bits_62; // @[fetch.scala 147:27]
  reg  valid_bits_63; // @[fetch.scala 147:27]
  reg  valid_bits_64; // @[fetch.scala 147:27]
  reg  valid_bits_65; // @[fetch.scala 147:27]
  reg  valid_bits_66; // @[fetch.scala 147:27]
  reg  valid_bits_67; // @[fetch.scala 147:27]
  reg  valid_bits_68; // @[fetch.scala 147:27]
  reg  valid_bits_69; // @[fetch.scala 147:27]
  reg  valid_bits_70; // @[fetch.scala 147:27]
  reg  valid_bits_71; // @[fetch.scala 147:27]
  reg  valid_bits_72; // @[fetch.scala 147:27]
  reg  valid_bits_73; // @[fetch.scala 147:27]
  reg  valid_bits_74; // @[fetch.scala 147:27]
  reg  valid_bits_75; // @[fetch.scala 147:27]
  reg  valid_bits_76; // @[fetch.scala 147:27]
  reg  valid_bits_77; // @[fetch.scala 147:27]
  reg  valid_bits_78; // @[fetch.scala 147:27]
  reg  valid_bits_79; // @[fetch.scala 147:27]
  reg  valid_bits_80; // @[fetch.scala 147:27]
  reg  valid_bits_81; // @[fetch.scala 147:27]
  reg  valid_bits_82; // @[fetch.scala 147:27]
  reg  valid_bits_83; // @[fetch.scala 147:27]
  reg  valid_bits_84; // @[fetch.scala 147:27]
  reg  valid_bits_85; // @[fetch.scala 147:27]
  reg  valid_bits_86; // @[fetch.scala 147:27]
  reg  valid_bits_87; // @[fetch.scala 147:27]
  reg  valid_bits_88; // @[fetch.scala 147:27]
  reg  valid_bits_89; // @[fetch.scala 147:27]
  reg  valid_bits_90; // @[fetch.scala 147:27]
  reg  valid_bits_91; // @[fetch.scala 147:27]
  reg  valid_bits_92; // @[fetch.scala 147:27]
  reg  valid_bits_93; // @[fetch.scala 147:27]
  reg  valid_bits_94; // @[fetch.scala 147:27]
  reg  valid_bits_95; // @[fetch.scala 147:27]
  reg  valid_bits_96; // @[fetch.scala 147:27]
  reg  valid_bits_97; // @[fetch.scala 147:27]
  reg  valid_bits_98; // @[fetch.scala 147:27]
  reg  valid_bits_99; // @[fetch.scala 147:27]
  reg  valid_bits_100; // @[fetch.scala 147:27]
  reg  valid_bits_101; // @[fetch.scala 147:27]
  reg  valid_bits_102; // @[fetch.scala 147:27]
  reg  valid_bits_103; // @[fetch.scala 147:27]
  reg  valid_bits_104; // @[fetch.scala 147:27]
  reg  valid_bits_105; // @[fetch.scala 147:27]
  reg  valid_bits_106; // @[fetch.scala 147:27]
  reg  valid_bits_107; // @[fetch.scala 147:27]
  reg  valid_bits_108; // @[fetch.scala 147:27]
  reg  valid_bits_109; // @[fetch.scala 147:27]
  reg  valid_bits_110; // @[fetch.scala 147:27]
  reg  valid_bits_111; // @[fetch.scala 147:27]
  reg  valid_bits_112; // @[fetch.scala 147:27]
  reg  valid_bits_113; // @[fetch.scala 147:27]
  reg  valid_bits_114; // @[fetch.scala 147:27]
  reg  valid_bits_115; // @[fetch.scala 147:27]
  reg  valid_bits_116; // @[fetch.scala 147:27]
  reg  valid_bits_117; // @[fetch.scala 147:27]
  reg  valid_bits_118; // @[fetch.scala 147:27]
  reg  valid_bits_119; // @[fetch.scala 147:27]
  reg  valid_bits_120; // @[fetch.scala 147:27]
  reg  valid_bits_121; // @[fetch.scala 147:27]
  reg  valid_bits_122; // @[fetch.scala 147:27]
  reg  valid_bits_123; // @[fetch.scala 147:27]
  reg  valid_bits_124; // @[fetch.scala 147:27]
  reg  valid_bits_125; // @[fetch.scala 147:27]
  reg  valid_bits_126; // @[fetch.scala 147:27]
  reg  valid_bits_127; // @[fetch.scala 147:27]
  reg  valid_bits_128; // @[fetch.scala 147:27]
  reg  valid_bits_129; // @[fetch.scala 147:27]
  reg  valid_bits_130; // @[fetch.scala 147:27]
  reg  valid_bits_131; // @[fetch.scala 147:27]
  reg  valid_bits_132; // @[fetch.scala 147:27]
  reg  valid_bits_133; // @[fetch.scala 147:27]
  reg  valid_bits_134; // @[fetch.scala 147:27]
  reg  valid_bits_135; // @[fetch.scala 147:27]
  reg  valid_bits_136; // @[fetch.scala 147:27]
  reg  valid_bits_137; // @[fetch.scala 147:27]
  reg  valid_bits_138; // @[fetch.scala 147:27]
  reg  valid_bits_139; // @[fetch.scala 147:27]
  reg  valid_bits_140; // @[fetch.scala 147:27]
  reg  valid_bits_141; // @[fetch.scala 147:27]
  reg  valid_bits_142; // @[fetch.scala 147:27]
  reg  valid_bits_143; // @[fetch.scala 147:27]
  reg  valid_bits_144; // @[fetch.scala 147:27]
  reg  valid_bits_145; // @[fetch.scala 147:27]
  reg  valid_bits_146; // @[fetch.scala 147:27]
  reg  valid_bits_147; // @[fetch.scala 147:27]
  reg  valid_bits_148; // @[fetch.scala 147:27]
  reg  valid_bits_149; // @[fetch.scala 147:27]
  reg  valid_bits_150; // @[fetch.scala 147:27]
  reg  valid_bits_151; // @[fetch.scala 147:27]
  reg  valid_bits_152; // @[fetch.scala 147:27]
  reg  valid_bits_153; // @[fetch.scala 147:27]
  reg  valid_bits_154; // @[fetch.scala 147:27]
  reg  valid_bits_155; // @[fetch.scala 147:27]
  reg  valid_bits_156; // @[fetch.scala 147:27]
  reg  valid_bits_157; // @[fetch.scala 147:27]
  reg  valid_bits_158; // @[fetch.scala 147:27]
  reg  valid_bits_159; // @[fetch.scala 147:27]
  reg  valid_bits_160; // @[fetch.scala 147:27]
  reg  valid_bits_161; // @[fetch.scala 147:27]
  reg  valid_bits_162; // @[fetch.scala 147:27]
  reg  valid_bits_163; // @[fetch.scala 147:27]
  reg  valid_bits_164; // @[fetch.scala 147:27]
  reg  valid_bits_165; // @[fetch.scala 147:27]
  reg  valid_bits_166; // @[fetch.scala 147:27]
  reg  valid_bits_167; // @[fetch.scala 147:27]
  reg  valid_bits_168; // @[fetch.scala 147:27]
  reg  valid_bits_169; // @[fetch.scala 147:27]
  reg  valid_bits_170; // @[fetch.scala 147:27]
  reg  valid_bits_171; // @[fetch.scala 147:27]
  reg  valid_bits_172; // @[fetch.scala 147:27]
  reg  valid_bits_173; // @[fetch.scala 147:27]
  reg  valid_bits_174; // @[fetch.scala 147:27]
  reg  valid_bits_175; // @[fetch.scala 147:27]
  reg  valid_bits_176; // @[fetch.scala 147:27]
  reg  valid_bits_177; // @[fetch.scala 147:27]
  reg  valid_bits_178; // @[fetch.scala 147:27]
  reg  valid_bits_179; // @[fetch.scala 147:27]
  reg  valid_bits_180; // @[fetch.scala 147:27]
  reg  valid_bits_181; // @[fetch.scala 147:27]
  reg  valid_bits_182; // @[fetch.scala 147:27]
  reg  valid_bits_183; // @[fetch.scala 147:27]
  reg  valid_bits_184; // @[fetch.scala 147:27]
  reg  valid_bits_185; // @[fetch.scala 147:27]
  reg  valid_bits_186; // @[fetch.scala 147:27]
  reg  valid_bits_187; // @[fetch.scala 147:27]
  reg  valid_bits_188; // @[fetch.scala 147:27]
  reg  valid_bits_189; // @[fetch.scala 147:27]
  reg  valid_bits_190; // @[fetch.scala 147:27]
  reg  valid_bits_191; // @[fetch.scala 147:27]
  reg  valid_bits_192; // @[fetch.scala 147:27]
  reg  valid_bits_193; // @[fetch.scala 147:27]
  reg  valid_bits_194; // @[fetch.scala 147:27]
  reg  valid_bits_195; // @[fetch.scala 147:27]
  reg  valid_bits_196; // @[fetch.scala 147:27]
  reg  valid_bits_197; // @[fetch.scala 147:27]
  reg  valid_bits_198; // @[fetch.scala 147:27]
  reg  valid_bits_199; // @[fetch.scala 147:27]
  reg  valid_bits_200; // @[fetch.scala 147:27]
  reg  valid_bits_201; // @[fetch.scala 147:27]
  reg  valid_bits_202; // @[fetch.scala 147:27]
  reg  valid_bits_203; // @[fetch.scala 147:27]
  reg  valid_bits_204; // @[fetch.scala 147:27]
  reg  valid_bits_205; // @[fetch.scala 147:27]
  reg  valid_bits_206; // @[fetch.scala 147:27]
  reg  valid_bits_207; // @[fetch.scala 147:27]
  reg  valid_bits_208; // @[fetch.scala 147:27]
  reg  valid_bits_209; // @[fetch.scala 147:27]
  reg  valid_bits_210; // @[fetch.scala 147:27]
  reg  valid_bits_211; // @[fetch.scala 147:27]
  reg  valid_bits_212; // @[fetch.scala 147:27]
  reg  valid_bits_213; // @[fetch.scala 147:27]
  reg  valid_bits_214; // @[fetch.scala 147:27]
  reg  valid_bits_215; // @[fetch.scala 147:27]
  reg  valid_bits_216; // @[fetch.scala 147:27]
  reg  valid_bits_217; // @[fetch.scala 147:27]
  reg  valid_bits_218; // @[fetch.scala 147:27]
  reg  valid_bits_219; // @[fetch.scala 147:27]
  reg  valid_bits_220; // @[fetch.scala 147:27]
  reg  valid_bits_221; // @[fetch.scala 147:27]
  reg  valid_bits_222; // @[fetch.scala 147:27]
  reg  valid_bits_223; // @[fetch.scala 147:27]
  reg  valid_bits_224; // @[fetch.scala 147:27]
  reg  valid_bits_225; // @[fetch.scala 147:27]
  reg  valid_bits_226; // @[fetch.scala 147:27]
  reg  valid_bits_227; // @[fetch.scala 147:27]
  reg  valid_bits_228; // @[fetch.scala 147:27]
  reg  valid_bits_229; // @[fetch.scala 147:27]
  reg  valid_bits_230; // @[fetch.scala 147:27]
  reg  valid_bits_231; // @[fetch.scala 147:27]
  reg  valid_bits_232; // @[fetch.scala 147:27]
  reg  valid_bits_233; // @[fetch.scala 147:27]
  reg  valid_bits_234; // @[fetch.scala 147:27]
  reg  valid_bits_235; // @[fetch.scala 147:27]
  reg  valid_bits_236; // @[fetch.scala 147:27]
  reg  valid_bits_237; // @[fetch.scala 147:27]
  reg  valid_bits_238; // @[fetch.scala 147:27]
  reg  valid_bits_239; // @[fetch.scala 147:27]
  reg  valid_bits_240; // @[fetch.scala 147:27]
  reg  valid_bits_241; // @[fetch.scala 147:27]
  reg  valid_bits_242; // @[fetch.scala 147:27]
  reg  valid_bits_243; // @[fetch.scala 147:27]
  reg  valid_bits_244; // @[fetch.scala 147:27]
  reg  valid_bits_245; // @[fetch.scala 147:27]
  reg  valid_bits_246; // @[fetch.scala 147:27]
  reg  valid_bits_247; // @[fetch.scala 147:27]
  reg  valid_bits_248; // @[fetch.scala 147:27]
  reg  valid_bits_249; // @[fetch.scala 147:27]
  reg  valid_bits_250; // @[fetch.scala 147:27]
  reg  valid_bits_251; // @[fetch.scala 147:27]
  reg  valid_bits_252; // @[fetch.scala 147:27]
  reg  valid_bits_253; // @[fetch.scala 147:27]
  reg  valid_bits_254; // @[fetch.scala 147:27]
  reg  valid_bits_255; // @[fetch.scala 147:27]
  wire  _GEN_0 = 8'h0 == result_addr | valid_bits_0; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_1 = 8'h1 == result_addr | valid_bits_1; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_2 = 8'h2 == result_addr | valid_bits_2; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_3 = 8'h3 == result_addr | valid_bits_3; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_4 = 8'h4 == result_addr | valid_bits_4; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_5 = 8'h5 == result_addr | valid_bits_5; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_6 = 8'h6 == result_addr | valid_bits_6; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_7 = 8'h7 == result_addr | valid_bits_7; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_8 = 8'h8 == result_addr | valid_bits_8; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_9 = 8'h9 == result_addr | valid_bits_9; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_10 = 8'ha == result_addr | valid_bits_10; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_11 = 8'hb == result_addr | valid_bits_11; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_12 = 8'hc == result_addr | valid_bits_12; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_13 = 8'hd == result_addr | valid_bits_13; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_14 = 8'he == result_addr | valid_bits_14; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_15 = 8'hf == result_addr | valid_bits_15; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_16 = 8'h10 == result_addr | valid_bits_16; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_17 = 8'h11 == result_addr | valid_bits_17; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_18 = 8'h12 == result_addr | valid_bits_18; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_19 = 8'h13 == result_addr | valid_bits_19; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_20 = 8'h14 == result_addr | valid_bits_20; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_21 = 8'h15 == result_addr | valid_bits_21; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_22 = 8'h16 == result_addr | valid_bits_22; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_23 = 8'h17 == result_addr | valid_bits_23; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_24 = 8'h18 == result_addr | valid_bits_24; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_25 = 8'h19 == result_addr | valid_bits_25; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_26 = 8'h1a == result_addr | valid_bits_26; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_27 = 8'h1b == result_addr | valid_bits_27; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_28 = 8'h1c == result_addr | valid_bits_28; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_29 = 8'h1d == result_addr | valid_bits_29; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_30 = 8'h1e == result_addr | valid_bits_30; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_31 = 8'h1f == result_addr | valid_bits_31; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_32 = 8'h20 == result_addr | valid_bits_32; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_33 = 8'h21 == result_addr | valid_bits_33; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_34 = 8'h22 == result_addr | valid_bits_34; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_35 = 8'h23 == result_addr | valid_bits_35; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_36 = 8'h24 == result_addr | valid_bits_36; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_37 = 8'h25 == result_addr | valid_bits_37; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_38 = 8'h26 == result_addr | valid_bits_38; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_39 = 8'h27 == result_addr | valid_bits_39; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_40 = 8'h28 == result_addr | valid_bits_40; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_41 = 8'h29 == result_addr | valid_bits_41; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_42 = 8'h2a == result_addr | valid_bits_42; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_43 = 8'h2b == result_addr | valid_bits_43; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_44 = 8'h2c == result_addr | valid_bits_44; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_45 = 8'h2d == result_addr | valid_bits_45; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_46 = 8'h2e == result_addr | valid_bits_46; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_47 = 8'h2f == result_addr | valid_bits_47; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_48 = 8'h30 == result_addr | valid_bits_48; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_49 = 8'h31 == result_addr | valid_bits_49; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_50 = 8'h32 == result_addr | valid_bits_50; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_51 = 8'h33 == result_addr | valid_bits_51; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_52 = 8'h34 == result_addr | valid_bits_52; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_53 = 8'h35 == result_addr | valid_bits_53; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_54 = 8'h36 == result_addr | valid_bits_54; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_55 = 8'h37 == result_addr | valid_bits_55; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_56 = 8'h38 == result_addr | valid_bits_56; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_57 = 8'h39 == result_addr | valid_bits_57; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_58 = 8'h3a == result_addr | valid_bits_58; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_59 = 8'h3b == result_addr | valid_bits_59; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_60 = 8'h3c == result_addr | valid_bits_60; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_61 = 8'h3d == result_addr | valid_bits_61; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_62 = 8'h3e == result_addr | valid_bits_62; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_63 = 8'h3f == result_addr | valid_bits_63; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_64 = 8'h40 == result_addr | valid_bits_64; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_65 = 8'h41 == result_addr | valid_bits_65; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_66 = 8'h42 == result_addr | valid_bits_66; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_67 = 8'h43 == result_addr | valid_bits_67; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_68 = 8'h44 == result_addr | valid_bits_68; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_69 = 8'h45 == result_addr | valid_bits_69; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_70 = 8'h46 == result_addr | valid_bits_70; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_71 = 8'h47 == result_addr | valid_bits_71; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_72 = 8'h48 == result_addr | valid_bits_72; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_73 = 8'h49 == result_addr | valid_bits_73; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_74 = 8'h4a == result_addr | valid_bits_74; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_75 = 8'h4b == result_addr | valid_bits_75; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_76 = 8'h4c == result_addr | valid_bits_76; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_77 = 8'h4d == result_addr | valid_bits_77; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_78 = 8'h4e == result_addr | valid_bits_78; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_79 = 8'h4f == result_addr | valid_bits_79; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_80 = 8'h50 == result_addr | valid_bits_80; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_81 = 8'h51 == result_addr | valid_bits_81; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_82 = 8'h52 == result_addr | valid_bits_82; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_83 = 8'h53 == result_addr | valid_bits_83; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_84 = 8'h54 == result_addr | valid_bits_84; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_85 = 8'h55 == result_addr | valid_bits_85; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_86 = 8'h56 == result_addr | valid_bits_86; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_87 = 8'h57 == result_addr | valid_bits_87; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_88 = 8'h58 == result_addr | valid_bits_88; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_89 = 8'h59 == result_addr | valid_bits_89; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_90 = 8'h5a == result_addr | valid_bits_90; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_91 = 8'h5b == result_addr | valid_bits_91; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_92 = 8'h5c == result_addr | valid_bits_92; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_93 = 8'h5d == result_addr | valid_bits_93; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_94 = 8'h5e == result_addr | valid_bits_94; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_95 = 8'h5f == result_addr | valid_bits_95; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_96 = 8'h60 == result_addr | valid_bits_96; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_97 = 8'h61 == result_addr | valid_bits_97; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_98 = 8'h62 == result_addr | valid_bits_98; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_99 = 8'h63 == result_addr | valid_bits_99; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_100 = 8'h64 == result_addr | valid_bits_100; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_101 = 8'h65 == result_addr | valid_bits_101; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_102 = 8'h66 == result_addr | valid_bits_102; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_103 = 8'h67 == result_addr | valid_bits_103; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_104 = 8'h68 == result_addr | valid_bits_104; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_105 = 8'h69 == result_addr | valid_bits_105; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_106 = 8'h6a == result_addr | valid_bits_106; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_107 = 8'h6b == result_addr | valid_bits_107; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_108 = 8'h6c == result_addr | valid_bits_108; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_109 = 8'h6d == result_addr | valid_bits_109; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_110 = 8'h6e == result_addr | valid_bits_110; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_111 = 8'h6f == result_addr | valid_bits_111; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_112 = 8'h70 == result_addr | valid_bits_112; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_113 = 8'h71 == result_addr | valid_bits_113; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_114 = 8'h72 == result_addr | valid_bits_114; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_115 = 8'h73 == result_addr | valid_bits_115; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_116 = 8'h74 == result_addr | valid_bits_116; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_117 = 8'h75 == result_addr | valid_bits_117; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_118 = 8'h76 == result_addr | valid_bits_118; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_119 = 8'h77 == result_addr | valid_bits_119; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_120 = 8'h78 == result_addr | valid_bits_120; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_121 = 8'h79 == result_addr | valid_bits_121; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_122 = 8'h7a == result_addr | valid_bits_122; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_123 = 8'h7b == result_addr | valid_bits_123; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_124 = 8'h7c == result_addr | valid_bits_124; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_125 = 8'h7d == result_addr | valid_bits_125; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_126 = 8'h7e == result_addr | valid_bits_126; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_127 = 8'h7f == result_addr | valid_bits_127; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_128 = 8'h80 == result_addr | valid_bits_128; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_129 = 8'h81 == result_addr | valid_bits_129; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_130 = 8'h82 == result_addr | valid_bits_130; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_131 = 8'h83 == result_addr | valid_bits_131; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_132 = 8'h84 == result_addr | valid_bits_132; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_133 = 8'h85 == result_addr | valid_bits_133; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_134 = 8'h86 == result_addr | valid_bits_134; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_135 = 8'h87 == result_addr | valid_bits_135; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_136 = 8'h88 == result_addr | valid_bits_136; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_137 = 8'h89 == result_addr | valid_bits_137; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_138 = 8'h8a == result_addr | valid_bits_138; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_139 = 8'h8b == result_addr | valid_bits_139; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_140 = 8'h8c == result_addr | valid_bits_140; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_141 = 8'h8d == result_addr | valid_bits_141; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_142 = 8'h8e == result_addr | valid_bits_142; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_143 = 8'h8f == result_addr | valid_bits_143; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_144 = 8'h90 == result_addr | valid_bits_144; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_145 = 8'h91 == result_addr | valid_bits_145; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_146 = 8'h92 == result_addr | valid_bits_146; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_147 = 8'h93 == result_addr | valid_bits_147; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_148 = 8'h94 == result_addr | valid_bits_148; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_149 = 8'h95 == result_addr | valid_bits_149; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_150 = 8'h96 == result_addr | valid_bits_150; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_151 = 8'h97 == result_addr | valid_bits_151; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_152 = 8'h98 == result_addr | valid_bits_152; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_153 = 8'h99 == result_addr | valid_bits_153; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_154 = 8'h9a == result_addr | valid_bits_154; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_155 = 8'h9b == result_addr | valid_bits_155; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_156 = 8'h9c == result_addr | valid_bits_156; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_157 = 8'h9d == result_addr | valid_bits_157; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_158 = 8'h9e == result_addr | valid_bits_158; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_159 = 8'h9f == result_addr | valid_bits_159; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_160 = 8'ha0 == result_addr | valid_bits_160; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_161 = 8'ha1 == result_addr | valid_bits_161; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_162 = 8'ha2 == result_addr | valid_bits_162; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_163 = 8'ha3 == result_addr | valid_bits_163; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_164 = 8'ha4 == result_addr | valid_bits_164; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_165 = 8'ha5 == result_addr | valid_bits_165; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_166 = 8'ha6 == result_addr | valid_bits_166; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_167 = 8'ha7 == result_addr | valid_bits_167; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_168 = 8'ha8 == result_addr | valid_bits_168; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_169 = 8'ha9 == result_addr | valid_bits_169; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_170 = 8'haa == result_addr | valid_bits_170; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_171 = 8'hab == result_addr | valid_bits_171; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_172 = 8'hac == result_addr | valid_bits_172; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_173 = 8'had == result_addr | valid_bits_173; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_174 = 8'hae == result_addr | valid_bits_174; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_175 = 8'haf == result_addr | valid_bits_175; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_176 = 8'hb0 == result_addr | valid_bits_176; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_177 = 8'hb1 == result_addr | valid_bits_177; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_178 = 8'hb2 == result_addr | valid_bits_178; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_179 = 8'hb3 == result_addr | valid_bits_179; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_180 = 8'hb4 == result_addr | valid_bits_180; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_181 = 8'hb5 == result_addr | valid_bits_181; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_182 = 8'hb6 == result_addr | valid_bits_182; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_183 = 8'hb7 == result_addr | valid_bits_183; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_184 = 8'hb8 == result_addr | valid_bits_184; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_185 = 8'hb9 == result_addr | valid_bits_185; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_186 = 8'hba == result_addr | valid_bits_186; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_187 = 8'hbb == result_addr | valid_bits_187; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_188 = 8'hbc == result_addr | valid_bits_188; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_189 = 8'hbd == result_addr | valid_bits_189; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_190 = 8'hbe == result_addr | valid_bits_190; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_191 = 8'hbf == result_addr | valid_bits_191; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_192 = 8'hc0 == result_addr | valid_bits_192; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_193 = 8'hc1 == result_addr | valid_bits_193; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_194 = 8'hc2 == result_addr | valid_bits_194; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_195 = 8'hc3 == result_addr | valid_bits_195; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_196 = 8'hc4 == result_addr | valid_bits_196; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_197 = 8'hc5 == result_addr | valid_bits_197; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_198 = 8'hc6 == result_addr | valid_bits_198; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_199 = 8'hc7 == result_addr | valid_bits_199; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_200 = 8'hc8 == result_addr | valid_bits_200; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_201 = 8'hc9 == result_addr | valid_bits_201; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_202 = 8'hca == result_addr | valid_bits_202; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_203 = 8'hcb == result_addr | valid_bits_203; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_204 = 8'hcc == result_addr | valid_bits_204; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_205 = 8'hcd == result_addr | valid_bits_205; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_206 = 8'hce == result_addr | valid_bits_206; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_207 = 8'hcf == result_addr | valid_bits_207; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_208 = 8'hd0 == result_addr | valid_bits_208; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_209 = 8'hd1 == result_addr | valid_bits_209; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_210 = 8'hd2 == result_addr | valid_bits_210; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_211 = 8'hd3 == result_addr | valid_bits_211; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_212 = 8'hd4 == result_addr | valid_bits_212; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_213 = 8'hd5 == result_addr | valid_bits_213; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_214 = 8'hd6 == result_addr | valid_bits_214; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_215 = 8'hd7 == result_addr | valid_bits_215; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_216 = 8'hd8 == result_addr | valid_bits_216; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_217 = 8'hd9 == result_addr | valid_bits_217; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_218 = 8'hda == result_addr | valid_bits_218; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_219 = 8'hdb == result_addr | valid_bits_219; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_220 = 8'hdc == result_addr | valid_bits_220; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_221 = 8'hdd == result_addr | valid_bits_221; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_222 = 8'hde == result_addr | valid_bits_222; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_223 = 8'hdf == result_addr | valid_bits_223; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_224 = 8'he0 == result_addr | valid_bits_224; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_225 = 8'he1 == result_addr | valid_bits_225; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_226 = 8'he2 == result_addr | valid_bits_226; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_227 = 8'he3 == result_addr | valid_bits_227; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_228 = 8'he4 == result_addr | valid_bits_228; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_229 = 8'he5 == result_addr | valid_bits_229; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_230 = 8'he6 == result_addr | valid_bits_230; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_231 = 8'he7 == result_addr | valid_bits_231; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_232 = 8'he8 == result_addr | valid_bits_232; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_233 = 8'he9 == result_addr | valid_bits_233; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_234 = 8'hea == result_addr | valid_bits_234; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_235 = 8'heb == result_addr | valid_bits_235; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_236 = 8'hec == result_addr | valid_bits_236; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_237 = 8'hed == result_addr | valid_bits_237; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_238 = 8'hee == result_addr | valid_bits_238; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_239 = 8'hef == result_addr | valid_bits_239; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_240 = 8'hf0 == result_addr | valid_bits_240; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_241 = 8'hf1 == result_addr | valid_bits_241; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_242 = 8'hf2 == result_addr | valid_bits_242; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_243 = 8'hf3 == result_addr | valid_bits_243; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_244 = 8'hf4 == result_addr | valid_bits_244; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_245 = 8'hf5 == result_addr | valid_bits_245; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_246 = 8'hf6 == result_addr | valid_bits_246; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_247 = 8'hf7 == result_addr | valid_bits_247; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_248 = 8'hf8 == result_addr | valid_bits_248; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_249 = 8'hf9 == result_addr | valid_bits_249; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_250 = 8'hfa == result_addr | valid_bits_250; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_251 = 8'hfb == result_addr | valid_bits_251; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_252 = 8'hfc == result_addr | valid_bits_252; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_253 = 8'hfd == result_addr | valid_bits_253; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_254 = 8'hfe == result_addr | valid_bits_254; // @[fetch.scala 147:27 153:{31,31}]
  wire  _GEN_255 = 8'hff == result_addr | valid_bits_255; // @[fetch.scala 147:27 153:{31,31}]
  wire  _T_1 = ~(counters_MPORT_2_data == 2'h3); // @[fetch.scala 158:14]
  wire  _T_5 = ~(counters_MPORT_5_data == 2'h0); // @[fetch.scala 162:14]
  wire  _GEN_271 = io_branchres_branchTaken & _T_1; // @[fetch.scala 146:21 157:37]
  wire  _GEN_276 = io_branchres_branchTaken ? 1'h0 : 1'h1; // @[fetch.scala 146:21 157:37 162:24]
  wire  _GEN_279 = io_branchres_branchTaken ? 1'h0 : _T_5; // @[fetch.scala 146:21 157:37]
  wire  _GEN_1351 = 8'h1 == btb_addr ? valid_bits_1 : valid_bits_0; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1352 = 8'h2 == btb_addr ? valid_bits_2 : _GEN_1351; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1353 = 8'h3 == btb_addr ? valid_bits_3 : _GEN_1352; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1354 = 8'h4 == btb_addr ? valid_bits_4 : _GEN_1353; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1355 = 8'h5 == btb_addr ? valid_bits_5 : _GEN_1354; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1356 = 8'h6 == btb_addr ? valid_bits_6 : _GEN_1355; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1357 = 8'h7 == btb_addr ? valid_bits_7 : _GEN_1356; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1358 = 8'h8 == btb_addr ? valid_bits_8 : _GEN_1357; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1359 = 8'h9 == btb_addr ? valid_bits_9 : _GEN_1358; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1360 = 8'ha == btb_addr ? valid_bits_10 : _GEN_1359; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1361 = 8'hb == btb_addr ? valid_bits_11 : _GEN_1360; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1362 = 8'hc == btb_addr ? valid_bits_12 : _GEN_1361; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1363 = 8'hd == btb_addr ? valid_bits_13 : _GEN_1362; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1364 = 8'he == btb_addr ? valid_bits_14 : _GEN_1363; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1365 = 8'hf == btb_addr ? valid_bits_15 : _GEN_1364; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1366 = 8'h10 == btb_addr ? valid_bits_16 : _GEN_1365; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1367 = 8'h11 == btb_addr ? valid_bits_17 : _GEN_1366; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1368 = 8'h12 == btb_addr ? valid_bits_18 : _GEN_1367; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1369 = 8'h13 == btb_addr ? valid_bits_19 : _GEN_1368; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1370 = 8'h14 == btb_addr ? valid_bits_20 : _GEN_1369; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1371 = 8'h15 == btb_addr ? valid_bits_21 : _GEN_1370; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1372 = 8'h16 == btb_addr ? valid_bits_22 : _GEN_1371; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1373 = 8'h17 == btb_addr ? valid_bits_23 : _GEN_1372; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1374 = 8'h18 == btb_addr ? valid_bits_24 : _GEN_1373; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1375 = 8'h19 == btb_addr ? valid_bits_25 : _GEN_1374; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1376 = 8'h1a == btb_addr ? valid_bits_26 : _GEN_1375; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1377 = 8'h1b == btb_addr ? valid_bits_27 : _GEN_1376; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1378 = 8'h1c == btb_addr ? valid_bits_28 : _GEN_1377; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1379 = 8'h1d == btb_addr ? valid_bits_29 : _GEN_1378; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1380 = 8'h1e == btb_addr ? valid_bits_30 : _GEN_1379; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1381 = 8'h1f == btb_addr ? valid_bits_31 : _GEN_1380; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1382 = 8'h20 == btb_addr ? valid_bits_32 : _GEN_1381; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1383 = 8'h21 == btb_addr ? valid_bits_33 : _GEN_1382; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1384 = 8'h22 == btb_addr ? valid_bits_34 : _GEN_1383; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1385 = 8'h23 == btb_addr ? valid_bits_35 : _GEN_1384; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1386 = 8'h24 == btb_addr ? valid_bits_36 : _GEN_1385; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1387 = 8'h25 == btb_addr ? valid_bits_37 : _GEN_1386; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1388 = 8'h26 == btb_addr ? valid_bits_38 : _GEN_1387; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1389 = 8'h27 == btb_addr ? valid_bits_39 : _GEN_1388; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1390 = 8'h28 == btb_addr ? valid_bits_40 : _GEN_1389; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1391 = 8'h29 == btb_addr ? valid_bits_41 : _GEN_1390; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1392 = 8'h2a == btb_addr ? valid_bits_42 : _GEN_1391; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1393 = 8'h2b == btb_addr ? valid_bits_43 : _GEN_1392; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1394 = 8'h2c == btb_addr ? valid_bits_44 : _GEN_1393; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1395 = 8'h2d == btb_addr ? valid_bits_45 : _GEN_1394; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1396 = 8'h2e == btb_addr ? valid_bits_46 : _GEN_1395; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1397 = 8'h2f == btb_addr ? valid_bits_47 : _GEN_1396; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1398 = 8'h30 == btb_addr ? valid_bits_48 : _GEN_1397; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1399 = 8'h31 == btb_addr ? valid_bits_49 : _GEN_1398; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1400 = 8'h32 == btb_addr ? valid_bits_50 : _GEN_1399; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1401 = 8'h33 == btb_addr ? valid_bits_51 : _GEN_1400; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1402 = 8'h34 == btb_addr ? valid_bits_52 : _GEN_1401; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1403 = 8'h35 == btb_addr ? valid_bits_53 : _GEN_1402; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1404 = 8'h36 == btb_addr ? valid_bits_54 : _GEN_1403; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1405 = 8'h37 == btb_addr ? valid_bits_55 : _GEN_1404; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1406 = 8'h38 == btb_addr ? valid_bits_56 : _GEN_1405; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1407 = 8'h39 == btb_addr ? valid_bits_57 : _GEN_1406; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1408 = 8'h3a == btb_addr ? valid_bits_58 : _GEN_1407; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1409 = 8'h3b == btb_addr ? valid_bits_59 : _GEN_1408; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1410 = 8'h3c == btb_addr ? valid_bits_60 : _GEN_1409; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1411 = 8'h3d == btb_addr ? valid_bits_61 : _GEN_1410; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1412 = 8'h3e == btb_addr ? valid_bits_62 : _GEN_1411; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1413 = 8'h3f == btb_addr ? valid_bits_63 : _GEN_1412; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1414 = 8'h40 == btb_addr ? valid_bits_64 : _GEN_1413; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1415 = 8'h41 == btb_addr ? valid_bits_65 : _GEN_1414; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1416 = 8'h42 == btb_addr ? valid_bits_66 : _GEN_1415; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1417 = 8'h43 == btb_addr ? valid_bits_67 : _GEN_1416; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1418 = 8'h44 == btb_addr ? valid_bits_68 : _GEN_1417; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1419 = 8'h45 == btb_addr ? valid_bits_69 : _GEN_1418; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1420 = 8'h46 == btb_addr ? valid_bits_70 : _GEN_1419; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1421 = 8'h47 == btb_addr ? valid_bits_71 : _GEN_1420; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1422 = 8'h48 == btb_addr ? valid_bits_72 : _GEN_1421; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1423 = 8'h49 == btb_addr ? valid_bits_73 : _GEN_1422; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1424 = 8'h4a == btb_addr ? valid_bits_74 : _GEN_1423; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1425 = 8'h4b == btb_addr ? valid_bits_75 : _GEN_1424; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1426 = 8'h4c == btb_addr ? valid_bits_76 : _GEN_1425; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1427 = 8'h4d == btb_addr ? valid_bits_77 : _GEN_1426; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1428 = 8'h4e == btb_addr ? valid_bits_78 : _GEN_1427; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1429 = 8'h4f == btb_addr ? valid_bits_79 : _GEN_1428; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1430 = 8'h50 == btb_addr ? valid_bits_80 : _GEN_1429; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1431 = 8'h51 == btb_addr ? valid_bits_81 : _GEN_1430; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1432 = 8'h52 == btb_addr ? valid_bits_82 : _GEN_1431; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1433 = 8'h53 == btb_addr ? valid_bits_83 : _GEN_1432; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1434 = 8'h54 == btb_addr ? valid_bits_84 : _GEN_1433; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1435 = 8'h55 == btb_addr ? valid_bits_85 : _GEN_1434; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1436 = 8'h56 == btb_addr ? valid_bits_86 : _GEN_1435; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1437 = 8'h57 == btb_addr ? valid_bits_87 : _GEN_1436; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1438 = 8'h58 == btb_addr ? valid_bits_88 : _GEN_1437; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1439 = 8'h59 == btb_addr ? valid_bits_89 : _GEN_1438; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1440 = 8'h5a == btb_addr ? valid_bits_90 : _GEN_1439; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1441 = 8'h5b == btb_addr ? valid_bits_91 : _GEN_1440; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1442 = 8'h5c == btb_addr ? valid_bits_92 : _GEN_1441; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1443 = 8'h5d == btb_addr ? valid_bits_93 : _GEN_1442; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1444 = 8'h5e == btb_addr ? valid_bits_94 : _GEN_1443; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1445 = 8'h5f == btb_addr ? valid_bits_95 : _GEN_1444; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1446 = 8'h60 == btb_addr ? valid_bits_96 : _GEN_1445; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1447 = 8'h61 == btb_addr ? valid_bits_97 : _GEN_1446; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1448 = 8'h62 == btb_addr ? valid_bits_98 : _GEN_1447; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1449 = 8'h63 == btb_addr ? valid_bits_99 : _GEN_1448; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1450 = 8'h64 == btb_addr ? valid_bits_100 : _GEN_1449; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1451 = 8'h65 == btb_addr ? valid_bits_101 : _GEN_1450; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1452 = 8'h66 == btb_addr ? valid_bits_102 : _GEN_1451; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1453 = 8'h67 == btb_addr ? valid_bits_103 : _GEN_1452; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1454 = 8'h68 == btb_addr ? valid_bits_104 : _GEN_1453; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1455 = 8'h69 == btb_addr ? valid_bits_105 : _GEN_1454; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1456 = 8'h6a == btb_addr ? valid_bits_106 : _GEN_1455; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1457 = 8'h6b == btb_addr ? valid_bits_107 : _GEN_1456; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1458 = 8'h6c == btb_addr ? valid_bits_108 : _GEN_1457; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1459 = 8'h6d == btb_addr ? valid_bits_109 : _GEN_1458; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1460 = 8'h6e == btb_addr ? valid_bits_110 : _GEN_1459; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1461 = 8'h6f == btb_addr ? valid_bits_111 : _GEN_1460; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1462 = 8'h70 == btb_addr ? valid_bits_112 : _GEN_1461; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1463 = 8'h71 == btb_addr ? valid_bits_113 : _GEN_1462; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1464 = 8'h72 == btb_addr ? valid_bits_114 : _GEN_1463; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1465 = 8'h73 == btb_addr ? valid_bits_115 : _GEN_1464; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1466 = 8'h74 == btb_addr ? valid_bits_116 : _GEN_1465; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1467 = 8'h75 == btb_addr ? valid_bits_117 : _GEN_1466; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1468 = 8'h76 == btb_addr ? valid_bits_118 : _GEN_1467; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1469 = 8'h77 == btb_addr ? valid_bits_119 : _GEN_1468; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1470 = 8'h78 == btb_addr ? valid_bits_120 : _GEN_1469; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1471 = 8'h79 == btb_addr ? valid_bits_121 : _GEN_1470; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1472 = 8'h7a == btb_addr ? valid_bits_122 : _GEN_1471; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1473 = 8'h7b == btb_addr ? valid_bits_123 : _GEN_1472; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1474 = 8'h7c == btb_addr ? valid_bits_124 : _GEN_1473; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1475 = 8'h7d == btb_addr ? valid_bits_125 : _GEN_1474; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1476 = 8'h7e == btb_addr ? valid_bits_126 : _GEN_1475; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1477 = 8'h7f == btb_addr ? valid_bits_127 : _GEN_1476; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1478 = 8'h80 == btb_addr ? valid_bits_128 : _GEN_1477; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1479 = 8'h81 == btb_addr ? valid_bits_129 : _GEN_1478; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1480 = 8'h82 == btb_addr ? valid_bits_130 : _GEN_1479; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1481 = 8'h83 == btb_addr ? valid_bits_131 : _GEN_1480; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1482 = 8'h84 == btb_addr ? valid_bits_132 : _GEN_1481; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1483 = 8'h85 == btb_addr ? valid_bits_133 : _GEN_1482; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1484 = 8'h86 == btb_addr ? valid_bits_134 : _GEN_1483; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1485 = 8'h87 == btb_addr ? valid_bits_135 : _GEN_1484; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1486 = 8'h88 == btb_addr ? valid_bits_136 : _GEN_1485; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1487 = 8'h89 == btb_addr ? valid_bits_137 : _GEN_1486; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1488 = 8'h8a == btb_addr ? valid_bits_138 : _GEN_1487; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1489 = 8'h8b == btb_addr ? valid_bits_139 : _GEN_1488; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1490 = 8'h8c == btb_addr ? valid_bits_140 : _GEN_1489; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1491 = 8'h8d == btb_addr ? valid_bits_141 : _GEN_1490; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1492 = 8'h8e == btb_addr ? valid_bits_142 : _GEN_1491; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1493 = 8'h8f == btb_addr ? valid_bits_143 : _GEN_1492; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1494 = 8'h90 == btb_addr ? valid_bits_144 : _GEN_1493; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1495 = 8'h91 == btb_addr ? valid_bits_145 : _GEN_1494; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1496 = 8'h92 == btb_addr ? valid_bits_146 : _GEN_1495; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1497 = 8'h93 == btb_addr ? valid_bits_147 : _GEN_1496; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1498 = 8'h94 == btb_addr ? valid_bits_148 : _GEN_1497; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1499 = 8'h95 == btb_addr ? valid_bits_149 : _GEN_1498; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1500 = 8'h96 == btb_addr ? valid_bits_150 : _GEN_1499; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1501 = 8'h97 == btb_addr ? valid_bits_151 : _GEN_1500; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1502 = 8'h98 == btb_addr ? valid_bits_152 : _GEN_1501; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1503 = 8'h99 == btb_addr ? valid_bits_153 : _GEN_1502; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1504 = 8'h9a == btb_addr ? valid_bits_154 : _GEN_1503; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1505 = 8'h9b == btb_addr ? valid_bits_155 : _GEN_1504; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1506 = 8'h9c == btb_addr ? valid_bits_156 : _GEN_1505; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1507 = 8'h9d == btb_addr ? valid_bits_157 : _GEN_1506; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1508 = 8'h9e == btb_addr ? valid_bits_158 : _GEN_1507; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1509 = 8'h9f == btb_addr ? valid_bits_159 : _GEN_1508; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1510 = 8'ha0 == btb_addr ? valid_bits_160 : _GEN_1509; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1511 = 8'ha1 == btb_addr ? valid_bits_161 : _GEN_1510; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1512 = 8'ha2 == btb_addr ? valid_bits_162 : _GEN_1511; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1513 = 8'ha3 == btb_addr ? valid_bits_163 : _GEN_1512; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1514 = 8'ha4 == btb_addr ? valid_bits_164 : _GEN_1513; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1515 = 8'ha5 == btb_addr ? valid_bits_165 : _GEN_1514; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1516 = 8'ha6 == btb_addr ? valid_bits_166 : _GEN_1515; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1517 = 8'ha7 == btb_addr ? valid_bits_167 : _GEN_1516; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1518 = 8'ha8 == btb_addr ? valid_bits_168 : _GEN_1517; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1519 = 8'ha9 == btb_addr ? valid_bits_169 : _GEN_1518; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1520 = 8'haa == btb_addr ? valid_bits_170 : _GEN_1519; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1521 = 8'hab == btb_addr ? valid_bits_171 : _GEN_1520; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1522 = 8'hac == btb_addr ? valid_bits_172 : _GEN_1521; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1523 = 8'had == btb_addr ? valid_bits_173 : _GEN_1522; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1524 = 8'hae == btb_addr ? valid_bits_174 : _GEN_1523; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1525 = 8'haf == btb_addr ? valid_bits_175 : _GEN_1524; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1526 = 8'hb0 == btb_addr ? valid_bits_176 : _GEN_1525; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1527 = 8'hb1 == btb_addr ? valid_bits_177 : _GEN_1526; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1528 = 8'hb2 == btb_addr ? valid_bits_178 : _GEN_1527; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1529 = 8'hb3 == btb_addr ? valid_bits_179 : _GEN_1528; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1530 = 8'hb4 == btb_addr ? valid_bits_180 : _GEN_1529; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1531 = 8'hb5 == btb_addr ? valid_bits_181 : _GEN_1530; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1532 = 8'hb6 == btb_addr ? valid_bits_182 : _GEN_1531; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1533 = 8'hb7 == btb_addr ? valid_bits_183 : _GEN_1532; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1534 = 8'hb8 == btb_addr ? valid_bits_184 : _GEN_1533; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1535 = 8'hb9 == btb_addr ? valid_bits_185 : _GEN_1534; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1536 = 8'hba == btb_addr ? valid_bits_186 : _GEN_1535; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1537 = 8'hbb == btb_addr ? valid_bits_187 : _GEN_1536; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1538 = 8'hbc == btb_addr ? valid_bits_188 : _GEN_1537; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1539 = 8'hbd == btb_addr ? valid_bits_189 : _GEN_1538; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1540 = 8'hbe == btb_addr ? valid_bits_190 : _GEN_1539; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1541 = 8'hbf == btb_addr ? valid_bits_191 : _GEN_1540; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1542 = 8'hc0 == btb_addr ? valid_bits_192 : _GEN_1541; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1543 = 8'hc1 == btb_addr ? valid_bits_193 : _GEN_1542; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1544 = 8'hc2 == btb_addr ? valid_bits_194 : _GEN_1543; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1545 = 8'hc3 == btb_addr ? valid_bits_195 : _GEN_1544; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1546 = 8'hc4 == btb_addr ? valid_bits_196 : _GEN_1545; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1547 = 8'hc5 == btb_addr ? valid_bits_197 : _GEN_1546; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1548 = 8'hc6 == btb_addr ? valid_bits_198 : _GEN_1547; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1549 = 8'hc7 == btb_addr ? valid_bits_199 : _GEN_1548; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1550 = 8'hc8 == btb_addr ? valid_bits_200 : _GEN_1549; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1551 = 8'hc9 == btb_addr ? valid_bits_201 : _GEN_1550; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1552 = 8'hca == btb_addr ? valid_bits_202 : _GEN_1551; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1553 = 8'hcb == btb_addr ? valid_bits_203 : _GEN_1552; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1554 = 8'hcc == btb_addr ? valid_bits_204 : _GEN_1553; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1555 = 8'hcd == btb_addr ? valid_bits_205 : _GEN_1554; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1556 = 8'hce == btb_addr ? valid_bits_206 : _GEN_1555; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1557 = 8'hcf == btb_addr ? valid_bits_207 : _GEN_1556; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1558 = 8'hd0 == btb_addr ? valid_bits_208 : _GEN_1557; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1559 = 8'hd1 == btb_addr ? valid_bits_209 : _GEN_1558; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1560 = 8'hd2 == btb_addr ? valid_bits_210 : _GEN_1559; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1561 = 8'hd3 == btb_addr ? valid_bits_211 : _GEN_1560; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1562 = 8'hd4 == btb_addr ? valid_bits_212 : _GEN_1561; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1563 = 8'hd5 == btb_addr ? valid_bits_213 : _GEN_1562; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1564 = 8'hd6 == btb_addr ? valid_bits_214 : _GEN_1563; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1565 = 8'hd7 == btb_addr ? valid_bits_215 : _GEN_1564; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1566 = 8'hd8 == btb_addr ? valid_bits_216 : _GEN_1565; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1567 = 8'hd9 == btb_addr ? valid_bits_217 : _GEN_1566; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1568 = 8'hda == btb_addr ? valid_bits_218 : _GEN_1567; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1569 = 8'hdb == btb_addr ? valid_bits_219 : _GEN_1568; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1570 = 8'hdc == btb_addr ? valid_bits_220 : _GEN_1569; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1571 = 8'hdd == btb_addr ? valid_bits_221 : _GEN_1570; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1572 = 8'hde == btb_addr ? valid_bits_222 : _GEN_1571; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1573 = 8'hdf == btb_addr ? valid_bits_223 : _GEN_1572; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1574 = 8'he0 == btb_addr ? valid_bits_224 : _GEN_1573; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1575 = 8'he1 == btb_addr ? valid_bits_225 : _GEN_1574; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1576 = 8'he2 == btb_addr ? valid_bits_226 : _GEN_1575; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1577 = 8'he3 == btb_addr ? valid_bits_227 : _GEN_1576; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1578 = 8'he4 == btb_addr ? valid_bits_228 : _GEN_1577; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1579 = 8'he5 == btb_addr ? valid_bits_229 : _GEN_1578; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1580 = 8'he6 == btb_addr ? valid_bits_230 : _GEN_1579; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1581 = 8'he7 == btb_addr ? valid_bits_231 : _GEN_1580; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1582 = 8'he8 == btb_addr ? valid_bits_232 : _GEN_1581; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1583 = 8'he9 == btb_addr ? valid_bits_233 : _GEN_1582; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1584 = 8'hea == btb_addr ? valid_bits_234 : _GEN_1583; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1585 = 8'heb == btb_addr ? valid_bits_235 : _GEN_1584; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1586 = 8'hec == btb_addr ? valid_bits_236 : _GEN_1585; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1587 = 8'hed == btb_addr ? valid_bits_237 : _GEN_1586; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1588 = 8'hee == btb_addr ? valid_bits_238 : _GEN_1587; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1589 = 8'hef == btb_addr ? valid_bits_239 : _GEN_1588; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1590 = 8'hf0 == btb_addr ? valid_bits_240 : _GEN_1589; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1591 = 8'hf1 == btb_addr ? valid_bits_241 : _GEN_1590; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1592 = 8'hf2 == btb_addr ? valid_bits_242 : _GEN_1591; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1593 = 8'hf3 == btb_addr ? valid_bits_243 : _GEN_1592; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1594 = 8'hf4 == btb_addr ? valid_bits_244 : _GEN_1593; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1595 = 8'hf5 == btb_addr ? valid_bits_245 : _GEN_1594; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1596 = 8'hf6 == btb_addr ? valid_bits_246 : _GEN_1595; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1597 = 8'hf7 == btb_addr ? valid_bits_247 : _GEN_1596; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1598 = 8'hf8 == btb_addr ? valid_bits_248 : _GEN_1597; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1599 = 8'hf9 == btb_addr ? valid_bits_249 : _GEN_1598; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1600 = 8'hfa == btb_addr ? valid_bits_250 : _GEN_1599; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1601 = 8'hfb == btb_addr ? valid_bits_251 : _GEN_1600; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1602 = 8'hfc == btb_addr ? valid_bits_252 : _GEN_1601; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1603 = 8'hfd == btb_addr ? valid_bits_253 : _GEN_1602; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1604 = 8'hfe == btb_addr ? valid_bits_254 : _GEN_1603; // @[fetch.scala 173:{37,37}]
  wire  _GEN_1605 = 8'hff == btb_addr ? valid_bits_255 : _GEN_1604; // @[fetch.scala 173:{37,37}]
  wire  btb_hit = _GEN_1605 & tag_store_btb_hit_MPORT_data == tag; // @[fetch.scala 173:44]
  wire  prediction = counters_prediction_MPORT_data[1]; // @[fetch.scala 174:47]
  wire [63:0] _io_next_pc_T_2 = io_curr_pc + 64'h4; // @[fetch.scala 179:70]
  wire  _GEN_1606 = correct_history_en ? io_branchres_branchTaken : correct_history_output_0; // @[fetch.scala 184:29 185:39 191:41]
  wire  _GEN_1607 = correct_history_output_1; // @[fetch.scala 184:29 187:41 191:41]
  wire  _GEN_1608 = correct_history_output_2; // @[fetch.scala 184:29 187:41 191:41]
  wire  _GEN_1609 = correct_history_output_3; // @[fetch.scala 184:29 187:41 191:41]
  wire  _GEN_1610 = correct_history_output_4; // @[fetch.scala 184:29 187:41 191:41]
  shiftReg correct_history ( // @[fetch.scala 120:31]
    .clock(correct_history_clock),
    .reset(correct_history_reset),
    .in(correct_history_in),
    .en(correct_history_en),
    .output_0(correct_history_output_0),
    .output_1(correct_history_output_1),
    .output_2(correct_history_output_2),
    .output_3(correct_history_output_3),
    .output_4(correct_history_output_4)
  );
  updateShiftReg predicted_history ( // @[fetch.scala 121:33]
    .clock(predicted_history_clock),
    .reset(predicted_history_reset),
    .in(predicted_history_in),
    .en(predicted_history_en),
    .output_0(predicted_history_output_0),
    .output_1(predicted_history_output_1),
    .output_2(predicted_history_output_2),
    .output_3(predicted_history_output_3),
    .output_4(predicted_history_output_4),
    .updateVals_0(predicted_history_updateVals_0),
    .updateVals_1(predicted_history_updateVals_1),
    .updateVals_2(predicted_history_updateVals_2),
    .updateVals_3(predicted_history_updateVals_3),
    .updateVals_4(predicted_history_updateVals_4),
    .update(predicted_history_update)
  );
  assign btb_io_next_pc_MPORT_en = 1'h1;
  assign btb_io_next_pc_MPORT_addr = io_curr_pc[9:2];
  assign btb_io_next_pc_MPORT_data = btb[btb_io_next_pc_MPORT_addr]; // @[fetch.scala 145:16]
  assign btb_MPORT_1_data = io_branchres_pcAfterBrnach;
  assign btb_MPORT_1_addr = io_branchres_pc[9:2];
  assign btb_MPORT_1_mask = 1'h1;
  assign btb_MPORT_1_en = io_branchres_fired;
  assign counters_MPORT_2_en = io_branchres_fired & io_branchres_branchTaken;
  assign counters_MPORT_2_addr = {io_branchres_pc[7:2],_counterIndex_train_T_15};
  assign counters_MPORT_2_data = counters[counters_MPORT_2_addr]; // @[fetch.scala 146:21]
  assign counters_MPORT_4_en = io_branchres_fired & _GEN_271;
  assign counters_MPORT_4_addr = {io_branchres_pc[7:2],_counterIndex_train_T_15};
  assign counters_MPORT_4_data = counters[counters_MPORT_4_addr]; // @[fetch.scala 146:21]
  assign counters_MPORT_5_en = io_branchres_fired & _GEN_276;
  assign counters_MPORT_5_addr = {io_branchres_pc[7:2],_counterIndex_train_T_15};
  assign counters_MPORT_5_data = counters[counters_MPORT_5_addr]; // @[fetch.scala 146:21]
  assign counters_MPORT_7_en = io_branchres_fired & _GEN_279;
  assign counters_MPORT_7_addr = {io_branchres_pc[7:2],_counterIndex_train_T_15};
  assign counters_MPORT_7_data = counters[counters_MPORT_7_addr]; // @[fetch.scala 146:21]
  assign counters_prediction_MPORT_en = 1'h1;
  assign counters_prediction_MPORT_addr = {io_curr_pc[7:2],_counterIndex_pred_T_15};
  assign counters_prediction_MPORT_data = counters[counters_prediction_MPORT_addr]; // @[fetch.scala 146:21]
  assign counters_MPORT_3_data = counters_MPORT_4_data + 2'h1;
  assign counters_MPORT_3_addr = {io_branchres_pc[7:2],_counterIndex_train_T_15};
  assign counters_MPORT_3_mask = 1'h1;
  assign counters_MPORT_3_en = io_branchres_fired & _GEN_271;
  assign counters_MPORT_6_data = counters_MPORT_7_data - 2'h1;
  assign counters_MPORT_6_addr = {io_branchres_pc[7:2],_counterIndex_train_T_15};
  assign counters_MPORT_6_mask = 1'h1;
  assign counters_MPORT_6_en = io_branchres_fired & _GEN_279;
  assign tag_store_btb_hit_MPORT_en = 1'h1;
  assign tag_store_btb_hit_MPORT_addr = io_curr_pc[9:2];
  assign tag_store_btb_hit_MPORT_data = tag_store[tag_store_btb_hit_MPORT_addr]; // @[fetch.scala 148:22]
  assign tag_store_MPORT_data = io_branchres_pc[63:10];
  assign tag_store_MPORT_addr = io_branchres_pc[9:2];
  assign tag_store_MPORT_mask = 1'h1;
  assign tag_store_MPORT_en = io_branchres_fired;
  assign io_next_pc = btb_hit & prediction ? btb_io_next_pc_MPORT_data : _io_next_pc_T_2; // @[fetch.scala 179:20]
  assign correct_history_clock = clock;
  assign correct_history_reset = reset;
  assign correct_history_in = io_branchres_branchTaken; // @[fetch.scala 123:22]
  assign correct_history_en = io_branchres_fired; // @[fetch.scala 122:44]
  assign predicted_history_clock = clock;
  assign predicted_history_reset = reset;
  assign predicted_history_in = counters_prediction_MPORT_data[1]; // @[fetch.scala 174:47]
  assign predicted_history_en = ~mispredicted & btb_hit & requestSent; // @[fetch.scala 176:52]
  assign predicted_history_updateVals_0 = mispredicted ? _GEN_1606 : correct_history_output_0; // @[fetch.scala 182:22 126:37]
  assign predicted_history_updateVals_1 = mispredicted ? _GEN_1607 : correct_history_output_1; // @[fetch.scala 182:22 126:37]
  assign predicted_history_updateVals_2 = mispredicted ? _GEN_1608 : correct_history_output_2; // @[fetch.scala 182:22 126:37]
  assign predicted_history_updateVals_3 = mispredicted ? _GEN_1609 : correct_history_output_3; // @[fetch.scala 182:22 126:37]
  assign predicted_history_updateVals_4 = mispredicted ? _GEN_1610 : correct_history_output_4; // @[fetch.scala 182:22 126:37]
  assign predicted_history_update = mispredicted; // @[fetch.scala 182:22 183:30 195:30]
  always @(posedge clock) begin
    if (btb_MPORT_1_en & btb_MPORT_1_mask) begin
      btb[btb_MPORT_1_addr] <= btb_MPORT_1_data; // @[fetch.scala 145:16]
    end
    if (counters_MPORT_3_en & counters_MPORT_3_mask) begin
      counters[counters_MPORT_3_addr] <= counters_MPORT_3_data; // @[fetch.scala 146:21]
    end
    if (counters_MPORT_6_en & counters_MPORT_6_mask) begin
      counters[counters_MPORT_6_addr] <= counters_MPORT_6_data; // @[fetch.scala 146:21]
    end
    if (tag_store_MPORT_en & tag_store_MPORT_mask) begin
      tag_store[tag_store_MPORT_addr] <= tag_store_MPORT_data; // @[fetch.scala 148:22]
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_0 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_0 <= _GEN_0;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_1 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_1 <= _GEN_1;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_2 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_2 <= _GEN_2;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_3 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_3 <= _GEN_3;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_4 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_4 <= _GEN_4;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_5 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_5 <= _GEN_5;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_6 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_6 <= _GEN_6;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_7 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_7 <= _GEN_7;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_8 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_8 <= _GEN_8;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_9 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_9 <= _GEN_9;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_10 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_10 <= _GEN_10;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_11 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_11 <= _GEN_11;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_12 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_12 <= _GEN_12;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_13 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_13 <= _GEN_13;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_14 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_14 <= _GEN_14;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_15 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_15 <= _GEN_15;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_16 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_16 <= _GEN_16;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_17 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_17 <= _GEN_17;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_18 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_18 <= _GEN_18;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_19 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_19 <= _GEN_19;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_20 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_20 <= _GEN_20;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_21 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_21 <= _GEN_21;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_22 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_22 <= _GEN_22;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_23 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_23 <= _GEN_23;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_24 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_24 <= _GEN_24;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_25 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_25 <= _GEN_25;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_26 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_26 <= _GEN_26;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_27 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_27 <= _GEN_27;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_28 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_28 <= _GEN_28;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_29 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_29 <= _GEN_29;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_30 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_30 <= _GEN_30;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_31 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_31 <= _GEN_31;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_32 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_32 <= _GEN_32;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_33 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_33 <= _GEN_33;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_34 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_34 <= _GEN_34;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_35 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_35 <= _GEN_35;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_36 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_36 <= _GEN_36;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_37 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_37 <= _GEN_37;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_38 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_38 <= _GEN_38;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_39 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_39 <= _GEN_39;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_40 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_40 <= _GEN_40;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_41 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_41 <= _GEN_41;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_42 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_42 <= _GEN_42;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_43 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_43 <= _GEN_43;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_44 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_44 <= _GEN_44;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_45 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_45 <= _GEN_45;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_46 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_46 <= _GEN_46;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_47 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_47 <= _GEN_47;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_48 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_48 <= _GEN_48;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_49 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_49 <= _GEN_49;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_50 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_50 <= _GEN_50;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_51 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_51 <= _GEN_51;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_52 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_52 <= _GEN_52;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_53 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_53 <= _GEN_53;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_54 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_54 <= _GEN_54;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_55 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_55 <= _GEN_55;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_56 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_56 <= _GEN_56;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_57 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_57 <= _GEN_57;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_58 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_58 <= _GEN_58;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_59 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_59 <= _GEN_59;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_60 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_60 <= _GEN_60;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_61 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_61 <= _GEN_61;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_62 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_62 <= _GEN_62;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_63 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_63 <= _GEN_63;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_64 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_64 <= _GEN_64;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_65 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_65 <= _GEN_65;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_66 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_66 <= _GEN_66;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_67 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_67 <= _GEN_67;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_68 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_68 <= _GEN_68;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_69 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_69 <= _GEN_69;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_70 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_70 <= _GEN_70;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_71 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_71 <= _GEN_71;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_72 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_72 <= _GEN_72;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_73 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_73 <= _GEN_73;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_74 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_74 <= _GEN_74;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_75 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_75 <= _GEN_75;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_76 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_76 <= _GEN_76;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_77 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_77 <= _GEN_77;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_78 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_78 <= _GEN_78;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_79 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_79 <= _GEN_79;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_80 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_80 <= _GEN_80;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_81 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_81 <= _GEN_81;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_82 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_82 <= _GEN_82;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_83 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_83 <= _GEN_83;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_84 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_84 <= _GEN_84;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_85 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_85 <= _GEN_85;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_86 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_86 <= _GEN_86;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_87 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_87 <= _GEN_87;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_88 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_88 <= _GEN_88;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_89 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_89 <= _GEN_89;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_90 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_90 <= _GEN_90;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_91 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_91 <= _GEN_91;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_92 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_92 <= _GEN_92;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_93 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_93 <= _GEN_93;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_94 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_94 <= _GEN_94;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_95 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_95 <= _GEN_95;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_96 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_96 <= _GEN_96;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_97 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_97 <= _GEN_97;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_98 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_98 <= _GEN_98;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_99 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_99 <= _GEN_99;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_100 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_100 <= _GEN_100;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_101 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_101 <= _GEN_101;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_102 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_102 <= _GEN_102;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_103 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_103 <= _GEN_103;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_104 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_104 <= _GEN_104;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_105 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_105 <= _GEN_105;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_106 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_106 <= _GEN_106;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_107 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_107 <= _GEN_107;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_108 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_108 <= _GEN_108;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_109 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_109 <= _GEN_109;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_110 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_110 <= _GEN_110;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_111 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_111 <= _GEN_111;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_112 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_112 <= _GEN_112;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_113 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_113 <= _GEN_113;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_114 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_114 <= _GEN_114;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_115 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_115 <= _GEN_115;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_116 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_116 <= _GEN_116;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_117 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_117 <= _GEN_117;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_118 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_118 <= _GEN_118;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_119 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_119 <= _GEN_119;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_120 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_120 <= _GEN_120;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_121 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_121 <= _GEN_121;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_122 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_122 <= _GEN_122;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_123 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_123 <= _GEN_123;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_124 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_124 <= _GEN_124;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_125 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_125 <= _GEN_125;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_126 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_126 <= _GEN_126;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_127 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_127 <= _GEN_127;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_128 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_128 <= _GEN_128;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_129 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_129 <= _GEN_129;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_130 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_130 <= _GEN_130;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_131 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_131 <= _GEN_131;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_132 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_132 <= _GEN_132;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_133 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_133 <= _GEN_133;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_134 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_134 <= _GEN_134;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_135 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_135 <= _GEN_135;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_136 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_136 <= _GEN_136;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_137 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_137 <= _GEN_137;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_138 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_138 <= _GEN_138;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_139 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_139 <= _GEN_139;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_140 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_140 <= _GEN_140;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_141 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_141 <= _GEN_141;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_142 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_142 <= _GEN_142;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_143 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_143 <= _GEN_143;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_144 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_144 <= _GEN_144;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_145 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_145 <= _GEN_145;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_146 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_146 <= _GEN_146;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_147 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_147 <= _GEN_147;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_148 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_148 <= _GEN_148;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_149 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_149 <= _GEN_149;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_150 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_150 <= _GEN_150;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_151 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_151 <= _GEN_151;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_152 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_152 <= _GEN_152;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_153 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_153 <= _GEN_153;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_154 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_154 <= _GEN_154;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_155 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_155 <= _GEN_155;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_156 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_156 <= _GEN_156;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_157 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_157 <= _GEN_157;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_158 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_158 <= _GEN_158;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_159 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_159 <= _GEN_159;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_160 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_160 <= _GEN_160;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_161 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_161 <= _GEN_161;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_162 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_162 <= _GEN_162;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_163 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_163 <= _GEN_163;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_164 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_164 <= _GEN_164;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_165 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_165 <= _GEN_165;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_166 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_166 <= _GEN_166;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_167 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_167 <= _GEN_167;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_168 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_168 <= _GEN_168;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_169 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_169 <= _GEN_169;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_170 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_170 <= _GEN_170;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_171 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_171 <= _GEN_171;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_172 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_172 <= _GEN_172;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_173 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_173 <= _GEN_173;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_174 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_174 <= _GEN_174;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_175 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_175 <= _GEN_175;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_176 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_176 <= _GEN_176;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_177 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_177 <= _GEN_177;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_178 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_178 <= _GEN_178;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_179 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_179 <= _GEN_179;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_180 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_180 <= _GEN_180;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_181 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_181 <= _GEN_181;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_182 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_182 <= _GEN_182;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_183 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_183 <= _GEN_183;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_184 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_184 <= _GEN_184;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_185 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_185 <= _GEN_185;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_186 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_186 <= _GEN_186;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_187 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_187 <= _GEN_187;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_188 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_188 <= _GEN_188;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_189 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_189 <= _GEN_189;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_190 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_190 <= _GEN_190;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_191 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_191 <= _GEN_191;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_192 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_192 <= _GEN_192;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_193 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_193 <= _GEN_193;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_194 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_194 <= _GEN_194;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_195 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_195 <= _GEN_195;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_196 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_196 <= _GEN_196;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_197 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_197 <= _GEN_197;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_198 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_198 <= _GEN_198;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_199 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_199 <= _GEN_199;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_200 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_200 <= _GEN_200;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_201 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_201 <= _GEN_201;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_202 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_202 <= _GEN_202;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_203 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_203 <= _GEN_203;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_204 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_204 <= _GEN_204;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_205 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_205 <= _GEN_205;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_206 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_206 <= _GEN_206;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_207 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_207 <= _GEN_207;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_208 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_208 <= _GEN_208;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_209 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_209 <= _GEN_209;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_210 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_210 <= _GEN_210;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_211 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_211 <= _GEN_211;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_212 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_212 <= _GEN_212;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_213 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_213 <= _GEN_213;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_214 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_214 <= _GEN_214;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_215 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_215 <= _GEN_215;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_216 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_216 <= _GEN_216;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_217 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_217 <= _GEN_217;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_218 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_218 <= _GEN_218;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_219 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_219 <= _GEN_219;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_220 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_220 <= _GEN_220;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_221 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_221 <= _GEN_221;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_222 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_222 <= _GEN_222;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_223 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_223 <= _GEN_223;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_224 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_224 <= _GEN_224;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_225 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_225 <= _GEN_225;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_226 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_226 <= _GEN_226;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_227 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_227 <= _GEN_227;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_228 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_228 <= _GEN_228;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_229 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_229 <= _GEN_229;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_230 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_230 <= _GEN_230;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_231 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_231 <= _GEN_231;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_232 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_232 <= _GEN_232;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_233 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_233 <= _GEN_233;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_234 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_234 <= _GEN_234;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_235 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_235 <= _GEN_235;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_236 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_236 <= _GEN_236;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_237 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_237 <= _GEN_237;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_238 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_238 <= _GEN_238;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_239 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_239 <= _GEN_239;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_240 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_240 <= _GEN_240;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_241 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_241 <= _GEN_241;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_242 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_242 <= _GEN_242;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_243 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_243 <= _GEN_243;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_244 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_244 <= _GEN_244;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_245 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_245 <= _GEN_245;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_246 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_246 <= _GEN_246;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_247 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_247 <= _GEN_247;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_248 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_248 <= _GEN_248;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_249 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_249 <= _GEN_249;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_250 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_250 <= _GEN_250;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_251 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_251 <= _GEN_251;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_252 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_252 <= _GEN_252;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_253 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_253 <= _GEN_253;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_254 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_254 <= _GEN_254;
    end
    if (reset) begin // @[fetch.scala 147:27]
      valid_bits_255 <= 1'h0; // @[fetch.scala 147:27]
    end else if (io_branchres_fired) begin // @[fetch.scala 151:27]
      valid_bits_255 <= _GEN_255;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    btb[initvar] = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    counters[initvar] = _RAND_1[1:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    tag_store[initvar] = _RAND_2[53:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  valid_bits_0 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  valid_bits_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  valid_bits_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  valid_bits_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  valid_bits_4 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  valid_bits_5 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  valid_bits_6 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  valid_bits_7 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  valid_bits_8 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  valid_bits_9 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  valid_bits_10 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  valid_bits_11 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  valid_bits_12 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  valid_bits_13 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  valid_bits_14 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  valid_bits_15 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  valid_bits_16 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  valid_bits_17 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  valid_bits_18 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  valid_bits_19 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  valid_bits_20 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  valid_bits_21 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  valid_bits_22 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  valid_bits_23 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  valid_bits_24 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  valid_bits_25 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  valid_bits_26 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  valid_bits_27 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  valid_bits_28 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  valid_bits_29 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  valid_bits_30 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  valid_bits_31 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  valid_bits_32 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  valid_bits_33 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  valid_bits_34 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  valid_bits_35 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  valid_bits_36 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  valid_bits_37 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  valid_bits_38 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  valid_bits_39 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  valid_bits_40 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  valid_bits_41 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  valid_bits_42 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  valid_bits_43 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  valid_bits_44 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  valid_bits_45 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  valid_bits_46 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  valid_bits_47 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  valid_bits_48 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  valid_bits_49 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  valid_bits_50 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  valid_bits_51 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  valid_bits_52 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  valid_bits_53 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  valid_bits_54 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  valid_bits_55 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  valid_bits_56 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  valid_bits_57 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  valid_bits_58 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  valid_bits_59 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  valid_bits_60 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  valid_bits_61 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  valid_bits_62 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  valid_bits_63 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  valid_bits_64 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  valid_bits_65 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  valid_bits_66 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  valid_bits_67 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  valid_bits_68 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  valid_bits_69 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  valid_bits_70 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  valid_bits_71 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  valid_bits_72 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  valid_bits_73 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  valid_bits_74 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  valid_bits_75 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  valid_bits_76 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  valid_bits_77 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  valid_bits_78 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  valid_bits_79 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  valid_bits_80 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  valid_bits_81 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  valid_bits_82 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  valid_bits_83 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  valid_bits_84 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  valid_bits_85 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  valid_bits_86 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  valid_bits_87 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  valid_bits_88 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  valid_bits_89 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  valid_bits_90 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  valid_bits_91 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  valid_bits_92 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  valid_bits_93 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  valid_bits_94 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  valid_bits_95 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  valid_bits_96 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  valid_bits_97 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  valid_bits_98 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  valid_bits_99 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  valid_bits_100 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  valid_bits_101 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  valid_bits_102 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  valid_bits_103 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  valid_bits_104 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  valid_bits_105 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  valid_bits_106 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  valid_bits_107 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  valid_bits_108 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  valid_bits_109 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  valid_bits_110 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  valid_bits_111 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  valid_bits_112 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  valid_bits_113 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  valid_bits_114 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  valid_bits_115 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  valid_bits_116 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  valid_bits_117 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  valid_bits_118 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  valid_bits_119 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  valid_bits_120 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  valid_bits_121 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  valid_bits_122 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  valid_bits_123 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  valid_bits_124 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  valid_bits_125 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  valid_bits_126 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  valid_bits_127 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  valid_bits_128 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  valid_bits_129 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  valid_bits_130 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  valid_bits_131 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  valid_bits_132 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  valid_bits_133 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  valid_bits_134 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  valid_bits_135 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  valid_bits_136 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  valid_bits_137 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  valid_bits_138 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  valid_bits_139 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  valid_bits_140 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  valid_bits_141 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  valid_bits_142 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  valid_bits_143 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  valid_bits_144 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  valid_bits_145 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  valid_bits_146 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  valid_bits_147 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  valid_bits_148 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  valid_bits_149 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  valid_bits_150 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  valid_bits_151 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  valid_bits_152 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  valid_bits_153 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  valid_bits_154 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  valid_bits_155 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  valid_bits_156 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  valid_bits_157 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  valid_bits_158 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  valid_bits_159 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  valid_bits_160 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  valid_bits_161 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  valid_bits_162 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  valid_bits_163 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  valid_bits_164 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  valid_bits_165 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  valid_bits_166 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  valid_bits_167 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  valid_bits_168 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  valid_bits_169 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  valid_bits_170 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  valid_bits_171 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  valid_bits_172 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  valid_bits_173 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  valid_bits_174 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  valid_bits_175 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  valid_bits_176 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  valid_bits_177 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  valid_bits_178 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  valid_bits_179 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  valid_bits_180 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  valid_bits_181 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  valid_bits_182 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  valid_bits_183 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  valid_bits_184 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  valid_bits_185 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  valid_bits_186 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  valid_bits_187 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  valid_bits_188 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  valid_bits_189 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  valid_bits_190 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  valid_bits_191 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  valid_bits_192 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  valid_bits_193 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  valid_bits_194 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  valid_bits_195 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  valid_bits_196 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  valid_bits_197 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  valid_bits_198 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  valid_bits_199 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  valid_bits_200 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  valid_bits_201 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  valid_bits_202 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  valid_bits_203 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  valid_bits_204 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  valid_bits_205 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  valid_bits_206 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  valid_bits_207 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  valid_bits_208 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  valid_bits_209 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  valid_bits_210 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  valid_bits_211 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  valid_bits_212 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  valid_bits_213 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  valid_bits_214 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  valid_bits_215 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  valid_bits_216 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  valid_bits_217 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  valid_bits_218 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  valid_bits_219 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  valid_bits_220 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  valid_bits_221 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  valid_bits_222 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  valid_bits_223 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  valid_bits_224 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  valid_bits_225 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  valid_bits_226 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  valid_bits_227 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  valid_bits_228 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  valid_bits_229 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  valid_bits_230 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  valid_bits_231 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  valid_bits_232 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  valid_bits_233 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  valid_bits_234 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  valid_bits_235 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  valid_bits_236 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  valid_bits_237 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  valid_bits_238 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  valid_bits_239 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  valid_bits_240 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  valid_bits_241 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  valid_bits_242 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  valid_bits_243 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  valid_bits_244 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  valid_bits_245 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  valid_bits_246 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  valid_bits_247 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  valid_bits_248 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  valid_bits_249 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  valid_bits_250 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  valid_bits_251 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  valid_bits_252 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  valid_bits_253 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  valid_bits_254 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  valid_bits_255 = _RAND_258[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module regFifo(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [127:0] io_enq_bits,
  input          io_deq_ready,
  output         io_deq_valid,
  output [127:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] memReg [0:3]; // @[Fifo.scala 21:19]
  wire  memReg_io_deq_bits_MPORT_en; // @[Fifo.scala 21:19]
  wire [1:0] memReg_io_deq_bits_MPORT_addr; // @[Fifo.scala 21:19]
  wire [127:0] memReg_io_deq_bits_MPORT_data; // @[Fifo.scala 21:19]
  wire [127:0] memReg_MPORT_data; // @[Fifo.scala 21:19]
  wire [1:0] memReg_MPORT_addr; // @[Fifo.scala 21:19]
  wire  memReg_MPORT_mask; // @[Fifo.scala 21:19]
  wire  memReg_MPORT_en; // @[Fifo.scala 21:19]
  wire [127:0] memReg_MPORT_1_data; // @[Fifo.scala 21:19]
  wire [1:0] memReg_MPORT_1_addr; // @[Fifo.scala 21:19]
  wire  memReg_MPORT_1_mask; // @[Fifo.scala 21:19]
  wire  memReg_MPORT_1_en; // @[Fifo.scala 21:19]
  reg [1:0] readPtr; // @[Fifo.scala 12:26]
  wire [1:0] _nextVal_T_2 = readPtr + 2'h1; // @[Fifo.scala 13:60]
  wire [1:0] nextRead = readPtr == 2'h3 ? 2'h0 : _nextVal_T_2; // @[Fifo.scala 13:22]
  wire  _T = io_deq_ready & io_deq_valid; // @[Fifo.scala 30:21]
  wire  _T_1 = io_deq_ready & io_deq_valid & io_enq_valid; // @[Fifo.scala 30:37]
  wire  _T_2 = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready; // @[Fifo.scala 30:53]
  wire  _T_3 = io_enq_valid & io_enq_ready; // @[Fifo.scala 34:27]
  wire  _GEN_12 = io_enq_valid & io_enq_ready ? 1'h0 : _T; // @[Fifo.scala 34:44]
  wire  incrRead = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready | _GEN_12; // @[Fifo.scala 30:70 33:14]
  reg [1:0] writePtr; // @[Fifo.scala 12:26]
  wire [1:0] _nextVal_T_5 = writePtr + 2'h1; // @[Fifo.scala 13:60]
  wire [1:0] nextWrite = writePtr == 2'h3 ? 2'h0 : _nextVal_T_5; // @[Fifo.scala 13:22]
  wire  incrWrite = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready | _T_3; // @[Fifo.scala 30:70 32:15]
  reg  emptyReg; // @[Fifo.scala 26:25]
  reg  fullReg; // @[Fifo.scala 27:24]
  wire  _GEN_3 = _T ? nextRead == writePtr : emptyReg; // @[Fifo.scala 39:44 41:14 26:25]
  wire  _GEN_10 = io_enq_valid & io_enq_ready ? 1'h0 : _GEN_3; // @[Fifo.scala 34:44 36:14]
  wire  _GEN_25 = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready ? emptyReg : _GEN_10; // @[Fifo.scala 26:25 30:70]
  assign memReg_io_deq_bits_MPORT_en = 1'h1;
  assign memReg_io_deq_bits_MPORT_addr = readPtr;
  assign memReg_io_deq_bits_MPORT_data = memReg[memReg_io_deq_bits_MPORT_addr]; // @[Fifo.scala 21:19]
  assign memReg_MPORT_data = io_enq_bits;
  assign memReg_MPORT_addr = writePtr;
  assign memReg_MPORT_mask = 1'h1;
  assign memReg_MPORT_en = _T_1 & io_enq_ready;
  assign memReg_MPORT_1_data = io_enq_bits;
  assign memReg_MPORT_1_addr = writePtr;
  assign memReg_MPORT_1_mask = 1'h1;
  assign memReg_MPORT_1_en = _T_2 ? 1'h0 : _T_3;
  assign io_enq_ready = ~fullReg | io_deq_valid & io_deq_ready; // @[Fifo.scala 46:28]
  assign io_deq_valid = ~emptyReg; // @[Fifo.scala 47:19]
  assign io_deq_bits = memReg_io_deq_bits_MPORT_data; // @[Fifo.scala 45:15]
  always @(posedge clock) begin
    if (memReg_MPORT_en & memReg_MPORT_mask) begin
      memReg[memReg_MPORT_addr] <= memReg_MPORT_data; // @[Fifo.scala 21:19]
    end
    if (memReg_MPORT_1_en & memReg_MPORT_1_mask) begin
      memReg[memReg_MPORT_1_addr] <= memReg_MPORT_1_data; // @[Fifo.scala 21:19]
    end
    if (reset) begin // @[Fifo.scala 12:26]
      readPtr <= 2'h0; // @[Fifo.scala 12:26]
    end else if (incrRead) begin // @[Fifo.scala 14:17]
      if (readPtr == 2'h3) begin // @[Fifo.scala 13:22]
        readPtr <= 2'h0;
      end else begin
        readPtr <= _nextVal_T_2;
      end
    end
    if (reset) begin // @[Fifo.scala 12:26]
      writePtr <= 2'h0; // @[Fifo.scala 12:26]
    end else if (incrWrite) begin // @[Fifo.scala 14:17]
      if (writePtr == 2'h3) begin // @[Fifo.scala 13:22]
        writePtr <= 2'h0;
      end else begin
        writePtr <= _nextVal_T_5;
      end
    end
    emptyReg <= reset | _GEN_25; // @[Fifo.scala 26:{25,25}]
    if (reset) begin // @[Fifo.scala 27:24]
      fullReg <= 1'h0; // @[Fifo.scala 27:24]
    end else if (!(io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready)) begin // @[Fifo.scala 30:70]
      if (io_enq_valid & io_enq_ready) begin // @[Fifo.scala 34:44]
        fullReg <= nextWrite == readPtr; // @[Fifo.scala 37:13]
      end else if (_T) begin // @[Fifo.scala 39:44]
        fullReg <= 1'h0; // @[Fifo.scala 40:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    memReg[initvar] = _RAND_0[127:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  readPtr = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  writePtr = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  emptyReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  fullReg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module fetch(
  input         clock,
  input         reset,
  input         cache_req_ready,
  output        cache_req_valid,
  output [63:0] cache_req_bits,
  output        cache_resp_ready,
  input         cache_resp_valid,
  input  [31:0] cache_resp_bits,
  output        toDecode_ready,
  input         toDecode_fired,
  output [63:0] toDecode_pc,
  output [31:0] toDecode_instruction,
  input         toDecode_expected_valid,
  input  [63:0] toDecode_expected_pc,
  input         branchRes_fired,
  input         branchRes_branchTaken,
  input  [63:0] branchRes_pc,
  input  [63:0] branchRes_pcAfterBrnach,
  output        carryOutFence_ready,
  input         carryOutFence_fired,
  output        updateAllCachelines_ready,
  input         updateAllCachelines_fired,
  output        cachelinesUpdatesResp_ready,
  input         cachelinesUpdatesResp_fired
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  predictor_clock; // @[fetch.scala 256:25]
  wire  predictor_reset; // @[fetch.scala 256:25]
  wire  predictor_io_branchres_fired; // @[fetch.scala 256:25]
  wire  predictor_io_branchres_branchTaken; // @[fetch.scala 256:25]
  wire [63:0] predictor_io_branchres_pc; // @[fetch.scala 256:25]
  wire [63:0] predictor_io_branchres_pcAfterBrnach; // @[fetch.scala 256:25]
  wire [63:0] predictor_io_curr_pc; // @[fetch.scala 256:25]
  wire [63:0] predictor_io_next_pc; // @[fetch.scala 256:25]
  wire  predictor_requestSent; // @[fetch.scala 256:25]
  wire  predictor_mispredicted; // @[fetch.scala 256:25]
  wire  PC_fifo_clock; // @[fetch.scala 259:23]
  wire  PC_fifo_reset; // @[fetch.scala 259:23]
  wire  PC_fifo_io_enq_ready; // @[fetch.scala 259:23]
  wire  PC_fifo_io_enq_valid; // @[fetch.scala 259:23]
  wire [127:0] PC_fifo_io_enq_bits; // @[fetch.scala 259:23]
  wire  PC_fifo_io_deq_ready; // @[fetch.scala 259:23]
  wire  PC_fifo_io_deq_valid; // @[fetch.scala 259:23]
  wire [127:0] PC_fifo_io_deq_bits; // @[fetch.scala 259:23]
  reg [63:0] PC; // @[fetch.scala 247:19]
  reg  redirect_bit; // @[fetch.scala 248:28]
  reg  handle_fenceI; // @[fetch.scala 249:29]
  reg  clear_cache_req; // @[fetch.scala 250:31]
  reg  cache_cleared; // @[fetch.scala 251:29]
  reg  fence_pending; // @[fetch.scala 252:29]
  wire  _PC_fifo_io_enq_valid_T = cache_req_valid & cache_req_ready; // @[fetch.scala 263:43]
  wire  is_fenceI = toDecode_instruction[6:2] == 5'h3 & toDecode_instruction[14:13] == 2'h0 & toDecode_fired; // @[fetch.scala 268:102]
  wire  _T_1 = ~handle_fenceI; // @[fetch.scala 272:23]
  wire  _T_2 = ~clear_cache_req; // @[fetch.scala 275:26]
  wire  _T_3 = ~cache_cleared; // @[fetch.scala 275:49]
  wire  _T_5 = ~fence_pending; // @[fetch.scala 275:72]
  wire  redirect = ~(toDecode_expected_pc == toDecode_pc) & toDecode_expected_valid; // @[fetch.scala 302:55]
  wire  _T_19 = ~redirect_bit; // @[fetch.scala 305:20]
  wire  _T_20 = ~redirect_bit & PC_fifo_io_deq_valid; // @[fetch.scala 305:27]
  wire  _T_21 = ~PC_fifo_io_deq_valid; // @[fetch.scala 307:36]
  wire [127:0] _PC_T_1 = PC_fifo_io_deq_bits + 128'h4; // @[fetch.scala 316:31]
  wire [63:0] _GEN_11 = _PC_fifo_io_enq_valid_T ? predictor_io_next_pc : PC; // @[fetch.scala 247:19 317:49 318:8]
  wire [127:0] _GEN_12 = is_fenceI ? _PC_T_1 : {{64'd0}, _GEN_11}; // @[fetch.scala 315:25 316:8]
  wire [127:0] _GEN_13 = redirect_bit ? {{64'd0}, toDecode_expected_pc} : _GEN_12; // @[fetch.scala 313:28 314:8]
  reg  misPredicted; // @[fetch.scala 339:29]
  wire  _GEN_15 = _T_20 & redirect; // @[fetch.scala 340:51 341:18 343:18]
  wire [127:0] _GEN_17 = reset ? 128'h10000000 : _GEN_13; // @[fetch.scala 247:{19,19}]
  gshare_predictor predictor ( // @[fetch.scala 256:25]
    .clock(predictor_clock),
    .reset(predictor_reset),
    .io_branchres_fired(predictor_io_branchres_fired),
    .io_branchres_branchTaken(predictor_io_branchres_branchTaken),
    .io_branchres_pc(predictor_io_branchres_pc),
    .io_branchres_pcAfterBrnach(predictor_io_branchres_pcAfterBrnach),
    .io_curr_pc(predictor_io_curr_pc),
    .io_next_pc(predictor_io_next_pc),
    .requestSent(predictor_requestSent),
    .mispredicted(predictor_mispredicted)
  );
  regFifo PC_fifo ( // @[fetch.scala 259:23]
    .clock(PC_fifo_clock),
    .reset(PC_fifo_reset),
    .io_enq_ready(PC_fifo_io_enq_ready),
    .io_enq_valid(PC_fifo_io_enq_valid),
    .io_enq_bits(PC_fifo_io_enq_bits),
    .io_deq_ready(PC_fifo_io_deq_ready),
    .io_deq_valid(PC_fifo_io_deq_valid),
    .io_deq_bits(PC_fifo_io_deq_bits)
  );
  assign cache_req_valid = _T_19 & PC_fifo_io_enq_ready & ~is_fenceI & _T_1; // @[fetch.scala 323:79]
  assign cache_req_bits = PC; // @[fetch.scala 320:18]
  assign cache_resp_ready = handle_fenceI | (redirect_bit | toDecode_fired) & _T_1; // @[fetch.scala 324:20 347:{30,49}]
  assign toDecode_ready = redirect | redirect_bit | ~cache_resp_valid | _T_21 | handle_fenceI ? 1'h0 : 1'h1; // @[fetch.scala 328:109 329:20 331:20]
  assign toDecode_pc = PC_fifo_io_deq_bits[63:0]; // @[fetch.scala 265:15]
  assign toDecode_instruction = cache_resp_bits; // @[fetch.scala 334:24]
  assign carryOutFence_ready = fence_pending; // @[fetch.scala 292:23]
  assign updateAllCachelines_ready = clear_cache_req; // @[fetch.scala 325:29]
  assign cachelinesUpdatesResp_ready = cache_cleared; // @[fetch.scala 326:31]
  assign predictor_clock = clock;
  assign predictor_reset = reset;
  assign predictor_io_branchres_fired = branchRes_fired; // @[fetch.scala 257:26]
  assign predictor_io_branchres_branchTaken = branchRes_branchTaken; // @[fetch.scala 257:26]
  assign predictor_io_branchres_pc = branchRes_pc; // @[fetch.scala 257:26]
  assign predictor_io_branchres_pcAfterBrnach = branchRes_pcAfterBrnach; // @[fetch.scala 257:26]
  assign predictor_io_curr_pc = PC; // @[fetch.scala 258:24]
  assign predictor_requestSent = cache_req_valid & cache_req_ready; // @[fetch.scala 336:44]
  assign predictor_mispredicted = misPredicted; // @[fetch.scala 346:26]
  assign PC_fifo_clock = clock;
  assign PC_fifo_reset = handle_fenceI | reset; // @[fetch.scala 269:29 270:18]
  assign PC_fifo_io_enq_valid = cache_req_valid & cache_req_ready; // @[fetch.scala 263:43]
  assign PC_fifo_io_enq_bits = {{64'd0}, PC}; // @[fetch.scala 262:23]
  assign PC_fifo_io_deq_ready = cache_resp_valid & cache_resp_ready; // @[fetch.scala 264:44]
  always @(posedge clock) begin
    PC <= _GEN_17[63:0]; // @[fetch.scala 247:{19,19}]
    if (reset) begin // @[fetch.scala 248:28]
      redirect_bit <= 1'h0; // @[fetch.scala 248:28]
    end else if (~redirect_bit & PC_fifo_io_deq_valid) begin // @[fetch.scala 305:50]
      redirect_bit <= redirect; // @[fetch.scala 306:18]
    end else if (~PC_fifo_io_deq_valid) begin // @[fetch.scala 307:44]
      redirect_bit <= 1'h0; // @[fetch.scala 308:18]
    end
    if (reset) begin // @[fetch.scala 249:29]
      handle_fenceI <= 1'h0; // @[fetch.scala 249:29]
    end else if (~handle_fenceI) begin // @[fetch.scala 272:31]
      handle_fenceI <= is_fenceI; // @[fetch.scala 273:19]
    end else if (~clear_cache_req & ~cache_cleared & ~fence_pending) begin // @[fetch.scala 275:79]
      handle_fenceI <= 1'h0; // @[fetch.scala 276:21]
    end
    if (reset) begin // @[fetch.scala 250:31]
      clear_cache_req <= 1'h0; // @[fetch.scala 250:31]
    end else if (_T_2 & _T_1) begin // @[fetch.scala 280:54]
      clear_cache_req <= is_fenceI; // @[fetch.scala 281:21]
    end else if (updateAllCachelines_fired) begin // @[fetch.scala 282:40]
      clear_cache_req <= 1'h0; // @[fetch.scala 283:21]
    end
    if (reset) begin // @[fetch.scala 251:29]
      cache_cleared <= 1'h0; // @[fetch.scala 251:29]
    end else if (_T_3 & _T_1) begin // @[fetch.scala 286:54]
      cache_cleared <= is_fenceI; // @[fetch.scala 287:19]
    end else if (cachelinesUpdatesResp_fired) begin // @[fetch.scala 288:43]
      cache_cleared <= 1'h0; // @[fetch.scala 289:19]
    end
    if (reset) begin // @[fetch.scala 252:29]
      fence_pending <= 1'h0; // @[fetch.scala 252:29]
    end else if (_T_5 & _T_1) begin // @[fetch.scala 294:52]
      fence_pending <= is_fenceI; // @[fetch.scala 295:18]
    end else if (carryOutFence_fired) begin // @[fetch.scala 296:34]
      fence_pending <= 1'h0; // @[fetch.scala 297:18]
    end
    if (reset) begin // @[fetch.scala 339:29]
      misPredicted <= 1'h0; // @[fetch.scala 339:29]
    end else begin
      misPredicted <= _GEN_15;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  PC = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  redirect_bit = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  handle_fenceI = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  clear_cache_req = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  cache_cleared = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  fence_pending = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  misPredicted = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module core_Anon(
  input         clock,
  input         reset,
  output        fromFetch_ready,
  input         fromFetch_fired,
  input  [63:0] fromFetch_pc,
  input  [31:0] fromFetch_instruction,
  output        fromFetch_expected_valid,
  output [63:0] fromFetch_expected_pc,
  output        toExec_ready,
  input         toExec_fired,
  output [31:0] toExec_instruction,
  output [63:0] toExec_pc,
  output [5:0]  toExec_PRFDest,
  output [5:0]  toExec_rs1Addr,
  output        toExec_rs1Ready,
  output [5:0]  toExec_rs2Addr,
  output        toExec_rs2Ready,
  output [3:0]  toExec_branchMask,
  input         writeBackResult_fired,
  input  [31:0] writeBackResult_instruction,
  input  [4:0]  writeBackResult_rdAddr,
  input  [5:0]  writeBackResult_PRFDest,
  input  [63:0] writeBackResult_data,
  input  [5:0]  writeAddrPRF_exec1Addr,
  input  [5:0]  writeAddrPRF_exec2Addr,
  input  [5:0]  writeAddrPRF_exec3Addr,
  input         writeAddrPRF_exec1Valid,
  input         writeAddrPRF_exec2Valid,
  input         writeAddrPRF_exec3Valid,
  output        jumpAddrWrite_ready,
  input         jumpAddrWrite_fired,
  output [5:0]  jumpAddrWrite_PRFDest,
  output [63:0] jumpAddrWrite_linkAddr,
  output        branchPCs_branchPCReady,
  output [63:0] branchPCs_branchPC,
  output        branchPCs_predictedPCReady,
  output [63:0] branchPCs_predictedPC,
  output [3:0]  branchPCs_branchMask,
  input         branchEvalIn_fired,
  input         branchEvalIn_passFail,
  input  [3:0]  branchEvalIn_branchMask,
  input  [63:0] branchEvalIn_targetPC,
  input  [63:0] interruptedPC,
  output        canTakeInterrupt
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [63:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [63:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [63:0] _RAND_854;
  reg [63:0] _RAND_855;
  reg [63:0] _RAND_856;
  reg [63:0] _RAND_857;
  reg [63:0] _RAND_858;
  reg [63:0] _RAND_859;
  reg [63:0] _RAND_860;
  reg [63:0] _RAND_861;
  reg [63:0] _RAND_862;
  reg [63:0] _RAND_863;
  reg [63:0] _RAND_864;
  reg [63:0] _RAND_865;
  reg [63:0] _RAND_866;
  reg [63:0] _RAND_867;
  reg [63:0] _RAND_868;
  reg [63:0] _RAND_869;
  reg [63:0] _RAND_870;
  reg [63:0] _RAND_871;
  reg [63:0] _RAND_872;
  reg [63:0] _RAND_873;
  reg [63:0] _RAND_874;
  reg [63:0] _RAND_875;
  reg [63:0] _RAND_876;
  reg [63:0] _RAND_877;
  reg [63:0] _RAND_878;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] inputBuffer_pc; // @[decode.scala 107:28]
  reg [31:0] inputBuffer_instruction; // @[decode.scala 107:28]
  reg [31:0] outputBuffer_instruction; // @[decode.scala 116:29]
  reg [63:0] outputBuffer_pc; // @[decode.scala 116:29]
  reg [5:0] outputBuffer_PRFDest; // @[decode.scala 116:29]
  reg [5:0] outputBuffer_rs1Addr; // @[decode.scala 116:29]
  reg [5:0] outputBuffer_rs2Addr; // @[decode.scala 116:29]
  reg [63:0] outputBuffer_immediate; // @[decode.scala 116:29]
  reg  branchBuffer_branchPCReady; // @[decode.scala 138:29]
  reg  branchBuffer_predictedPCReady; // @[decode.scala 138:29]
  reg [63:0] branchBuffer_branchPC; // @[decode.scala 138:29]
  reg [63:0] branchBuffer_predictedPC; // @[decode.scala 138:29]
  reg  branchBuffer_branchMask_0; // @[decode.scala 138:29]
  reg  branchBuffer_branchMask_1; // @[decode.scala 138:29]
  reg  branchBuffer_branchMask_2; // @[decode.scala 138:29]
  reg  branchBuffer_branchMask_3; // @[decode.scala 138:29]
  reg [2:0] branchTracker; // @[decode.scala 173:30]
  reg [63:0] expectedPC; // @[decode.scala 183:27]
  reg  stateRegInputBuf; // @[decode.scala 187:34]
  reg  stateRegOutputBuf; // @[decode.scala 188:34]
  reg  stallReg; // @[decode.scala 190:25]
  reg [63:0] ecallPC; // @[decode.scala 191:20]
  reg  PRFValidList_0; // @[decode.scala 193:29]
  reg  PRFValidList_1; // @[decode.scala 193:29]
  reg  PRFValidList_2; // @[decode.scala 193:29]
  reg  PRFValidList_3; // @[decode.scala 193:29]
  reg  PRFValidList_4; // @[decode.scala 193:29]
  reg  PRFValidList_5; // @[decode.scala 193:29]
  reg  PRFValidList_6; // @[decode.scala 193:29]
  reg  PRFValidList_7; // @[decode.scala 193:29]
  reg  PRFValidList_8; // @[decode.scala 193:29]
  reg  PRFValidList_9; // @[decode.scala 193:29]
  reg  PRFValidList_10; // @[decode.scala 193:29]
  reg  PRFValidList_11; // @[decode.scala 193:29]
  reg  PRFValidList_12; // @[decode.scala 193:29]
  reg  PRFValidList_13; // @[decode.scala 193:29]
  reg  PRFValidList_14; // @[decode.scala 193:29]
  reg  PRFValidList_15; // @[decode.scala 193:29]
  reg  PRFValidList_16; // @[decode.scala 193:29]
  reg  PRFValidList_17; // @[decode.scala 193:29]
  reg  PRFValidList_18; // @[decode.scala 193:29]
  reg  PRFValidList_19; // @[decode.scala 193:29]
  reg  PRFValidList_20; // @[decode.scala 193:29]
  reg  PRFValidList_21; // @[decode.scala 193:29]
  reg  PRFValidList_22; // @[decode.scala 193:29]
  reg  PRFValidList_23; // @[decode.scala 193:29]
  reg  PRFValidList_24; // @[decode.scala 193:29]
  reg  PRFValidList_25; // @[decode.scala 193:29]
  reg  PRFValidList_26; // @[decode.scala 193:29]
  reg  PRFValidList_27; // @[decode.scala 193:29]
  reg  PRFValidList_28; // @[decode.scala 193:29]
  reg  PRFValidList_29; // @[decode.scala 193:29]
  reg  PRFValidList_30; // @[decode.scala 193:29]
  reg  PRFValidList_31; // @[decode.scala 193:29]
  reg  PRFValidList_32; // @[decode.scala 193:29]
  reg  PRFValidList_33; // @[decode.scala 193:29]
  reg  PRFValidList_34; // @[decode.scala 193:29]
  reg  PRFValidList_35; // @[decode.scala 193:29]
  reg  PRFValidList_36; // @[decode.scala 193:29]
  reg  PRFValidList_37; // @[decode.scala 193:29]
  reg  PRFValidList_38; // @[decode.scala 193:29]
  reg  PRFValidList_39; // @[decode.scala 193:29]
  reg  PRFValidList_40; // @[decode.scala 193:29]
  reg  PRFValidList_41; // @[decode.scala 193:29]
  reg  PRFValidList_42; // @[decode.scala 193:29]
  reg  PRFValidList_43; // @[decode.scala 193:29]
  reg  PRFValidList_44; // @[decode.scala 193:29]
  reg  PRFValidList_45; // @[decode.scala 193:29]
  reg  PRFValidList_46; // @[decode.scala 193:29]
  reg  PRFValidList_47; // @[decode.scala 193:29]
  reg  PRFValidList_48; // @[decode.scala 193:29]
  reg  PRFValidList_49; // @[decode.scala 193:29]
  reg  PRFValidList_50; // @[decode.scala 193:29]
  reg  PRFValidList_51; // @[decode.scala 193:29]
  reg  PRFValidList_52; // @[decode.scala 193:29]
  reg  PRFValidList_53; // @[decode.scala 193:29]
  reg  PRFValidList_54; // @[decode.scala 193:29]
  reg  PRFValidList_55; // @[decode.scala 193:29]
  reg  PRFValidList_56; // @[decode.scala 193:29]
  reg  PRFValidList_57; // @[decode.scala 193:29]
  reg  PRFValidList_58; // @[decode.scala 193:29]
  reg  PRFValidList_59; // @[decode.scala 193:29]
  reg  PRFValidList_60; // @[decode.scala 193:29]
  reg  PRFValidList_61; // @[decode.scala 193:29]
  reg  PRFValidList_62; // @[decode.scala 193:29]
  reg  PRFValidList_63; // @[decode.scala 193:29]
  wire  _T_424 = ~branchEvalIn_passFail; // @[decode.scala 761:34]
  wire  _T_425 = branchEvalIn_fired & ~branchEvalIn_passFail; // @[decode.scala 761:31]
  wire  _GEN_9096 = branchEvalIn_fired & ~branchEvalIn_passFail ? 1'h0 : 1'h1; // @[decode.scala 761:58 764:26 768:23]
  wire  _GEN_9098 = stallReg ? 1'h0 : _GEN_9096; // @[decode.scala 779:22 780:23]
  wire [4:0] rs1 = inputBuffer_instruction[19:15]; // @[decode.scala 290:16]
  reg [5:0] frontEndRegMap_31; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_30; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_29; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_28; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_27; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_26; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_25; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_24; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_23; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_22; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_21; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_20; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_19; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_18; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_17; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_16; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_15; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_14; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_13; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_12; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_11; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_10; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_9; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_8; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_7; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_6; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_5; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_4; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_3; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_2; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_1; // @[decode.scala 301:36]
  reg [5:0] frontEndRegMap_0; // @[decode.scala 301:36]
  wire [5:0] _GEN_209 = 5'h1 == rs1 ? frontEndRegMap_1 : frontEndRegMap_0; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_210 = 5'h2 == rs1 ? frontEndRegMap_2 : _GEN_209; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_211 = 5'h3 == rs1 ? frontEndRegMap_3 : _GEN_210; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_212 = 5'h4 == rs1 ? frontEndRegMap_4 : _GEN_211; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_213 = 5'h5 == rs1 ? frontEndRegMap_5 : _GEN_212; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_214 = 5'h6 == rs1 ? frontEndRegMap_6 : _GEN_213; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_215 = 5'h7 == rs1 ? frontEndRegMap_7 : _GEN_214; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_216 = 5'h8 == rs1 ? frontEndRegMap_8 : _GEN_215; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_217 = 5'h9 == rs1 ? frontEndRegMap_9 : _GEN_216; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_218 = 5'ha == rs1 ? frontEndRegMap_10 : _GEN_217; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_219 = 5'hb == rs1 ? frontEndRegMap_11 : _GEN_218; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_220 = 5'hc == rs1 ? frontEndRegMap_12 : _GEN_219; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_221 = 5'hd == rs1 ? frontEndRegMap_13 : _GEN_220; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_222 = 5'he == rs1 ? frontEndRegMap_14 : _GEN_221; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_223 = 5'hf == rs1 ? frontEndRegMap_15 : _GEN_222; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_224 = 5'h10 == rs1 ? frontEndRegMap_16 : _GEN_223; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_225 = 5'h11 == rs1 ? frontEndRegMap_17 : _GEN_224; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_226 = 5'h12 == rs1 ? frontEndRegMap_18 : _GEN_225; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_227 = 5'h13 == rs1 ? frontEndRegMap_19 : _GEN_226; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_228 = 5'h14 == rs1 ? frontEndRegMap_20 : _GEN_227; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_229 = 5'h15 == rs1 ? frontEndRegMap_21 : _GEN_228; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_230 = 5'h16 == rs1 ? frontEndRegMap_22 : _GEN_229; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_231 = 5'h17 == rs1 ? frontEndRegMap_23 : _GEN_230; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_232 = 5'h18 == rs1 ? frontEndRegMap_24 : _GEN_231; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_233 = 5'h19 == rs1 ? frontEndRegMap_25 : _GEN_232; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_234 = 5'h1a == rs1 ? frontEndRegMap_26 : _GEN_233; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_235 = 5'h1b == rs1 ? frontEndRegMap_27 : _GEN_234; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_236 = 5'h1c == rs1 ? frontEndRegMap_28 : _GEN_235; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_237 = 5'h1d == rs1 ? frontEndRegMap_29 : _GEN_236; // @[decode.scala 325:{12,12}]
  wire [5:0] _GEN_238 = 5'h1e == rs1 ? frontEndRegMap_30 : _GEN_237; // @[decode.scala 325:{12,12}]
  wire [5:0] rs1Addr = 5'h1f == rs1 ? frontEndRegMap_31 : _GEN_238; // @[decode.scala 325:{12,12}]
  reg  PRFFreeList_0; // @[decode.scala 303:36]
  reg  PRFFreeList_1; // @[decode.scala 303:36]
  reg  PRFFreeList_2; // @[decode.scala 303:36]
  reg  PRFFreeList_3; // @[decode.scala 303:36]
  reg  PRFFreeList_4; // @[decode.scala 303:36]
  reg  PRFFreeList_5; // @[decode.scala 303:36]
  reg  PRFFreeList_6; // @[decode.scala 303:36]
  reg  PRFFreeList_7; // @[decode.scala 303:36]
  reg  PRFFreeList_8; // @[decode.scala 303:36]
  reg  PRFFreeList_9; // @[decode.scala 303:36]
  reg  PRFFreeList_10; // @[decode.scala 303:36]
  reg  PRFFreeList_11; // @[decode.scala 303:36]
  reg  PRFFreeList_12; // @[decode.scala 303:36]
  reg  PRFFreeList_13; // @[decode.scala 303:36]
  reg  PRFFreeList_14; // @[decode.scala 303:36]
  reg  PRFFreeList_15; // @[decode.scala 303:36]
  reg  PRFFreeList_16; // @[decode.scala 303:36]
  reg  PRFFreeList_17; // @[decode.scala 303:36]
  reg  PRFFreeList_18; // @[decode.scala 303:36]
  reg  PRFFreeList_19; // @[decode.scala 303:36]
  reg  PRFFreeList_20; // @[decode.scala 303:36]
  reg  PRFFreeList_21; // @[decode.scala 303:36]
  reg  PRFFreeList_22; // @[decode.scala 303:36]
  reg  PRFFreeList_23; // @[decode.scala 303:36]
  reg  PRFFreeList_24; // @[decode.scala 303:36]
  reg  PRFFreeList_25; // @[decode.scala 303:36]
  reg  PRFFreeList_26; // @[decode.scala 303:36]
  reg  PRFFreeList_27; // @[decode.scala 303:36]
  reg  PRFFreeList_28; // @[decode.scala 303:36]
  reg  PRFFreeList_29; // @[decode.scala 303:36]
  reg  PRFFreeList_30; // @[decode.scala 303:36]
  reg  PRFFreeList_31; // @[decode.scala 303:36]
  reg  PRFFreeList_32; // @[decode.scala 303:36]
  reg  PRFFreeList_33; // @[decode.scala 303:36]
  reg  PRFFreeList_34; // @[decode.scala 303:36]
  reg  PRFFreeList_35; // @[decode.scala 303:36]
  reg  PRFFreeList_36; // @[decode.scala 303:36]
  reg  PRFFreeList_37; // @[decode.scala 303:36]
  reg  PRFFreeList_38; // @[decode.scala 303:36]
  reg  PRFFreeList_39; // @[decode.scala 303:36]
  reg  PRFFreeList_40; // @[decode.scala 303:36]
  reg  PRFFreeList_41; // @[decode.scala 303:36]
  reg  PRFFreeList_42; // @[decode.scala 303:36]
  reg  PRFFreeList_43; // @[decode.scala 303:36]
  reg  PRFFreeList_44; // @[decode.scala 303:36]
  reg  PRFFreeList_45; // @[decode.scala 303:36]
  reg  PRFFreeList_46; // @[decode.scala 303:36]
  reg  PRFFreeList_47; // @[decode.scala 303:36]
  reg  PRFFreeList_48; // @[decode.scala 303:36]
  reg  PRFFreeList_49; // @[decode.scala 303:36]
  reg  PRFFreeList_50; // @[decode.scala 303:36]
  reg  PRFFreeList_51; // @[decode.scala 303:36]
  reg  PRFFreeList_52; // @[decode.scala 303:36]
  reg  PRFFreeList_53; // @[decode.scala 303:36]
  reg  PRFFreeList_54; // @[decode.scala 303:36]
  reg  PRFFreeList_55; // @[decode.scala 303:36]
  reg  PRFFreeList_56; // @[decode.scala 303:36]
  reg  PRFFreeList_57; // @[decode.scala 303:36]
  reg  PRFFreeList_58; // @[decode.scala 303:36]
  reg  PRFFreeList_59; // @[decode.scala 303:36]
  reg  PRFFreeList_60; // @[decode.scala 303:36]
  reg  PRFFreeList_61; // @[decode.scala 303:36]
  reg  PRFFreeList_62; // @[decode.scala 303:36]
  wire [5:0] _freeRegAddr_T = PRFFreeList_62 ? 6'h3e : 6'h3f; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_1 = PRFFreeList_61 ? 6'h3d : _freeRegAddr_T; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_2 = PRFFreeList_60 ? 6'h3c : _freeRegAddr_T_1; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_3 = PRFFreeList_59 ? 6'h3b : _freeRegAddr_T_2; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_4 = PRFFreeList_58 ? 6'h3a : _freeRegAddr_T_3; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_5 = PRFFreeList_57 ? 6'h39 : _freeRegAddr_T_4; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_6 = PRFFreeList_56 ? 6'h38 : _freeRegAddr_T_5; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_7 = PRFFreeList_55 ? 6'h37 : _freeRegAddr_T_6; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_8 = PRFFreeList_54 ? 6'h36 : _freeRegAddr_T_7; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_9 = PRFFreeList_53 ? 6'h35 : _freeRegAddr_T_8; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_10 = PRFFreeList_52 ? 6'h34 : _freeRegAddr_T_9; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_11 = PRFFreeList_51 ? 6'h33 : _freeRegAddr_T_10; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_12 = PRFFreeList_50 ? 6'h32 : _freeRegAddr_T_11; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_13 = PRFFreeList_49 ? 6'h31 : _freeRegAddr_T_12; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_14 = PRFFreeList_48 ? 6'h30 : _freeRegAddr_T_13; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_15 = PRFFreeList_47 ? 6'h2f : _freeRegAddr_T_14; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_16 = PRFFreeList_46 ? 6'h2e : _freeRegAddr_T_15; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_17 = PRFFreeList_45 ? 6'h2d : _freeRegAddr_T_16; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_18 = PRFFreeList_44 ? 6'h2c : _freeRegAddr_T_17; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_19 = PRFFreeList_43 ? 6'h2b : _freeRegAddr_T_18; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_20 = PRFFreeList_42 ? 6'h2a : _freeRegAddr_T_19; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_21 = PRFFreeList_41 ? 6'h29 : _freeRegAddr_T_20; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_22 = PRFFreeList_40 ? 6'h28 : _freeRegAddr_T_21; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_23 = PRFFreeList_39 ? 6'h27 : _freeRegAddr_T_22; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_24 = PRFFreeList_38 ? 6'h26 : _freeRegAddr_T_23; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_25 = PRFFreeList_37 ? 6'h25 : _freeRegAddr_T_24; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_26 = PRFFreeList_36 ? 6'h24 : _freeRegAddr_T_25; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_27 = PRFFreeList_35 ? 6'h23 : _freeRegAddr_T_26; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_28 = PRFFreeList_34 ? 6'h22 : _freeRegAddr_T_27; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_29 = PRFFreeList_33 ? 6'h21 : _freeRegAddr_T_28; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_30 = PRFFreeList_32 ? 6'h20 : _freeRegAddr_T_29; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_31 = PRFFreeList_31 ? 6'h1f : _freeRegAddr_T_30; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_32 = PRFFreeList_30 ? 6'h1e : _freeRegAddr_T_31; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_33 = PRFFreeList_29 ? 6'h1d : _freeRegAddr_T_32; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_34 = PRFFreeList_28 ? 6'h1c : _freeRegAddr_T_33; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_35 = PRFFreeList_27 ? 6'h1b : _freeRegAddr_T_34; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_36 = PRFFreeList_26 ? 6'h1a : _freeRegAddr_T_35; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_37 = PRFFreeList_25 ? 6'h19 : _freeRegAddr_T_36; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_38 = PRFFreeList_24 ? 6'h18 : _freeRegAddr_T_37; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_39 = PRFFreeList_23 ? 6'h17 : _freeRegAddr_T_38; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_40 = PRFFreeList_22 ? 6'h16 : _freeRegAddr_T_39; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_41 = PRFFreeList_21 ? 6'h15 : _freeRegAddr_T_40; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_42 = PRFFreeList_20 ? 6'h14 : _freeRegAddr_T_41; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_43 = PRFFreeList_19 ? 6'h13 : _freeRegAddr_T_42; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_44 = PRFFreeList_18 ? 6'h12 : _freeRegAddr_T_43; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_45 = PRFFreeList_17 ? 6'h11 : _freeRegAddr_T_44; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_46 = PRFFreeList_16 ? 6'h10 : _freeRegAddr_T_45; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_47 = PRFFreeList_15 ? 6'hf : _freeRegAddr_T_46; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_48 = PRFFreeList_14 ? 6'he : _freeRegAddr_T_47; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_49 = PRFFreeList_13 ? 6'hd : _freeRegAddr_T_48; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_50 = PRFFreeList_12 ? 6'hc : _freeRegAddr_T_49; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_51 = PRFFreeList_11 ? 6'hb : _freeRegAddr_T_50; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_52 = PRFFreeList_10 ? 6'ha : _freeRegAddr_T_51; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_53 = PRFFreeList_9 ? 6'h9 : _freeRegAddr_T_52; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_54 = PRFFreeList_8 ? 6'h8 : _freeRegAddr_T_53; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_55 = PRFFreeList_7 ? 6'h7 : _freeRegAddr_T_54; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_56 = PRFFreeList_6 ? 6'h6 : _freeRegAddr_T_55; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_57 = PRFFreeList_5 ? 6'h5 : _freeRegAddr_T_56; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_58 = PRFFreeList_4 ? 6'h4 : _freeRegAddr_T_57; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_59 = PRFFreeList_3 ? 6'h3 : _freeRegAddr_T_58; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_60 = PRFFreeList_2 ? 6'h2 : _freeRegAddr_T_59; // @[Mux.scala 47:70]
  wire [5:0] _freeRegAddr_T_61 = PRFFreeList_1 ? 6'h1 : _freeRegAddr_T_60; // @[Mux.scala 47:70]
  wire [5:0] freeRegAddr = PRFFreeList_0 ? 6'h0 : _freeRegAddr_T_61; // @[Mux.scala 47:70]
  wire  _T_19 = rs1Addr == freeRegAddr; // @[decode.scala 333:16]
  wire [4:0] rs2 = inputBuffer_instruction[24:20]; // @[decode.scala 291:16]
  wire [5:0] _GEN_241 = 5'h1 == rs2 ? frontEndRegMap_1 : frontEndRegMap_0; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_242 = 5'h2 == rs2 ? frontEndRegMap_2 : _GEN_241; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_243 = 5'h3 == rs2 ? frontEndRegMap_3 : _GEN_242; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_244 = 5'h4 == rs2 ? frontEndRegMap_4 : _GEN_243; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_245 = 5'h5 == rs2 ? frontEndRegMap_5 : _GEN_244; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_246 = 5'h6 == rs2 ? frontEndRegMap_6 : _GEN_245; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_247 = 5'h7 == rs2 ? frontEndRegMap_7 : _GEN_246; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_248 = 5'h8 == rs2 ? frontEndRegMap_8 : _GEN_247; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_249 = 5'h9 == rs2 ? frontEndRegMap_9 : _GEN_248; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_250 = 5'ha == rs2 ? frontEndRegMap_10 : _GEN_249; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_251 = 5'hb == rs2 ? frontEndRegMap_11 : _GEN_250; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_252 = 5'hc == rs2 ? frontEndRegMap_12 : _GEN_251; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_253 = 5'hd == rs2 ? frontEndRegMap_13 : _GEN_252; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_254 = 5'he == rs2 ? frontEndRegMap_14 : _GEN_253; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_255 = 5'hf == rs2 ? frontEndRegMap_15 : _GEN_254; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_256 = 5'h10 == rs2 ? frontEndRegMap_16 : _GEN_255; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_257 = 5'h11 == rs2 ? frontEndRegMap_17 : _GEN_256; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_258 = 5'h12 == rs2 ? frontEndRegMap_18 : _GEN_257; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_259 = 5'h13 == rs2 ? frontEndRegMap_19 : _GEN_258; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_260 = 5'h14 == rs2 ? frontEndRegMap_20 : _GEN_259; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_261 = 5'h15 == rs2 ? frontEndRegMap_21 : _GEN_260; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_262 = 5'h16 == rs2 ? frontEndRegMap_22 : _GEN_261; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_263 = 5'h17 == rs2 ? frontEndRegMap_23 : _GEN_262; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_264 = 5'h18 == rs2 ? frontEndRegMap_24 : _GEN_263; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_265 = 5'h19 == rs2 ? frontEndRegMap_25 : _GEN_264; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_266 = 5'h1a == rs2 ? frontEndRegMap_26 : _GEN_265; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_267 = 5'h1b == rs2 ? frontEndRegMap_27 : _GEN_266; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_268 = 5'h1c == rs2 ? frontEndRegMap_28 : _GEN_267; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_269 = 5'h1d == rs2 ? frontEndRegMap_29 : _GEN_268; // @[decode.scala 326:{12,12}]
  wire [5:0] _GEN_270 = 5'h1e == rs2 ? frontEndRegMap_30 : _GEN_269; // @[decode.scala 326:{12,12}]
  wire [5:0] rs2Addr = 5'h1f == rs2 ? frontEndRegMap_31 : _GEN_270; // @[decode.scala 326:{12,12}]
  wire  _T_20 = rs2Addr == freeRegAddr; // @[decode.scala 333:43]
  wire [6:0] opcode = inputBuffer_instruction[6:0]; // @[decode.scala 289:16]
  wire  _T_5 = 7'h6f == opcode; // @[decode.scala 329:69]
  wire  _T_6 = 7'h67 == opcode; // @[decode.scala 329:69]
  wire  _T_7 = 7'h63 == opcode; // @[decode.scala 329:69]
  wire  _T_18 = freeRegAddr == 6'h3f | (7'h6f == opcode | 7'h67 == opcode | 7'h63 == opcode) & (
    branchBuffer_branchMask_0 & branchBuffer_branchMask_1 & branchBuffer_branchMask_2 & branchBuffer_branchMask_3); // @[decode.scala 329:29]
  wire  stall = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr | _T_18; // @[decode.scala 333:60 334:11]
  wire  _T_431 = opcode == 7'h63; // @[decode.scala 790:56]
  wire  _T_432 = opcode == 7'h6f; // @[decode.scala 790:78]
  wire  _T_434 = opcode == 7'h67; // @[decode.scala 790:99]
  wire  _T_435 = opcode == 7'h63 | opcode == 7'h6f | opcode == 7'h67; // @[decode.scala 790:89]
  wire  _T_438 = ~stall & ~(branchEvalIn_fired & (opcode == 7'h63 | opcode == 7'h6f | opcode == 7'h67)); // @[decode.scala 790:21]
  wire  _GEN_9127 = _T_425 ? 1'h0 : toExec_fired; // @[decode.scala 828:58 831:27]
  wire  readyOutputBuf = ~stateRegOutputBuf ? _GEN_9096 : stateRegOutputBuf & _GEN_9127; // @[decode.scala 813:29]
  wire  _GEN_9103 = ~stall & ~(branchEvalIn_fired & (opcode == 7'h63 | opcode == 7'h6f | opcode == 7'h67)) &
    readyOutputBuf; // @[decode.scala 790:114]
  wire  _GEN_9107 = _T_425 ? 1'h0 : _GEN_9103; // @[decode.scala 784:58 787:26]
  wire  _GEN_9109 = stallReg ? 1'h0 : _GEN_9107; // @[decode.scala 804:22 805:23]
  wire  readyInputBuf = ~stateRegInputBuf ? _GEN_9098 : stateRegInputBuf & _GEN_9109; // @[decode.scala 759:28]
  wire  _GEN_0 = fromFetch_instruction[6:0] == 7'h73 | stallReg; // @[decode.scala 199:97 200:16 190:25]
  wire  _GEN_4 = fromFetch_fired & readyInputBuf ? _GEN_0 : stallReg; // @[decode.scala 190:25 196:42]
  wire  _GEN_9106 = _T_425 ? 1'h0 : _T_438; // @[decode.scala 784:58 786:26]
  wire  validInputBuf = ~stateRegInputBuf ? 1'h0 : stateRegInputBuf & _GEN_9106; // @[decode.scala 759:28]
  wire  _T_3 = validInputBuf & readyOutputBuf; // @[decode.scala 206:22]
  wire [2:0] _GEN_188 = 7'hf == opcode ? 3'h6 : 3'h0; // @[utils.scala 10:20 48:17]
  wire [2:0] _GEN_189 = 7'h73 == opcode ? 3'h1 : _GEN_188; // @[utils.scala 10:20 45:17]
  wire [2:0] _GEN_190 = 7'h3b == opcode ? 3'h0 : _GEN_189; // @[utils.scala 10:20 42:17]
  wire [2:0] _GEN_191 = 7'h33 == opcode ? 3'h0 : _GEN_190; // @[utils.scala 10:20 39:17]
  wire [2:0] _GEN_192 = 7'h1b == opcode ? 3'h1 : _GEN_191; // @[utils.scala 10:20 36:17]
  wire [2:0] _GEN_193 = 7'h13 == opcode ? 3'h1 : _GEN_192; // @[utils.scala 10:20 33:17]
  wire [2:0] _GEN_194 = 7'h23 == opcode ? 3'h2 : _GEN_193; // @[utils.scala 10:20 30:17]
  wire [2:0] _GEN_195 = 7'h3 == opcode ? 3'h1 : _GEN_194; // @[utils.scala 10:20 27:17]
  wire [2:0] _GEN_196 = _T_7 ? 3'h3 : _GEN_195; // @[utils.scala 10:20 24:17]
  wire [2:0] _GEN_197 = _T_6 ? 3'h1 : _GEN_196; // @[utils.scala 10:20 21:17]
  wire [2:0] _GEN_198 = _T_5 ? 3'h5 : _GEN_197; // @[utils.scala 10:20 18:17]
  wire [2:0] _GEN_199 = 7'h17 == opcode ? 3'h4 : _GEN_198; // @[utils.scala 10:20 15:17]
  wire [2:0] insType_insType = 7'h37 == opcode ? 3'h4 : _GEN_199; // @[utils.scala 10:20 12:17]
  wire [52:0] _immediate_immediate_T_2 = inputBuffer_instruction[31] ? 53'h1fffffffffffff : 53'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _immediate_immediate_T_4 = {_immediate_immediate_T_2,inputBuffer_instruction[30:20]}; // @[Cat.scala 33:92]
  wire [63:0] _immediate_immediate_T_10 = {_immediate_immediate_T_2,inputBuffer_instruction[30:25],
    inputBuffer_instruction[11:7]}; // @[Cat.scala 33:92]
  wire [64:0] _immediate_immediate_T_17 = {_immediate_immediate_T_2,inputBuffer_instruction[7],inputBuffer_instruction[
    30:25],inputBuffer_instruction[11:8],1'h0}; // @[Cat.scala 33:92]
  wire [31:0] _immediate_immediate_T_20 = inputBuffer_instruction[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _immediate_immediate_T_22 = {_immediate_immediate_T_20,inputBuffer_instruction[31:12],12'h0}; // @[Cat.scala 33:92]
  wire [43:0] _immediate_immediate_T_25 = inputBuffer_instruction[31] ? 44'hfffffffffff : 44'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _immediate_immediate_T_30 = {_immediate_immediate_T_25,inputBuffer_instruction[19:12],
    inputBuffer_instruction[20],inputBuffer_instruction[30:25],inputBuffer_instruction[24:21],1'h0}; // @[Cat.scala 33:92]
  wire [63:0] _GEN_203 = 3'h5 == insType_insType ? _immediate_immediate_T_30 : 64'h0; // @[utils.scala 59:29 73:19]
  wire [63:0] _GEN_204 = 3'h4 == insType_insType ? _immediate_immediate_T_22 : _GEN_203; // @[utils.scala 59:29 70:19]
  wire [64:0] _GEN_205 = 3'h3 == insType_insType ? _immediate_immediate_T_17 : {{1'd0}, _GEN_204}; // @[utils.scala 59:29 67:19]
  wire [64:0] _GEN_206 = 3'h2 == insType_insType ? {{1'd0}, _immediate_immediate_T_10} : _GEN_205; // @[utils.scala 59:29 64:19]
  wire [64:0] _GEN_207 = 3'h1 == insType_insType ? {{1'd0}, _immediate_immediate_T_4} : _GEN_206; // @[utils.scala 59:29 61:19]
  wire [63:0] immediate_immediate = _GEN_207[63:0];
  reg [3:0] branchPCMask; // @[decode.scala 219:29]
  reg  branchReg; // @[decode.scala 220:29]
  reg [63:0] csrReadDataReg; // @[decode.scala 234:31]
  reg [11:0] csrAddrReg; // @[decode.scala 236:27]
  reg [63:0] csrImmReg; // @[decode.scala 237:26]
  wire  _GEN_13 = 6'h1 == outputBuffer_rs1Addr ? PRFValidList_1 : PRFValidList_0; // @[decode.scala 248:{22,22}]
  wire  _GEN_14 = 6'h2 == outputBuffer_rs1Addr ? PRFValidList_2 : _GEN_13; // @[decode.scala 248:{22,22}]
  wire  _GEN_15 = 6'h3 == outputBuffer_rs1Addr ? PRFValidList_3 : _GEN_14; // @[decode.scala 248:{22,22}]
  wire  _GEN_16 = 6'h4 == outputBuffer_rs1Addr ? PRFValidList_4 : _GEN_15; // @[decode.scala 248:{22,22}]
  wire  _GEN_17 = 6'h5 == outputBuffer_rs1Addr ? PRFValidList_5 : _GEN_16; // @[decode.scala 248:{22,22}]
  wire  _GEN_18 = 6'h6 == outputBuffer_rs1Addr ? PRFValidList_6 : _GEN_17; // @[decode.scala 248:{22,22}]
  wire  _GEN_19 = 6'h7 == outputBuffer_rs1Addr ? PRFValidList_7 : _GEN_18; // @[decode.scala 248:{22,22}]
  wire  _GEN_20 = 6'h8 == outputBuffer_rs1Addr ? PRFValidList_8 : _GEN_19; // @[decode.scala 248:{22,22}]
  wire  _GEN_21 = 6'h9 == outputBuffer_rs1Addr ? PRFValidList_9 : _GEN_20; // @[decode.scala 248:{22,22}]
  wire  _GEN_22 = 6'ha == outputBuffer_rs1Addr ? PRFValidList_10 : _GEN_21; // @[decode.scala 248:{22,22}]
  wire  _GEN_23 = 6'hb == outputBuffer_rs1Addr ? PRFValidList_11 : _GEN_22; // @[decode.scala 248:{22,22}]
  wire  _GEN_24 = 6'hc == outputBuffer_rs1Addr ? PRFValidList_12 : _GEN_23; // @[decode.scala 248:{22,22}]
  wire  _GEN_25 = 6'hd == outputBuffer_rs1Addr ? PRFValidList_13 : _GEN_24; // @[decode.scala 248:{22,22}]
  wire  _GEN_26 = 6'he == outputBuffer_rs1Addr ? PRFValidList_14 : _GEN_25; // @[decode.scala 248:{22,22}]
  wire  _GEN_27 = 6'hf == outputBuffer_rs1Addr ? PRFValidList_15 : _GEN_26; // @[decode.scala 248:{22,22}]
  wire  _GEN_28 = 6'h10 == outputBuffer_rs1Addr ? PRFValidList_16 : _GEN_27; // @[decode.scala 248:{22,22}]
  wire  _GEN_29 = 6'h11 == outputBuffer_rs1Addr ? PRFValidList_17 : _GEN_28; // @[decode.scala 248:{22,22}]
  wire  _GEN_30 = 6'h12 == outputBuffer_rs1Addr ? PRFValidList_18 : _GEN_29; // @[decode.scala 248:{22,22}]
  wire  _GEN_31 = 6'h13 == outputBuffer_rs1Addr ? PRFValidList_19 : _GEN_30; // @[decode.scala 248:{22,22}]
  wire  _GEN_32 = 6'h14 == outputBuffer_rs1Addr ? PRFValidList_20 : _GEN_31; // @[decode.scala 248:{22,22}]
  wire  _GEN_33 = 6'h15 == outputBuffer_rs1Addr ? PRFValidList_21 : _GEN_32; // @[decode.scala 248:{22,22}]
  wire  _GEN_34 = 6'h16 == outputBuffer_rs1Addr ? PRFValidList_22 : _GEN_33; // @[decode.scala 248:{22,22}]
  wire  _GEN_35 = 6'h17 == outputBuffer_rs1Addr ? PRFValidList_23 : _GEN_34; // @[decode.scala 248:{22,22}]
  wire  _GEN_36 = 6'h18 == outputBuffer_rs1Addr ? PRFValidList_24 : _GEN_35; // @[decode.scala 248:{22,22}]
  wire  _GEN_37 = 6'h19 == outputBuffer_rs1Addr ? PRFValidList_25 : _GEN_36; // @[decode.scala 248:{22,22}]
  wire  _GEN_38 = 6'h1a == outputBuffer_rs1Addr ? PRFValidList_26 : _GEN_37; // @[decode.scala 248:{22,22}]
  wire  _GEN_39 = 6'h1b == outputBuffer_rs1Addr ? PRFValidList_27 : _GEN_38; // @[decode.scala 248:{22,22}]
  wire  _GEN_40 = 6'h1c == outputBuffer_rs1Addr ? PRFValidList_28 : _GEN_39; // @[decode.scala 248:{22,22}]
  wire  _GEN_41 = 6'h1d == outputBuffer_rs1Addr ? PRFValidList_29 : _GEN_40; // @[decode.scala 248:{22,22}]
  wire  _GEN_42 = 6'h1e == outputBuffer_rs1Addr ? PRFValidList_30 : _GEN_41; // @[decode.scala 248:{22,22}]
  wire  _GEN_43 = 6'h1f == outputBuffer_rs1Addr ? PRFValidList_31 : _GEN_42; // @[decode.scala 248:{22,22}]
  wire  _GEN_44 = 6'h20 == outputBuffer_rs1Addr ? PRFValidList_32 : _GEN_43; // @[decode.scala 248:{22,22}]
  wire  _GEN_45 = 6'h21 == outputBuffer_rs1Addr ? PRFValidList_33 : _GEN_44; // @[decode.scala 248:{22,22}]
  wire  _GEN_46 = 6'h22 == outputBuffer_rs1Addr ? PRFValidList_34 : _GEN_45; // @[decode.scala 248:{22,22}]
  wire  _GEN_47 = 6'h23 == outputBuffer_rs1Addr ? PRFValidList_35 : _GEN_46; // @[decode.scala 248:{22,22}]
  wire  _GEN_48 = 6'h24 == outputBuffer_rs1Addr ? PRFValidList_36 : _GEN_47; // @[decode.scala 248:{22,22}]
  wire  _GEN_49 = 6'h25 == outputBuffer_rs1Addr ? PRFValidList_37 : _GEN_48; // @[decode.scala 248:{22,22}]
  wire  _GEN_50 = 6'h26 == outputBuffer_rs1Addr ? PRFValidList_38 : _GEN_49; // @[decode.scala 248:{22,22}]
  wire  _GEN_51 = 6'h27 == outputBuffer_rs1Addr ? PRFValidList_39 : _GEN_50; // @[decode.scala 248:{22,22}]
  wire  _GEN_52 = 6'h28 == outputBuffer_rs1Addr ? PRFValidList_40 : _GEN_51; // @[decode.scala 248:{22,22}]
  wire  _GEN_53 = 6'h29 == outputBuffer_rs1Addr ? PRFValidList_41 : _GEN_52; // @[decode.scala 248:{22,22}]
  wire  _GEN_54 = 6'h2a == outputBuffer_rs1Addr ? PRFValidList_42 : _GEN_53; // @[decode.scala 248:{22,22}]
  wire  _GEN_55 = 6'h2b == outputBuffer_rs1Addr ? PRFValidList_43 : _GEN_54; // @[decode.scala 248:{22,22}]
  wire  _GEN_56 = 6'h2c == outputBuffer_rs1Addr ? PRFValidList_44 : _GEN_55; // @[decode.scala 248:{22,22}]
  wire  _GEN_57 = 6'h2d == outputBuffer_rs1Addr ? PRFValidList_45 : _GEN_56; // @[decode.scala 248:{22,22}]
  wire  _GEN_58 = 6'h2e == outputBuffer_rs1Addr ? PRFValidList_46 : _GEN_57; // @[decode.scala 248:{22,22}]
  wire  _GEN_59 = 6'h2f == outputBuffer_rs1Addr ? PRFValidList_47 : _GEN_58; // @[decode.scala 248:{22,22}]
  wire  _GEN_60 = 6'h30 == outputBuffer_rs1Addr ? PRFValidList_48 : _GEN_59; // @[decode.scala 248:{22,22}]
  wire  _GEN_61 = 6'h31 == outputBuffer_rs1Addr ? PRFValidList_49 : _GEN_60; // @[decode.scala 248:{22,22}]
  wire  _GEN_62 = 6'h32 == outputBuffer_rs1Addr ? PRFValidList_50 : _GEN_61; // @[decode.scala 248:{22,22}]
  wire  _GEN_63 = 6'h33 == outputBuffer_rs1Addr ? PRFValidList_51 : _GEN_62; // @[decode.scala 248:{22,22}]
  wire  _GEN_64 = 6'h34 == outputBuffer_rs1Addr ? PRFValidList_52 : _GEN_63; // @[decode.scala 248:{22,22}]
  wire  _GEN_65 = 6'h35 == outputBuffer_rs1Addr ? PRFValidList_53 : _GEN_64; // @[decode.scala 248:{22,22}]
  wire  _GEN_66 = 6'h36 == outputBuffer_rs1Addr ? PRFValidList_54 : _GEN_65; // @[decode.scala 248:{22,22}]
  wire  _GEN_67 = 6'h37 == outputBuffer_rs1Addr ? PRFValidList_55 : _GEN_66; // @[decode.scala 248:{22,22}]
  wire  _GEN_68 = 6'h38 == outputBuffer_rs1Addr ? PRFValidList_56 : _GEN_67; // @[decode.scala 248:{22,22}]
  wire  _GEN_69 = 6'h39 == outputBuffer_rs1Addr ? PRFValidList_57 : _GEN_68; // @[decode.scala 248:{22,22}]
  wire  _GEN_70 = 6'h3a == outputBuffer_rs1Addr ? PRFValidList_58 : _GEN_69; // @[decode.scala 248:{22,22}]
  wire  _GEN_71 = 6'h3b == outputBuffer_rs1Addr ? PRFValidList_59 : _GEN_70; // @[decode.scala 248:{22,22}]
  wire  _GEN_72 = 6'h3c == outputBuffer_rs1Addr ? PRFValidList_60 : _GEN_71; // @[decode.scala 248:{22,22}]
  wire  _GEN_73 = 6'h3d == outputBuffer_rs1Addr ? PRFValidList_61 : _GEN_72; // @[decode.scala 248:{22,22}]
  wire  _GEN_74 = 6'h3e == outputBuffer_rs1Addr ? PRFValidList_62 : _GEN_73; // @[decode.scala 248:{22,22}]
  wire [2:0] _GEN_77 = 7'hf == outputBuffer_instruction[6:0] ? 3'h6 : 3'h0; // @[utils.scala 10:20 48:17]
  wire [2:0] _GEN_78 = 7'h73 == outputBuffer_instruction[6:0] ? 3'h1 : _GEN_77; // @[utils.scala 10:20 45:17]
  wire [2:0] _GEN_79 = 7'h3b == outputBuffer_instruction[6:0] ? 3'h0 : _GEN_78; // @[utils.scala 10:20 42:17]
  wire [2:0] _GEN_80 = 7'h33 == outputBuffer_instruction[6:0] ? 3'h0 : _GEN_79; // @[utils.scala 10:20 39:17]
  wire [2:0] _GEN_81 = 7'h1b == outputBuffer_instruction[6:0] ? 3'h1 : _GEN_80; // @[utils.scala 10:20 36:17]
  wire [2:0] _GEN_82 = 7'h13 == outputBuffer_instruction[6:0] ? 3'h1 : _GEN_81; // @[utils.scala 10:20 33:17]
  wire [2:0] _GEN_83 = 7'h23 == outputBuffer_instruction[6:0] ? 3'h2 : _GEN_82; // @[utils.scala 10:20 30:17]
  wire [2:0] _GEN_84 = 7'h3 == outputBuffer_instruction[6:0] ? 3'h1 : _GEN_83; // @[utils.scala 10:20 27:17]
  wire [2:0] _GEN_85 = 7'h63 == outputBuffer_instruction[6:0] ? 3'h3 : _GEN_84; // @[utils.scala 10:20 24:17]
  wire [2:0] _GEN_86 = 7'h67 == outputBuffer_instruction[6:0] ? 3'h1 : _GEN_85; // @[utils.scala 10:20 21:17]
  wire [2:0] _GEN_87 = 7'h6f == outputBuffer_instruction[6:0] ? 3'h5 : _GEN_86; // @[utils.scala 10:20 18:17]
  wire [2:0] _GEN_88 = 7'h17 == outputBuffer_instruction[6:0] ? 3'h4 : _GEN_87; // @[utils.scala 10:20 15:17]
  wire [2:0] toExec_rs2Ready_insType = 7'h37 == outputBuffer_instruction[6:0] ? 3'h4 : _GEN_88; // @[utils.scala 10:20 12:17]
  wire  _GEN_119 = 6'h1 == outputBuffer_rs2Addr ? PRFValidList_1 : PRFValidList_0; // @[decode.scala 250:{60,60}]
  wire  _GEN_120 = 6'h2 == outputBuffer_rs2Addr ? PRFValidList_2 : _GEN_119; // @[decode.scala 250:{60,60}]
  wire  _GEN_121 = 6'h3 == outputBuffer_rs2Addr ? PRFValidList_3 : _GEN_120; // @[decode.scala 250:{60,60}]
  wire  _GEN_122 = 6'h4 == outputBuffer_rs2Addr ? PRFValidList_4 : _GEN_121; // @[decode.scala 250:{60,60}]
  wire  _GEN_123 = 6'h5 == outputBuffer_rs2Addr ? PRFValidList_5 : _GEN_122; // @[decode.scala 250:{60,60}]
  wire  _GEN_124 = 6'h6 == outputBuffer_rs2Addr ? PRFValidList_6 : _GEN_123; // @[decode.scala 250:{60,60}]
  wire  _GEN_125 = 6'h7 == outputBuffer_rs2Addr ? PRFValidList_7 : _GEN_124; // @[decode.scala 250:{60,60}]
  wire  _GEN_126 = 6'h8 == outputBuffer_rs2Addr ? PRFValidList_8 : _GEN_125; // @[decode.scala 250:{60,60}]
  wire  _GEN_127 = 6'h9 == outputBuffer_rs2Addr ? PRFValidList_9 : _GEN_126; // @[decode.scala 250:{60,60}]
  wire  _GEN_128 = 6'ha == outputBuffer_rs2Addr ? PRFValidList_10 : _GEN_127; // @[decode.scala 250:{60,60}]
  wire  _GEN_129 = 6'hb == outputBuffer_rs2Addr ? PRFValidList_11 : _GEN_128; // @[decode.scala 250:{60,60}]
  wire  _GEN_130 = 6'hc == outputBuffer_rs2Addr ? PRFValidList_12 : _GEN_129; // @[decode.scala 250:{60,60}]
  wire  _GEN_131 = 6'hd == outputBuffer_rs2Addr ? PRFValidList_13 : _GEN_130; // @[decode.scala 250:{60,60}]
  wire  _GEN_132 = 6'he == outputBuffer_rs2Addr ? PRFValidList_14 : _GEN_131; // @[decode.scala 250:{60,60}]
  wire  _GEN_133 = 6'hf == outputBuffer_rs2Addr ? PRFValidList_15 : _GEN_132; // @[decode.scala 250:{60,60}]
  wire  _GEN_134 = 6'h10 == outputBuffer_rs2Addr ? PRFValidList_16 : _GEN_133; // @[decode.scala 250:{60,60}]
  wire  _GEN_135 = 6'h11 == outputBuffer_rs2Addr ? PRFValidList_17 : _GEN_134; // @[decode.scala 250:{60,60}]
  wire  _GEN_136 = 6'h12 == outputBuffer_rs2Addr ? PRFValidList_18 : _GEN_135; // @[decode.scala 250:{60,60}]
  wire  _GEN_137 = 6'h13 == outputBuffer_rs2Addr ? PRFValidList_19 : _GEN_136; // @[decode.scala 250:{60,60}]
  wire  _GEN_138 = 6'h14 == outputBuffer_rs2Addr ? PRFValidList_20 : _GEN_137; // @[decode.scala 250:{60,60}]
  wire  _GEN_139 = 6'h15 == outputBuffer_rs2Addr ? PRFValidList_21 : _GEN_138; // @[decode.scala 250:{60,60}]
  wire  _GEN_140 = 6'h16 == outputBuffer_rs2Addr ? PRFValidList_22 : _GEN_139; // @[decode.scala 250:{60,60}]
  wire  _GEN_141 = 6'h17 == outputBuffer_rs2Addr ? PRFValidList_23 : _GEN_140; // @[decode.scala 250:{60,60}]
  wire  _GEN_142 = 6'h18 == outputBuffer_rs2Addr ? PRFValidList_24 : _GEN_141; // @[decode.scala 250:{60,60}]
  wire  _GEN_143 = 6'h19 == outputBuffer_rs2Addr ? PRFValidList_25 : _GEN_142; // @[decode.scala 250:{60,60}]
  wire  _GEN_144 = 6'h1a == outputBuffer_rs2Addr ? PRFValidList_26 : _GEN_143; // @[decode.scala 250:{60,60}]
  wire  _GEN_145 = 6'h1b == outputBuffer_rs2Addr ? PRFValidList_27 : _GEN_144; // @[decode.scala 250:{60,60}]
  wire  _GEN_146 = 6'h1c == outputBuffer_rs2Addr ? PRFValidList_28 : _GEN_145; // @[decode.scala 250:{60,60}]
  wire  _GEN_147 = 6'h1d == outputBuffer_rs2Addr ? PRFValidList_29 : _GEN_146; // @[decode.scala 250:{60,60}]
  wire  _GEN_148 = 6'h1e == outputBuffer_rs2Addr ? PRFValidList_30 : _GEN_147; // @[decode.scala 250:{60,60}]
  wire  _GEN_149 = 6'h1f == outputBuffer_rs2Addr ? PRFValidList_31 : _GEN_148; // @[decode.scala 250:{60,60}]
  wire  _GEN_150 = 6'h20 == outputBuffer_rs2Addr ? PRFValidList_32 : _GEN_149; // @[decode.scala 250:{60,60}]
  wire  _GEN_151 = 6'h21 == outputBuffer_rs2Addr ? PRFValidList_33 : _GEN_150; // @[decode.scala 250:{60,60}]
  wire  _GEN_152 = 6'h22 == outputBuffer_rs2Addr ? PRFValidList_34 : _GEN_151; // @[decode.scala 250:{60,60}]
  wire  _GEN_153 = 6'h23 == outputBuffer_rs2Addr ? PRFValidList_35 : _GEN_152; // @[decode.scala 250:{60,60}]
  wire  _GEN_154 = 6'h24 == outputBuffer_rs2Addr ? PRFValidList_36 : _GEN_153; // @[decode.scala 250:{60,60}]
  wire  _GEN_155 = 6'h25 == outputBuffer_rs2Addr ? PRFValidList_37 : _GEN_154; // @[decode.scala 250:{60,60}]
  wire  _GEN_156 = 6'h26 == outputBuffer_rs2Addr ? PRFValidList_38 : _GEN_155; // @[decode.scala 250:{60,60}]
  wire  _GEN_157 = 6'h27 == outputBuffer_rs2Addr ? PRFValidList_39 : _GEN_156; // @[decode.scala 250:{60,60}]
  wire  _GEN_158 = 6'h28 == outputBuffer_rs2Addr ? PRFValidList_40 : _GEN_157; // @[decode.scala 250:{60,60}]
  wire  _GEN_159 = 6'h29 == outputBuffer_rs2Addr ? PRFValidList_41 : _GEN_158; // @[decode.scala 250:{60,60}]
  wire  _GEN_160 = 6'h2a == outputBuffer_rs2Addr ? PRFValidList_42 : _GEN_159; // @[decode.scala 250:{60,60}]
  wire  _GEN_161 = 6'h2b == outputBuffer_rs2Addr ? PRFValidList_43 : _GEN_160; // @[decode.scala 250:{60,60}]
  wire  _GEN_162 = 6'h2c == outputBuffer_rs2Addr ? PRFValidList_44 : _GEN_161; // @[decode.scala 250:{60,60}]
  wire  _GEN_163 = 6'h2d == outputBuffer_rs2Addr ? PRFValidList_45 : _GEN_162; // @[decode.scala 250:{60,60}]
  wire  _GEN_164 = 6'h2e == outputBuffer_rs2Addr ? PRFValidList_46 : _GEN_163; // @[decode.scala 250:{60,60}]
  wire  _GEN_165 = 6'h2f == outputBuffer_rs2Addr ? PRFValidList_47 : _GEN_164; // @[decode.scala 250:{60,60}]
  wire  _GEN_166 = 6'h30 == outputBuffer_rs2Addr ? PRFValidList_48 : _GEN_165; // @[decode.scala 250:{60,60}]
  wire  _GEN_167 = 6'h31 == outputBuffer_rs2Addr ? PRFValidList_49 : _GEN_166; // @[decode.scala 250:{60,60}]
  wire  _GEN_168 = 6'h32 == outputBuffer_rs2Addr ? PRFValidList_50 : _GEN_167; // @[decode.scala 250:{60,60}]
  wire  _GEN_169 = 6'h33 == outputBuffer_rs2Addr ? PRFValidList_51 : _GEN_168; // @[decode.scala 250:{60,60}]
  wire  _GEN_170 = 6'h34 == outputBuffer_rs2Addr ? PRFValidList_52 : _GEN_169; // @[decode.scala 250:{60,60}]
  wire  _GEN_171 = 6'h35 == outputBuffer_rs2Addr ? PRFValidList_53 : _GEN_170; // @[decode.scala 250:{60,60}]
  wire  _GEN_172 = 6'h36 == outputBuffer_rs2Addr ? PRFValidList_54 : _GEN_171; // @[decode.scala 250:{60,60}]
  wire  _GEN_173 = 6'h37 == outputBuffer_rs2Addr ? PRFValidList_55 : _GEN_172; // @[decode.scala 250:{60,60}]
  wire  _GEN_174 = 6'h38 == outputBuffer_rs2Addr ? PRFValidList_56 : _GEN_173; // @[decode.scala 250:{60,60}]
  wire  _GEN_175 = 6'h39 == outputBuffer_rs2Addr ? PRFValidList_57 : _GEN_174; // @[decode.scala 250:{60,60}]
  wire  _GEN_176 = 6'h3a == outputBuffer_rs2Addr ? PRFValidList_58 : _GEN_175; // @[decode.scala 250:{60,60}]
  wire  _GEN_177 = 6'h3b == outputBuffer_rs2Addr ? PRFValidList_59 : _GEN_176; // @[decode.scala 250:{60,60}]
  wire  _GEN_178 = 6'h3c == outputBuffer_rs2Addr ? PRFValidList_60 : _GEN_177; // @[decode.scala 250:{60,60}]
  wire  _GEN_179 = 6'h3d == outputBuffer_rs2Addr ? PRFValidList_61 : _GEN_178; // @[decode.scala 250:{60,60}]
  wire  _GEN_180 = 6'h3e == outputBuffer_rs2Addr ? PRFValidList_62 : _GEN_179; // @[decode.scala 250:{60,60}]
  wire  _GEN_181 = 6'h3f == outputBuffer_rs2Addr ? PRFValidList_63 : _GEN_180; // @[decode.scala 250:{60,60}]
  wire [1:0] toExec_branchMask_lo = {branchBuffer_branchMask_1,branchBuffer_branchMask_0}; // @[decode.scala 252:49]
  wire [1:0] toExec_branchMask_hi = {branchBuffer_branchMask_3,branchBuffer_branchMask_2}; // @[decode.scala 252:49]
  wire [3:0] _toExec_branchMask_T = {branchBuffer_branchMask_3,branchBuffer_branchMask_2,branchBuffer_branchMask_1,
    branchBuffer_branchMask_0}; // @[decode.scala 252:49]
  wire  _fromFetch_expected_valid_T = expectedPC != 64'h0; // @[decode.scala 255:42]
  wire  unconditionalJumps = outputBuffer_instruction[6:0] == 7'h6f | outputBuffer_instruction[6:0] == 7'h67 |
    outputBuffer_instruction[6:0] == 7'h37 | outputBuffer_instruction[6:0] == 7'h17; // @[decode.scala 298:154]
  wire  csrIns = outputBuffer_instruction[6:0] == 7'h73 & outputBuffer_instruction[14:12] != 3'h0; // @[decode.scala 299:56]
  wire  validOutputBuf = ~stateRegOutputBuf ? 1'h0 : stateRegOutputBuf & _GEN_9096; // @[decode.scala 813:29]
  wire [31:0] _jumpAddrWrite_linkAddr_T_2 = outputBuffer_instruction[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _jumpAddrWrite_linkAddr_T_4 = {_jumpAddrWrite_linkAddr_T_2,outputBuffer_instruction[31:12],12'h0}; // @[Cat.scala 33:92]
  wire [63:0] _jumpAddrWrite_linkAddr_T_6 = outputBuffer_pc + _jumpAddrWrite_linkAddr_T_4; // @[decode.scala 262:24]
  wire [63:0] _jumpAddrWrite_linkAddr_T_13 = outputBuffer_pc + 64'h4; // @[decode.scala 265:23]
  wire [63:0] _GEN_183 = 2'h1 == outputBuffer_instruction[6:5] ? _jumpAddrWrite_linkAddr_T_4 :
    _jumpAddrWrite_linkAddr_T_6; // @[decode.scala 261:{28,28}]
  wire [63:0] _GEN_184 = 2'h2 == outputBuffer_instruction[6:5] ? 64'h0 : _GEN_183; // @[decode.scala 261:{28,28}]
  wire [63:0] _GEN_185 = 2'h3 == outputBuffer_instruction[6:5] ? _jumpAddrWrite_linkAddr_T_13 : _GEN_184; // @[decode.scala 261:{28,28}]
  wire [2:0] fun3 = inputBuffer_instruction[14:12]; // @[decode.scala 293:16]
  reg [5:0] architecturalRegMap_0; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_1; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_2; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_3; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_4; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_5; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_6; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_7; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_8; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_9; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_10; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_11; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_12; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_13; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_14; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_15; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_16; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_17; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_18; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_19; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_20; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_21; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_22; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_23; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_24; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_25; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_26; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_27; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_28; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_29; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_30; // @[decode.scala 302:36]
  reg [5:0] architecturalRegMap_31; // @[decode.scala 302:36]
  reg [5:0] reservedRegMap1_0; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_1; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_2; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_3; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_4; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_5; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_6; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_7; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_8; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_9; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_10; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_11; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_12; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_13; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_14; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_15; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_16; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_17; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_18; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_19; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_20; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_21; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_22; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_23; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_24; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_25; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_26; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_27; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_28; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_29; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_30; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap1_31; // @[decode.scala 310:28]
  reg [5:0] reservedRegMap2_0; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_1; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_2; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_3; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_4; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_5; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_6; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_7; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_8; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_9; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_10; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_11; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_12; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_13; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_14; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_15; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_16; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_17; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_18; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_19; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_20; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_21; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_22; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_23; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_24; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_25; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_26; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_27; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_28; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_29; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_30; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap2_31; // @[decode.scala 311:28]
  reg [5:0] reservedRegMap3_0; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_1; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_2; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_3; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_4; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_5; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_6; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_7; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_8; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_9; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_10; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_11; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_12; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_13; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_14; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_15; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_16; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_17; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_18; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_19; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_20; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_21; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_22; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_23; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_24; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_25; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_26; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_27; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_28; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_29; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_30; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap3_31; // @[decode.scala 312:28]
  reg [5:0] reservedRegMap4_0; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_1; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_2; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_3; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_4; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_5; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_6; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_7; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_8; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_9; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_10; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_11; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_12; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_13; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_14; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_15; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_16; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_17; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_18; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_19; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_20; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_21; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_22; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_23; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_24; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_25; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_26; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_27; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_28; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_29; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_30; // @[decode.scala 313:28]
  reg [5:0] reservedRegMap4_31; // @[decode.scala 313:28]
  reg  reservedFreeList1_0; // @[decode.scala 315:30]
  reg  reservedFreeList1_1; // @[decode.scala 315:30]
  reg  reservedFreeList1_2; // @[decode.scala 315:30]
  reg  reservedFreeList1_3; // @[decode.scala 315:30]
  reg  reservedFreeList1_4; // @[decode.scala 315:30]
  reg  reservedFreeList1_5; // @[decode.scala 315:30]
  reg  reservedFreeList1_6; // @[decode.scala 315:30]
  reg  reservedFreeList1_7; // @[decode.scala 315:30]
  reg  reservedFreeList1_8; // @[decode.scala 315:30]
  reg  reservedFreeList1_9; // @[decode.scala 315:30]
  reg  reservedFreeList1_10; // @[decode.scala 315:30]
  reg  reservedFreeList1_11; // @[decode.scala 315:30]
  reg  reservedFreeList1_12; // @[decode.scala 315:30]
  reg  reservedFreeList1_13; // @[decode.scala 315:30]
  reg  reservedFreeList1_14; // @[decode.scala 315:30]
  reg  reservedFreeList1_15; // @[decode.scala 315:30]
  reg  reservedFreeList1_16; // @[decode.scala 315:30]
  reg  reservedFreeList1_17; // @[decode.scala 315:30]
  reg  reservedFreeList1_18; // @[decode.scala 315:30]
  reg  reservedFreeList1_19; // @[decode.scala 315:30]
  reg  reservedFreeList1_20; // @[decode.scala 315:30]
  reg  reservedFreeList1_21; // @[decode.scala 315:30]
  reg  reservedFreeList1_22; // @[decode.scala 315:30]
  reg  reservedFreeList1_23; // @[decode.scala 315:30]
  reg  reservedFreeList1_24; // @[decode.scala 315:30]
  reg  reservedFreeList1_25; // @[decode.scala 315:30]
  reg  reservedFreeList1_26; // @[decode.scala 315:30]
  reg  reservedFreeList1_27; // @[decode.scala 315:30]
  reg  reservedFreeList1_28; // @[decode.scala 315:30]
  reg  reservedFreeList1_29; // @[decode.scala 315:30]
  reg  reservedFreeList1_30; // @[decode.scala 315:30]
  reg  reservedFreeList1_31; // @[decode.scala 315:30]
  reg  reservedFreeList1_32; // @[decode.scala 315:30]
  reg  reservedFreeList1_33; // @[decode.scala 315:30]
  reg  reservedFreeList1_34; // @[decode.scala 315:30]
  reg  reservedFreeList1_35; // @[decode.scala 315:30]
  reg  reservedFreeList1_36; // @[decode.scala 315:30]
  reg  reservedFreeList1_37; // @[decode.scala 315:30]
  reg  reservedFreeList1_38; // @[decode.scala 315:30]
  reg  reservedFreeList1_39; // @[decode.scala 315:30]
  reg  reservedFreeList1_40; // @[decode.scala 315:30]
  reg  reservedFreeList1_41; // @[decode.scala 315:30]
  reg  reservedFreeList1_42; // @[decode.scala 315:30]
  reg  reservedFreeList1_43; // @[decode.scala 315:30]
  reg  reservedFreeList1_44; // @[decode.scala 315:30]
  reg  reservedFreeList1_45; // @[decode.scala 315:30]
  reg  reservedFreeList1_46; // @[decode.scala 315:30]
  reg  reservedFreeList1_47; // @[decode.scala 315:30]
  reg  reservedFreeList1_48; // @[decode.scala 315:30]
  reg  reservedFreeList1_49; // @[decode.scala 315:30]
  reg  reservedFreeList1_50; // @[decode.scala 315:30]
  reg  reservedFreeList1_51; // @[decode.scala 315:30]
  reg  reservedFreeList1_52; // @[decode.scala 315:30]
  reg  reservedFreeList1_53; // @[decode.scala 315:30]
  reg  reservedFreeList1_54; // @[decode.scala 315:30]
  reg  reservedFreeList1_55; // @[decode.scala 315:30]
  reg  reservedFreeList1_56; // @[decode.scala 315:30]
  reg  reservedFreeList1_57; // @[decode.scala 315:30]
  reg  reservedFreeList1_58; // @[decode.scala 315:30]
  reg  reservedFreeList1_59; // @[decode.scala 315:30]
  reg  reservedFreeList1_60; // @[decode.scala 315:30]
  reg  reservedFreeList1_61; // @[decode.scala 315:30]
  reg  reservedFreeList1_62; // @[decode.scala 315:30]
  reg  reservedFreeList2_0; // @[decode.scala 316:30]
  reg  reservedFreeList2_1; // @[decode.scala 316:30]
  reg  reservedFreeList2_2; // @[decode.scala 316:30]
  reg  reservedFreeList2_3; // @[decode.scala 316:30]
  reg  reservedFreeList2_4; // @[decode.scala 316:30]
  reg  reservedFreeList2_5; // @[decode.scala 316:30]
  reg  reservedFreeList2_6; // @[decode.scala 316:30]
  reg  reservedFreeList2_7; // @[decode.scala 316:30]
  reg  reservedFreeList2_8; // @[decode.scala 316:30]
  reg  reservedFreeList2_9; // @[decode.scala 316:30]
  reg  reservedFreeList2_10; // @[decode.scala 316:30]
  reg  reservedFreeList2_11; // @[decode.scala 316:30]
  reg  reservedFreeList2_12; // @[decode.scala 316:30]
  reg  reservedFreeList2_13; // @[decode.scala 316:30]
  reg  reservedFreeList2_14; // @[decode.scala 316:30]
  reg  reservedFreeList2_15; // @[decode.scala 316:30]
  reg  reservedFreeList2_16; // @[decode.scala 316:30]
  reg  reservedFreeList2_17; // @[decode.scala 316:30]
  reg  reservedFreeList2_18; // @[decode.scala 316:30]
  reg  reservedFreeList2_19; // @[decode.scala 316:30]
  reg  reservedFreeList2_20; // @[decode.scala 316:30]
  reg  reservedFreeList2_21; // @[decode.scala 316:30]
  reg  reservedFreeList2_22; // @[decode.scala 316:30]
  reg  reservedFreeList2_23; // @[decode.scala 316:30]
  reg  reservedFreeList2_24; // @[decode.scala 316:30]
  reg  reservedFreeList2_25; // @[decode.scala 316:30]
  reg  reservedFreeList2_26; // @[decode.scala 316:30]
  reg  reservedFreeList2_27; // @[decode.scala 316:30]
  reg  reservedFreeList2_28; // @[decode.scala 316:30]
  reg  reservedFreeList2_29; // @[decode.scala 316:30]
  reg  reservedFreeList2_30; // @[decode.scala 316:30]
  reg  reservedFreeList2_31; // @[decode.scala 316:30]
  reg  reservedFreeList2_32; // @[decode.scala 316:30]
  reg  reservedFreeList2_33; // @[decode.scala 316:30]
  reg  reservedFreeList2_34; // @[decode.scala 316:30]
  reg  reservedFreeList2_35; // @[decode.scala 316:30]
  reg  reservedFreeList2_36; // @[decode.scala 316:30]
  reg  reservedFreeList2_37; // @[decode.scala 316:30]
  reg  reservedFreeList2_38; // @[decode.scala 316:30]
  reg  reservedFreeList2_39; // @[decode.scala 316:30]
  reg  reservedFreeList2_40; // @[decode.scala 316:30]
  reg  reservedFreeList2_41; // @[decode.scala 316:30]
  reg  reservedFreeList2_42; // @[decode.scala 316:30]
  reg  reservedFreeList2_43; // @[decode.scala 316:30]
  reg  reservedFreeList2_44; // @[decode.scala 316:30]
  reg  reservedFreeList2_45; // @[decode.scala 316:30]
  reg  reservedFreeList2_46; // @[decode.scala 316:30]
  reg  reservedFreeList2_47; // @[decode.scala 316:30]
  reg  reservedFreeList2_48; // @[decode.scala 316:30]
  reg  reservedFreeList2_49; // @[decode.scala 316:30]
  reg  reservedFreeList2_50; // @[decode.scala 316:30]
  reg  reservedFreeList2_51; // @[decode.scala 316:30]
  reg  reservedFreeList2_52; // @[decode.scala 316:30]
  reg  reservedFreeList2_53; // @[decode.scala 316:30]
  reg  reservedFreeList2_54; // @[decode.scala 316:30]
  reg  reservedFreeList2_55; // @[decode.scala 316:30]
  reg  reservedFreeList2_56; // @[decode.scala 316:30]
  reg  reservedFreeList2_57; // @[decode.scala 316:30]
  reg  reservedFreeList2_58; // @[decode.scala 316:30]
  reg  reservedFreeList2_59; // @[decode.scala 316:30]
  reg  reservedFreeList2_60; // @[decode.scala 316:30]
  reg  reservedFreeList2_61; // @[decode.scala 316:30]
  reg  reservedFreeList2_62; // @[decode.scala 316:30]
  reg  reservedFreeList3_0; // @[decode.scala 317:30]
  reg  reservedFreeList3_1; // @[decode.scala 317:30]
  reg  reservedFreeList3_2; // @[decode.scala 317:30]
  reg  reservedFreeList3_3; // @[decode.scala 317:30]
  reg  reservedFreeList3_4; // @[decode.scala 317:30]
  reg  reservedFreeList3_5; // @[decode.scala 317:30]
  reg  reservedFreeList3_6; // @[decode.scala 317:30]
  reg  reservedFreeList3_7; // @[decode.scala 317:30]
  reg  reservedFreeList3_8; // @[decode.scala 317:30]
  reg  reservedFreeList3_9; // @[decode.scala 317:30]
  reg  reservedFreeList3_10; // @[decode.scala 317:30]
  reg  reservedFreeList3_11; // @[decode.scala 317:30]
  reg  reservedFreeList3_12; // @[decode.scala 317:30]
  reg  reservedFreeList3_13; // @[decode.scala 317:30]
  reg  reservedFreeList3_14; // @[decode.scala 317:30]
  reg  reservedFreeList3_15; // @[decode.scala 317:30]
  reg  reservedFreeList3_16; // @[decode.scala 317:30]
  reg  reservedFreeList3_17; // @[decode.scala 317:30]
  reg  reservedFreeList3_18; // @[decode.scala 317:30]
  reg  reservedFreeList3_19; // @[decode.scala 317:30]
  reg  reservedFreeList3_20; // @[decode.scala 317:30]
  reg  reservedFreeList3_21; // @[decode.scala 317:30]
  reg  reservedFreeList3_22; // @[decode.scala 317:30]
  reg  reservedFreeList3_23; // @[decode.scala 317:30]
  reg  reservedFreeList3_24; // @[decode.scala 317:30]
  reg  reservedFreeList3_25; // @[decode.scala 317:30]
  reg  reservedFreeList3_26; // @[decode.scala 317:30]
  reg  reservedFreeList3_27; // @[decode.scala 317:30]
  reg  reservedFreeList3_28; // @[decode.scala 317:30]
  reg  reservedFreeList3_29; // @[decode.scala 317:30]
  reg  reservedFreeList3_30; // @[decode.scala 317:30]
  reg  reservedFreeList3_31; // @[decode.scala 317:30]
  reg  reservedFreeList3_32; // @[decode.scala 317:30]
  reg  reservedFreeList3_33; // @[decode.scala 317:30]
  reg  reservedFreeList3_34; // @[decode.scala 317:30]
  reg  reservedFreeList3_35; // @[decode.scala 317:30]
  reg  reservedFreeList3_36; // @[decode.scala 317:30]
  reg  reservedFreeList3_37; // @[decode.scala 317:30]
  reg  reservedFreeList3_38; // @[decode.scala 317:30]
  reg  reservedFreeList3_39; // @[decode.scala 317:30]
  reg  reservedFreeList3_40; // @[decode.scala 317:30]
  reg  reservedFreeList3_41; // @[decode.scala 317:30]
  reg  reservedFreeList3_42; // @[decode.scala 317:30]
  reg  reservedFreeList3_43; // @[decode.scala 317:30]
  reg  reservedFreeList3_44; // @[decode.scala 317:30]
  reg  reservedFreeList3_45; // @[decode.scala 317:30]
  reg  reservedFreeList3_46; // @[decode.scala 317:30]
  reg  reservedFreeList3_47; // @[decode.scala 317:30]
  reg  reservedFreeList3_48; // @[decode.scala 317:30]
  reg  reservedFreeList3_49; // @[decode.scala 317:30]
  reg  reservedFreeList3_50; // @[decode.scala 317:30]
  reg  reservedFreeList3_51; // @[decode.scala 317:30]
  reg  reservedFreeList3_52; // @[decode.scala 317:30]
  reg  reservedFreeList3_53; // @[decode.scala 317:30]
  reg  reservedFreeList3_54; // @[decode.scala 317:30]
  reg  reservedFreeList3_55; // @[decode.scala 317:30]
  reg  reservedFreeList3_56; // @[decode.scala 317:30]
  reg  reservedFreeList3_57; // @[decode.scala 317:30]
  reg  reservedFreeList3_58; // @[decode.scala 317:30]
  reg  reservedFreeList3_59; // @[decode.scala 317:30]
  reg  reservedFreeList3_60; // @[decode.scala 317:30]
  reg  reservedFreeList3_61; // @[decode.scala 317:30]
  reg  reservedFreeList3_62; // @[decode.scala 317:30]
  reg  reservedFreeList4_0; // @[decode.scala 318:30]
  reg  reservedFreeList4_1; // @[decode.scala 318:30]
  reg  reservedFreeList4_2; // @[decode.scala 318:30]
  reg  reservedFreeList4_3; // @[decode.scala 318:30]
  reg  reservedFreeList4_4; // @[decode.scala 318:30]
  reg  reservedFreeList4_5; // @[decode.scala 318:30]
  reg  reservedFreeList4_6; // @[decode.scala 318:30]
  reg  reservedFreeList4_7; // @[decode.scala 318:30]
  reg  reservedFreeList4_8; // @[decode.scala 318:30]
  reg  reservedFreeList4_9; // @[decode.scala 318:30]
  reg  reservedFreeList4_10; // @[decode.scala 318:30]
  reg  reservedFreeList4_11; // @[decode.scala 318:30]
  reg  reservedFreeList4_12; // @[decode.scala 318:30]
  reg  reservedFreeList4_13; // @[decode.scala 318:30]
  reg  reservedFreeList4_14; // @[decode.scala 318:30]
  reg  reservedFreeList4_15; // @[decode.scala 318:30]
  reg  reservedFreeList4_16; // @[decode.scala 318:30]
  reg  reservedFreeList4_17; // @[decode.scala 318:30]
  reg  reservedFreeList4_18; // @[decode.scala 318:30]
  reg  reservedFreeList4_19; // @[decode.scala 318:30]
  reg  reservedFreeList4_20; // @[decode.scala 318:30]
  reg  reservedFreeList4_21; // @[decode.scala 318:30]
  reg  reservedFreeList4_22; // @[decode.scala 318:30]
  reg  reservedFreeList4_23; // @[decode.scala 318:30]
  reg  reservedFreeList4_24; // @[decode.scala 318:30]
  reg  reservedFreeList4_25; // @[decode.scala 318:30]
  reg  reservedFreeList4_26; // @[decode.scala 318:30]
  reg  reservedFreeList4_27; // @[decode.scala 318:30]
  reg  reservedFreeList4_28; // @[decode.scala 318:30]
  reg  reservedFreeList4_29; // @[decode.scala 318:30]
  reg  reservedFreeList4_30; // @[decode.scala 318:30]
  reg  reservedFreeList4_31; // @[decode.scala 318:30]
  reg  reservedFreeList4_32; // @[decode.scala 318:30]
  reg  reservedFreeList4_33; // @[decode.scala 318:30]
  reg  reservedFreeList4_34; // @[decode.scala 318:30]
  reg  reservedFreeList4_35; // @[decode.scala 318:30]
  reg  reservedFreeList4_36; // @[decode.scala 318:30]
  reg  reservedFreeList4_37; // @[decode.scala 318:30]
  reg  reservedFreeList4_38; // @[decode.scala 318:30]
  reg  reservedFreeList4_39; // @[decode.scala 318:30]
  reg  reservedFreeList4_40; // @[decode.scala 318:30]
  reg  reservedFreeList4_41; // @[decode.scala 318:30]
  reg  reservedFreeList4_42; // @[decode.scala 318:30]
  reg  reservedFreeList4_43; // @[decode.scala 318:30]
  reg  reservedFreeList4_44; // @[decode.scala 318:30]
  reg  reservedFreeList4_45; // @[decode.scala 318:30]
  reg  reservedFreeList4_46; // @[decode.scala 318:30]
  reg  reservedFreeList4_47; // @[decode.scala 318:30]
  reg  reservedFreeList4_48; // @[decode.scala 318:30]
  reg  reservedFreeList4_49; // @[decode.scala 318:30]
  reg  reservedFreeList4_50; // @[decode.scala 318:30]
  reg  reservedFreeList4_51; // @[decode.scala 318:30]
  reg  reservedFreeList4_52; // @[decode.scala 318:30]
  reg  reservedFreeList4_53; // @[decode.scala 318:30]
  reg  reservedFreeList4_54; // @[decode.scala 318:30]
  reg  reservedFreeList4_55; // @[decode.scala 318:30]
  reg  reservedFreeList4_56; // @[decode.scala 318:30]
  reg  reservedFreeList4_57; // @[decode.scala 318:30]
  reg  reservedFreeList4_58; // @[decode.scala 318:30]
  reg  reservedFreeList4_59; // @[decode.scala 318:30]
  reg  reservedFreeList4_60; // @[decode.scala 318:30]
  reg  reservedFreeList4_61; // @[decode.scala 318:30]
  reg  reservedFreeList4_62; // @[decode.scala 318:30]
  reg  reservedValidList1_0; // @[decode.scala 320:31]
  reg  reservedValidList1_1; // @[decode.scala 320:31]
  reg  reservedValidList1_2; // @[decode.scala 320:31]
  reg  reservedValidList1_3; // @[decode.scala 320:31]
  reg  reservedValidList1_4; // @[decode.scala 320:31]
  reg  reservedValidList1_5; // @[decode.scala 320:31]
  reg  reservedValidList1_6; // @[decode.scala 320:31]
  reg  reservedValidList1_7; // @[decode.scala 320:31]
  reg  reservedValidList1_8; // @[decode.scala 320:31]
  reg  reservedValidList1_9; // @[decode.scala 320:31]
  reg  reservedValidList1_10; // @[decode.scala 320:31]
  reg  reservedValidList1_11; // @[decode.scala 320:31]
  reg  reservedValidList1_12; // @[decode.scala 320:31]
  reg  reservedValidList1_13; // @[decode.scala 320:31]
  reg  reservedValidList1_14; // @[decode.scala 320:31]
  reg  reservedValidList1_15; // @[decode.scala 320:31]
  reg  reservedValidList1_16; // @[decode.scala 320:31]
  reg  reservedValidList1_17; // @[decode.scala 320:31]
  reg  reservedValidList1_18; // @[decode.scala 320:31]
  reg  reservedValidList1_19; // @[decode.scala 320:31]
  reg  reservedValidList1_20; // @[decode.scala 320:31]
  reg  reservedValidList1_21; // @[decode.scala 320:31]
  reg  reservedValidList1_22; // @[decode.scala 320:31]
  reg  reservedValidList1_23; // @[decode.scala 320:31]
  reg  reservedValidList1_24; // @[decode.scala 320:31]
  reg  reservedValidList1_25; // @[decode.scala 320:31]
  reg  reservedValidList1_26; // @[decode.scala 320:31]
  reg  reservedValidList1_27; // @[decode.scala 320:31]
  reg  reservedValidList1_28; // @[decode.scala 320:31]
  reg  reservedValidList1_29; // @[decode.scala 320:31]
  reg  reservedValidList1_30; // @[decode.scala 320:31]
  reg  reservedValidList1_31; // @[decode.scala 320:31]
  reg  reservedValidList1_32; // @[decode.scala 320:31]
  reg  reservedValidList1_33; // @[decode.scala 320:31]
  reg  reservedValidList1_34; // @[decode.scala 320:31]
  reg  reservedValidList1_35; // @[decode.scala 320:31]
  reg  reservedValidList1_36; // @[decode.scala 320:31]
  reg  reservedValidList1_37; // @[decode.scala 320:31]
  reg  reservedValidList1_38; // @[decode.scala 320:31]
  reg  reservedValidList1_39; // @[decode.scala 320:31]
  reg  reservedValidList1_40; // @[decode.scala 320:31]
  reg  reservedValidList1_41; // @[decode.scala 320:31]
  reg  reservedValidList1_42; // @[decode.scala 320:31]
  reg  reservedValidList1_43; // @[decode.scala 320:31]
  reg  reservedValidList1_44; // @[decode.scala 320:31]
  reg  reservedValidList1_45; // @[decode.scala 320:31]
  reg  reservedValidList1_46; // @[decode.scala 320:31]
  reg  reservedValidList1_47; // @[decode.scala 320:31]
  reg  reservedValidList1_48; // @[decode.scala 320:31]
  reg  reservedValidList1_49; // @[decode.scala 320:31]
  reg  reservedValidList1_50; // @[decode.scala 320:31]
  reg  reservedValidList1_51; // @[decode.scala 320:31]
  reg  reservedValidList1_52; // @[decode.scala 320:31]
  reg  reservedValidList1_53; // @[decode.scala 320:31]
  reg  reservedValidList1_54; // @[decode.scala 320:31]
  reg  reservedValidList1_55; // @[decode.scala 320:31]
  reg  reservedValidList1_56; // @[decode.scala 320:31]
  reg  reservedValidList1_57; // @[decode.scala 320:31]
  reg  reservedValidList1_58; // @[decode.scala 320:31]
  reg  reservedValidList1_59; // @[decode.scala 320:31]
  reg  reservedValidList1_60; // @[decode.scala 320:31]
  reg  reservedValidList1_61; // @[decode.scala 320:31]
  reg  reservedValidList1_62; // @[decode.scala 320:31]
  reg  reservedValidList1_63; // @[decode.scala 320:31]
  reg  reservedValidList2_0; // @[decode.scala 321:31]
  reg  reservedValidList2_1; // @[decode.scala 321:31]
  reg  reservedValidList2_2; // @[decode.scala 321:31]
  reg  reservedValidList2_3; // @[decode.scala 321:31]
  reg  reservedValidList2_4; // @[decode.scala 321:31]
  reg  reservedValidList2_5; // @[decode.scala 321:31]
  reg  reservedValidList2_6; // @[decode.scala 321:31]
  reg  reservedValidList2_7; // @[decode.scala 321:31]
  reg  reservedValidList2_8; // @[decode.scala 321:31]
  reg  reservedValidList2_9; // @[decode.scala 321:31]
  reg  reservedValidList2_10; // @[decode.scala 321:31]
  reg  reservedValidList2_11; // @[decode.scala 321:31]
  reg  reservedValidList2_12; // @[decode.scala 321:31]
  reg  reservedValidList2_13; // @[decode.scala 321:31]
  reg  reservedValidList2_14; // @[decode.scala 321:31]
  reg  reservedValidList2_15; // @[decode.scala 321:31]
  reg  reservedValidList2_16; // @[decode.scala 321:31]
  reg  reservedValidList2_17; // @[decode.scala 321:31]
  reg  reservedValidList2_18; // @[decode.scala 321:31]
  reg  reservedValidList2_19; // @[decode.scala 321:31]
  reg  reservedValidList2_20; // @[decode.scala 321:31]
  reg  reservedValidList2_21; // @[decode.scala 321:31]
  reg  reservedValidList2_22; // @[decode.scala 321:31]
  reg  reservedValidList2_23; // @[decode.scala 321:31]
  reg  reservedValidList2_24; // @[decode.scala 321:31]
  reg  reservedValidList2_25; // @[decode.scala 321:31]
  reg  reservedValidList2_26; // @[decode.scala 321:31]
  reg  reservedValidList2_27; // @[decode.scala 321:31]
  reg  reservedValidList2_28; // @[decode.scala 321:31]
  reg  reservedValidList2_29; // @[decode.scala 321:31]
  reg  reservedValidList2_30; // @[decode.scala 321:31]
  reg  reservedValidList2_31; // @[decode.scala 321:31]
  reg  reservedValidList2_32; // @[decode.scala 321:31]
  reg  reservedValidList2_33; // @[decode.scala 321:31]
  reg  reservedValidList2_34; // @[decode.scala 321:31]
  reg  reservedValidList2_35; // @[decode.scala 321:31]
  reg  reservedValidList2_36; // @[decode.scala 321:31]
  reg  reservedValidList2_37; // @[decode.scala 321:31]
  reg  reservedValidList2_38; // @[decode.scala 321:31]
  reg  reservedValidList2_39; // @[decode.scala 321:31]
  reg  reservedValidList2_40; // @[decode.scala 321:31]
  reg  reservedValidList2_41; // @[decode.scala 321:31]
  reg  reservedValidList2_42; // @[decode.scala 321:31]
  reg  reservedValidList2_43; // @[decode.scala 321:31]
  reg  reservedValidList2_44; // @[decode.scala 321:31]
  reg  reservedValidList2_45; // @[decode.scala 321:31]
  reg  reservedValidList2_46; // @[decode.scala 321:31]
  reg  reservedValidList2_47; // @[decode.scala 321:31]
  reg  reservedValidList2_48; // @[decode.scala 321:31]
  reg  reservedValidList2_49; // @[decode.scala 321:31]
  reg  reservedValidList2_50; // @[decode.scala 321:31]
  reg  reservedValidList2_51; // @[decode.scala 321:31]
  reg  reservedValidList2_52; // @[decode.scala 321:31]
  reg  reservedValidList2_53; // @[decode.scala 321:31]
  reg  reservedValidList2_54; // @[decode.scala 321:31]
  reg  reservedValidList2_55; // @[decode.scala 321:31]
  reg  reservedValidList2_56; // @[decode.scala 321:31]
  reg  reservedValidList2_57; // @[decode.scala 321:31]
  reg  reservedValidList2_58; // @[decode.scala 321:31]
  reg  reservedValidList2_59; // @[decode.scala 321:31]
  reg  reservedValidList2_60; // @[decode.scala 321:31]
  reg  reservedValidList2_61; // @[decode.scala 321:31]
  reg  reservedValidList2_62; // @[decode.scala 321:31]
  reg  reservedValidList2_63; // @[decode.scala 321:31]
  reg  reservedValidList3_0; // @[decode.scala 322:31]
  reg  reservedValidList3_1; // @[decode.scala 322:31]
  reg  reservedValidList3_2; // @[decode.scala 322:31]
  reg  reservedValidList3_3; // @[decode.scala 322:31]
  reg  reservedValidList3_4; // @[decode.scala 322:31]
  reg  reservedValidList3_5; // @[decode.scala 322:31]
  reg  reservedValidList3_6; // @[decode.scala 322:31]
  reg  reservedValidList3_7; // @[decode.scala 322:31]
  reg  reservedValidList3_8; // @[decode.scala 322:31]
  reg  reservedValidList3_9; // @[decode.scala 322:31]
  reg  reservedValidList3_10; // @[decode.scala 322:31]
  reg  reservedValidList3_11; // @[decode.scala 322:31]
  reg  reservedValidList3_12; // @[decode.scala 322:31]
  reg  reservedValidList3_13; // @[decode.scala 322:31]
  reg  reservedValidList3_14; // @[decode.scala 322:31]
  reg  reservedValidList3_15; // @[decode.scala 322:31]
  reg  reservedValidList3_16; // @[decode.scala 322:31]
  reg  reservedValidList3_17; // @[decode.scala 322:31]
  reg  reservedValidList3_18; // @[decode.scala 322:31]
  reg  reservedValidList3_19; // @[decode.scala 322:31]
  reg  reservedValidList3_20; // @[decode.scala 322:31]
  reg  reservedValidList3_21; // @[decode.scala 322:31]
  reg  reservedValidList3_22; // @[decode.scala 322:31]
  reg  reservedValidList3_23; // @[decode.scala 322:31]
  reg  reservedValidList3_24; // @[decode.scala 322:31]
  reg  reservedValidList3_25; // @[decode.scala 322:31]
  reg  reservedValidList3_26; // @[decode.scala 322:31]
  reg  reservedValidList3_27; // @[decode.scala 322:31]
  reg  reservedValidList3_28; // @[decode.scala 322:31]
  reg  reservedValidList3_29; // @[decode.scala 322:31]
  reg  reservedValidList3_30; // @[decode.scala 322:31]
  reg  reservedValidList3_31; // @[decode.scala 322:31]
  reg  reservedValidList3_32; // @[decode.scala 322:31]
  reg  reservedValidList3_33; // @[decode.scala 322:31]
  reg  reservedValidList3_34; // @[decode.scala 322:31]
  reg  reservedValidList3_35; // @[decode.scala 322:31]
  reg  reservedValidList3_36; // @[decode.scala 322:31]
  reg  reservedValidList3_37; // @[decode.scala 322:31]
  reg  reservedValidList3_38; // @[decode.scala 322:31]
  reg  reservedValidList3_39; // @[decode.scala 322:31]
  reg  reservedValidList3_40; // @[decode.scala 322:31]
  reg  reservedValidList3_41; // @[decode.scala 322:31]
  reg  reservedValidList3_42; // @[decode.scala 322:31]
  reg  reservedValidList3_43; // @[decode.scala 322:31]
  reg  reservedValidList3_44; // @[decode.scala 322:31]
  reg  reservedValidList3_45; // @[decode.scala 322:31]
  reg  reservedValidList3_46; // @[decode.scala 322:31]
  reg  reservedValidList3_47; // @[decode.scala 322:31]
  reg  reservedValidList3_48; // @[decode.scala 322:31]
  reg  reservedValidList3_49; // @[decode.scala 322:31]
  reg  reservedValidList3_50; // @[decode.scala 322:31]
  reg  reservedValidList3_51; // @[decode.scala 322:31]
  reg  reservedValidList3_52; // @[decode.scala 322:31]
  reg  reservedValidList3_53; // @[decode.scala 322:31]
  reg  reservedValidList3_54; // @[decode.scala 322:31]
  reg  reservedValidList3_55; // @[decode.scala 322:31]
  reg  reservedValidList3_56; // @[decode.scala 322:31]
  reg  reservedValidList3_57; // @[decode.scala 322:31]
  reg  reservedValidList3_58; // @[decode.scala 322:31]
  reg  reservedValidList3_59; // @[decode.scala 322:31]
  reg  reservedValidList3_60; // @[decode.scala 322:31]
  reg  reservedValidList3_61; // @[decode.scala 322:31]
  reg  reservedValidList3_62; // @[decode.scala 322:31]
  reg  reservedValidList3_63; // @[decode.scala 322:31]
  reg  reservedValidList4_0; // @[decode.scala 323:31]
  reg  reservedValidList4_1; // @[decode.scala 323:31]
  reg  reservedValidList4_2; // @[decode.scala 323:31]
  reg  reservedValidList4_3; // @[decode.scala 323:31]
  reg  reservedValidList4_4; // @[decode.scala 323:31]
  reg  reservedValidList4_5; // @[decode.scala 323:31]
  reg  reservedValidList4_6; // @[decode.scala 323:31]
  reg  reservedValidList4_7; // @[decode.scala 323:31]
  reg  reservedValidList4_8; // @[decode.scala 323:31]
  reg  reservedValidList4_9; // @[decode.scala 323:31]
  reg  reservedValidList4_10; // @[decode.scala 323:31]
  reg  reservedValidList4_11; // @[decode.scala 323:31]
  reg  reservedValidList4_12; // @[decode.scala 323:31]
  reg  reservedValidList4_13; // @[decode.scala 323:31]
  reg  reservedValidList4_14; // @[decode.scala 323:31]
  reg  reservedValidList4_15; // @[decode.scala 323:31]
  reg  reservedValidList4_16; // @[decode.scala 323:31]
  reg  reservedValidList4_17; // @[decode.scala 323:31]
  reg  reservedValidList4_18; // @[decode.scala 323:31]
  reg  reservedValidList4_19; // @[decode.scala 323:31]
  reg  reservedValidList4_20; // @[decode.scala 323:31]
  reg  reservedValidList4_21; // @[decode.scala 323:31]
  reg  reservedValidList4_22; // @[decode.scala 323:31]
  reg  reservedValidList4_23; // @[decode.scala 323:31]
  reg  reservedValidList4_24; // @[decode.scala 323:31]
  reg  reservedValidList4_25; // @[decode.scala 323:31]
  reg  reservedValidList4_26; // @[decode.scala 323:31]
  reg  reservedValidList4_27; // @[decode.scala 323:31]
  reg  reservedValidList4_28; // @[decode.scala 323:31]
  reg  reservedValidList4_29; // @[decode.scala 323:31]
  reg  reservedValidList4_30; // @[decode.scala 323:31]
  reg  reservedValidList4_31; // @[decode.scala 323:31]
  reg  reservedValidList4_32; // @[decode.scala 323:31]
  reg  reservedValidList4_33; // @[decode.scala 323:31]
  reg  reservedValidList4_34; // @[decode.scala 323:31]
  reg  reservedValidList4_35; // @[decode.scala 323:31]
  reg  reservedValidList4_36; // @[decode.scala 323:31]
  reg  reservedValidList4_37; // @[decode.scala 323:31]
  reg  reservedValidList4_38; // @[decode.scala 323:31]
  reg  reservedValidList4_39; // @[decode.scala 323:31]
  reg  reservedValidList4_40; // @[decode.scala 323:31]
  reg  reservedValidList4_41; // @[decode.scala 323:31]
  reg  reservedValidList4_42; // @[decode.scala 323:31]
  reg  reservedValidList4_43; // @[decode.scala 323:31]
  reg  reservedValidList4_44; // @[decode.scala 323:31]
  reg  reservedValidList4_45; // @[decode.scala 323:31]
  reg  reservedValidList4_46; // @[decode.scala 323:31]
  reg  reservedValidList4_47; // @[decode.scala 323:31]
  reg  reservedValidList4_48; // @[decode.scala 323:31]
  reg  reservedValidList4_49; // @[decode.scala 323:31]
  reg  reservedValidList4_50; // @[decode.scala 323:31]
  reg  reservedValidList4_51; // @[decode.scala 323:31]
  reg  reservedValidList4_52; // @[decode.scala 323:31]
  reg  reservedValidList4_53; // @[decode.scala 323:31]
  reg  reservedValidList4_54; // @[decode.scala 323:31]
  reg  reservedValidList4_55; // @[decode.scala 323:31]
  reg  reservedValidList4_56; // @[decode.scala 323:31]
  reg  reservedValidList4_57; // @[decode.scala 323:31]
  reg  reservedValidList4_58; // @[decode.scala 323:31]
  reg  reservedValidList4_59; // @[decode.scala 323:31]
  reg  reservedValidList4_60; // @[decode.scala 323:31]
  reg  reservedValidList4_61; // @[decode.scala 323:31]
  reg  reservedValidList4_62; // @[decode.scala 323:31]
  reg  reservedValidList4_63; // @[decode.scala 323:31]
  wire  _GEN_273 = 6'h0 == rs1Addr ? 1'h0 : PRFFreeList_0; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_274 = 6'h1 == rs1Addr ? 1'h0 : PRFFreeList_1; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_275 = 6'h2 == rs1Addr ? 1'h0 : PRFFreeList_2; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_276 = 6'h3 == rs1Addr ? 1'h0 : PRFFreeList_3; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_277 = 6'h4 == rs1Addr ? 1'h0 : PRFFreeList_4; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_278 = 6'h5 == rs1Addr ? 1'h0 : PRFFreeList_5; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_279 = 6'h6 == rs1Addr ? 1'h0 : PRFFreeList_6; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_280 = 6'h7 == rs1Addr ? 1'h0 : PRFFreeList_7; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_281 = 6'h8 == rs1Addr ? 1'h0 : PRFFreeList_8; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_282 = 6'h9 == rs1Addr ? 1'h0 : PRFFreeList_9; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_283 = 6'ha == rs1Addr ? 1'h0 : PRFFreeList_10; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_284 = 6'hb == rs1Addr ? 1'h0 : PRFFreeList_11; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_285 = 6'hc == rs1Addr ? 1'h0 : PRFFreeList_12; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_286 = 6'hd == rs1Addr ? 1'h0 : PRFFreeList_13; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_287 = 6'he == rs1Addr ? 1'h0 : PRFFreeList_14; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_288 = 6'hf == rs1Addr ? 1'h0 : PRFFreeList_15; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_289 = 6'h10 == rs1Addr ? 1'h0 : PRFFreeList_16; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_290 = 6'h11 == rs1Addr ? 1'h0 : PRFFreeList_17; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_291 = 6'h12 == rs1Addr ? 1'h0 : PRFFreeList_18; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_292 = 6'h13 == rs1Addr ? 1'h0 : PRFFreeList_19; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_293 = 6'h14 == rs1Addr ? 1'h0 : PRFFreeList_20; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_294 = 6'h15 == rs1Addr ? 1'h0 : PRFFreeList_21; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_295 = 6'h16 == rs1Addr ? 1'h0 : PRFFreeList_22; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_296 = 6'h17 == rs1Addr ? 1'h0 : PRFFreeList_23; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_297 = 6'h18 == rs1Addr ? 1'h0 : PRFFreeList_24; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_298 = 6'h19 == rs1Addr ? 1'h0 : PRFFreeList_25; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_299 = 6'h1a == rs1Addr ? 1'h0 : PRFFreeList_26; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_300 = 6'h1b == rs1Addr ? 1'h0 : PRFFreeList_27; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_301 = 6'h1c == rs1Addr ? 1'h0 : PRFFreeList_28; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_302 = 6'h1d == rs1Addr ? 1'h0 : PRFFreeList_29; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_303 = 6'h1e == rs1Addr ? 1'h0 : PRFFreeList_30; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_304 = 6'h1f == rs1Addr ? 1'h0 : PRFFreeList_31; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_305 = 6'h20 == rs1Addr ? 1'h0 : PRFFreeList_32; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_306 = 6'h21 == rs1Addr ? 1'h0 : PRFFreeList_33; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_307 = 6'h22 == rs1Addr ? 1'h0 : PRFFreeList_34; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_308 = 6'h23 == rs1Addr ? 1'h0 : PRFFreeList_35; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_309 = 6'h24 == rs1Addr ? 1'h0 : PRFFreeList_36; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_310 = 6'h25 == rs1Addr ? 1'h0 : PRFFreeList_37; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_311 = 6'h26 == rs1Addr ? 1'h0 : PRFFreeList_38; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_312 = 6'h27 == rs1Addr ? 1'h0 : PRFFreeList_39; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_313 = 6'h28 == rs1Addr ? 1'h0 : PRFFreeList_40; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_314 = 6'h29 == rs1Addr ? 1'h0 : PRFFreeList_41; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_315 = 6'h2a == rs1Addr ? 1'h0 : PRFFreeList_42; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_316 = 6'h2b == rs1Addr ? 1'h0 : PRFFreeList_43; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_317 = 6'h2c == rs1Addr ? 1'h0 : PRFFreeList_44; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_318 = 6'h2d == rs1Addr ? 1'h0 : PRFFreeList_45; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_319 = 6'h2e == rs1Addr ? 1'h0 : PRFFreeList_46; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_320 = 6'h2f == rs1Addr ? 1'h0 : PRFFreeList_47; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_321 = 6'h30 == rs1Addr ? 1'h0 : PRFFreeList_48; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_322 = 6'h31 == rs1Addr ? 1'h0 : PRFFreeList_49; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_323 = 6'h32 == rs1Addr ? 1'h0 : PRFFreeList_50; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_324 = 6'h33 == rs1Addr ? 1'h0 : PRFFreeList_51; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_325 = 6'h34 == rs1Addr ? 1'h0 : PRFFreeList_52; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_326 = 6'h35 == rs1Addr ? 1'h0 : PRFFreeList_53; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_327 = 6'h36 == rs1Addr ? 1'h0 : PRFFreeList_54; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_328 = 6'h37 == rs1Addr ? 1'h0 : PRFFreeList_55; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_329 = 6'h38 == rs1Addr ? 1'h0 : PRFFreeList_56; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_330 = 6'h39 == rs1Addr ? 1'h0 : PRFFreeList_57; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_331 = 6'h3a == rs1Addr ? 1'h0 : PRFFreeList_58; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_332 = 6'h3b == rs1Addr ? 1'h0 : PRFFreeList_59; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_333 = 6'h3c == rs1Addr ? 1'h0 : PRFFreeList_60; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_334 = 6'h3d == rs1Addr ? 1'h0 : PRFFreeList_61; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_335 = 6'h3e == rs1Addr ? 1'h0 : PRFFreeList_62; // @[decode.scala 336:{28,28} 303:36]
  wire  _GEN_337 = 6'h0 == rs2Addr ? 1'h0 : PRFFreeList_0; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_338 = 6'h1 == rs2Addr ? 1'h0 : PRFFreeList_1; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_339 = 6'h2 == rs2Addr ? 1'h0 : PRFFreeList_2; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_340 = 6'h3 == rs2Addr ? 1'h0 : PRFFreeList_3; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_341 = 6'h4 == rs2Addr ? 1'h0 : PRFFreeList_4; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_342 = 6'h5 == rs2Addr ? 1'h0 : PRFFreeList_5; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_343 = 6'h6 == rs2Addr ? 1'h0 : PRFFreeList_6; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_344 = 6'h7 == rs2Addr ? 1'h0 : PRFFreeList_7; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_345 = 6'h8 == rs2Addr ? 1'h0 : PRFFreeList_8; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_346 = 6'h9 == rs2Addr ? 1'h0 : PRFFreeList_9; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_347 = 6'ha == rs2Addr ? 1'h0 : PRFFreeList_10; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_348 = 6'hb == rs2Addr ? 1'h0 : PRFFreeList_11; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_349 = 6'hc == rs2Addr ? 1'h0 : PRFFreeList_12; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_350 = 6'hd == rs2Addr ? 1'h0 : PRFFreeList_13; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_351 = 6'he == rs2Addr ? 1'h0 : PRFFreeList_14; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_352 = 6'hf == rs2Addr ? 1'h0 : PRFFreeList_15; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_353 = 6'h10 == rs2Addr ? 1'h0 : PRFFreeList_16; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_354 = 6'h11 == rs2Addr ? 1'h0 : PRFFreeList_17; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_355 = 6'h12 == rs2Addr ? 1'h0 : PRFFreeList_18; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_356 = 6'h13 == rs2Addr ? 1'h0 : PRFFreeList_19; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_357 = 6'h14 == rs2Addr ? 1'h0 : PRFFreeList_20; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_358 = 6'h15 == rs2Addr ? 1'h0 : PRFFreeList_21; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_359 = 6'h16 == rs2Addr ? 1'h0 : PRFFreeList_22; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_360 = 6'h17 == rs2Addr ? 1'h0 : PRFFreeList_23; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_361 = 6'h18 == rs2Addr ? 1'h0 : PRFFreeList_24; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_362 = 6'h19 == rs2Addr ? 1'h0 : PRFFreeList_25; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_363 = 6'h1a == rs2Addr ? 1'h0 : PRFFreeList_26; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_364 = 6'h1b == rs2Addr ? 1'h0 : PRFFreeList_27; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_365 = 6'h1c == rs2Addr ? 1'h0 : PRFFreeList_28; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_366 = 6'h1d == rs2Addr ? 1'h0 : PRFFreeList_29; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_367 = 6'h1e == rs2Addr ? 1'h0 : PRFFreeList_30; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_368 = 6'h1f == rs2Addr ? 1'h0 : PRFFreeList_31; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_369 = 6'h20 == rs2Addr ? 1'h0 : PRFFreeList_32; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_370 = 6'h21 == rs2Addr ? 1'h0 : PRFFreeList_33; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_371 = 6'h22 == rs2Addr ? 1'h0 : PRFFreeList_34; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_372 = 6'h23 == rs2Addr ? 1'h0 : PRFFreeList_35; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_373 = 6'h24 == rs2Addr ? 1'h0 : PRFFreeList_36; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_374 = 6'h25 == rs2Addr ? 1'h0 : PRFFreeList_37; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_375 = 6'h26 == rs2Addr ? 1'h0 : PRFFreeList_38; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_376 = 6'h27 == rs2Addr ? 1'h0 : PRFFreeList_39; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_377 = 6'h28 == rs2Addr ? 1'h0 : PRFFreeList_40; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_378 = 6'h29 == rs2Addr ? 1'h0 : PRFFreeList_41; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_379 = 6'h2a == rs2Addr ? 1'h0 : PRFFreeList_42; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_380 = 6'h2b == rs2Addr ? 1'h0 : PRFFreeList_43; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_381 = 6'h2c == rs2Addr ? 1'h0 : PRFFreeList_44; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_382 = 6'h2d == rs2Addr ? 1'h0 : PRFFreeList_45; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_383 = 6'h2e == rs2Addr ? 1'h0 : PRFFreeList_46; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_384 = 6'h2f == rs2Addr ? 1'h0 : PRFFreeList_47; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_385 = 6'h30 == rs2Addr ? 1'h0 : PRFFreeList_48; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_386 = 6'h31 == rs2Addr ? 1'h0 : PRFFreeList_49; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_387 = 6'h32 == rs2Addr ? 1'h0 : PRFFreeList_50; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_388 = 6'h33 == rs2Addr ? 1'h0 : PRFFreeList_51; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_389 = 6'h34 == rs2Addr ? 1'h0 : PRFFreeList_52; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_390 = 6'h35 == rs2Addr ? 1'h0 : PRFFreeList_53; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_391 = 6'h36 == rs2Addr ? 1'h0 : PRFFreeList_54; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_392 = 6'h37 == rs2Addr ? 1'h0 : PRFFreeList_55; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_393 = 6'h38 == rs2Addr ? 1'h0 : PRFFreeList_56; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_394 = 6'h39 == rs2Addr ? 1'h0 : PRFFreeList_57; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_395 = 6'h3a == rs2Addr ? 1'h0 : PRFFreeList_58; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_396 = 6'h3b == rs2Addr ? 1'h0 : PRFFreeList_59; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_397 = 6'h3c == rs2Addr ? 1'h0 : PRFFreeList_60; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_398 = 6'h3d == rs2Addr ? 1'h0 : PRFFreeList_61; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_399 = 6'h3e == rs2Addr ? 1'h0 : PRFFreeList_62; // @[decode.scala 338:{28,28} 303:36]
  wire  _GEN_401 = _T_20 ? _GEN_337 : PRFFreeList_0; // @[decode.scala 303:36 337:41]
  wire  _GEN_402 = _T_20 ? _GEN_338 : PRFFreeList_1; // @[decode.scala 303:36 337:41]
  wire  _GEN_403 = _T_20 ? _GEN_339 : PRFFreeList_2; // @[decode.scala 303:36 337:41]
  wire  _GEN_404 = _T_20 ? _GEN_340 : PRFFreeList_3; // @[decode.scala 303:36 337:41]
  wire  _GEN_405 = _T_20 ? _GEN_341 : PRFFreeList_4; // @[decode.scala 303:36 337:41]
  wire  _GEN_406 = _T_20 ? _GEN_342 : PRFFreeList_5; // @[decode.scala 303:36 337:41]
  wire  _GEN_407 = _T_20 ? _GEN_343 : PRFFreeList_6; // @[decode.scala 303:36 337:41]
  wire  _GEN_408 = _T_20 ? _GEN_344 : PRFFreeList_7; // @[decode.scala 303:36 337:41]
  wire  _GEN_409 = _T_20 ? _GEN_345 : PRFFreeList_8; // @[decode.scala 303:36 337:41]
  wire  _GEN_410 = _T_20 ? _GEN_346 : PRFFreeList_9; // @[decode.scala 303:36 337:41]
  wire  _GEN_411 = _T_20 ? _GEN_347 : PRFFreeList_10; // @[decode.scala 303:36 337:41]
  wire  _GEN_412 = _T_20 ? _GEN_348 : PRFFreeList_11; // @[decode.scala 303:36 337:41]
  wire  _GEN_413 = _T_20 ? _GEN_349 : PRFFreeList_12; // @[decode.scala 303:36 337:41]
  wire  _GEN_414 = _T_20 ? _GEN_350 : PRFFreeList_13; // @[decode.scala 303:36 337:41]
  wire  _GEN_415 = _T_20 ? _GEN_351 : PRFFreeList_14; // @[decode.scala 303:36 337:41]
  wire  _GEN_416 = _T_20 ? _GEN_352 : PRFFreeList_15; // @[decode.scala 303:36 337:41]
  wire  _GEN_417 = _T_20 ? _GEN_353 : PRFFreeList_16; // @[decode.scala 303:36 337:41]
  wire  _GEN_418 = _T_20 ? _GEN_354 : PRFFreeList_17; // @[decode.scala 303:36 337:41]
  wire  _GEN_419 = _T_20 ? _GEN_355 : PRFFreeList_18; // @[decode.scala 303:36 337:41]
  wire  _GEN_420 = _T_20 ? _GEN_356 : PRFFreeList_19; // @[decode.scala 303:36 337:41]
  wire  _GEN_421 = _T_20 ? _GEN_357 : PRFFreeList_20; // @[decode.scala 303:36 337:41]
  wire  _GEN_422 = _T_20 ? _GEN_358 : PRFFreeList_21; // @[decode.scala 303:36 337:41]
  wire  _GEN_423 = _T_20 ? _GEN_359 : PRFFreeList_22; // @[decode.scala 303:36 337:41]
  wire  _GEN_424 = _T_20 ? _GEN_360 : PRFFreeList_23; // @[decode.scala 303:36 337:41]
  wire  _GEN_425 = _T_20 ? _GEN_361 : PRFFreeList_24; // @[decode.scala 303:36 337:41]
  wire  _GEN_426 = _T_20 ? _GEN_362 : PRFFreeList_25; // @[decode.scala 303:36 337:41]
  wire  _GEN_427 = _T_20 ? _GEN_363 : PRFFreeList_26; // @[decode.scala 303:36 337:41]
  wire  _GEN_428 = _T_20 ? _GEN_364 : PRFFreeList_27; // @[decode.scala 303:36 337:41]
  wire  _GEN_429 = _T_20 ? _GEN_365 : PRFFreeList_28; // @[decode.scala 303:36 337:41]
  wire  _GEN_430 = _T_20 ? _GEN_366 : PRFFreeList_29; // @[decode.scala 303:36 337:41]
  wire  _GEN_431 = _T_20 ? _GEN_367 : PRFFreeList_30; // @[decode.scala 303:36 337:41]
  wire  _GEN_432 = _T_20 ? _GEN_368 : PRFFreeList_31; // @[decode.scala 303:36 337:41]
  wire  _GEN_433 = _T_20 ? _GEN_369 : PRFFreeList_32; // @[decode.scala 303:36 337:41]
  wire  _GEN_434 = _T_20 ? _GEN_370 : PRFFreeList_33; // @[decode.scala 303:36 337:41]
  wire  _GEN_435 = _T_20 ? _GEN_371 : PRFFreeList_34; // @[decode.scala 303:36 337:41]
  wire  _GEN_436 = _T_20 ? _GEN_372 : PRFFreeList_35; // @[decode.scala 303:36 337:41]
  wire  _GEN_437 = _T_20 ? _GEN_373 : PRFFreeList_36; // @[decode.scala 303:36 337:41]
  wire  _GEN_438 = _T_20 ? _GEN_374 : PRFFreeList_37; // @[decode.scala 303:36 337:41]
  wire  _GEN_439 = _T_20 ? _GEN_375 : PRFFreeList_38; // @[decode.scala 303:36 337:41]
  wire  _GEN_440 = _T_20 ? _GEN_376 : PRFFreeList_39; // @[decode.scala 303:36 337:41]
  wire  _GEN_441 = _T_20 ? _GEN_377 : PRFFreeList_40; // @[decode.scala 303:36 337:41]
  wire  _GEN_442 = _T_20 ? _GEN_378 : PRFFreeList_41; // @[decode.scala 303:36 337:41]
  wire  _GEN_443 = _T_20 ? _GEN_379 : PRFFreeList_42; // @[decode.scala 303:36 337:41]
  wire  _GEN_444 = _T_20 ? _GEN_380 : PRFFreeList_43; // @[decode.scala 303:36 337:41]
  wire  _GEN_445 = _T_20 ? _GEN_381 : PRFFreeList_44; // @[decode.scala 303:36 337:41]
  wire  _GEN_446 = _T_20 ? _GEN_382 : PRFFreeList_45; // @[decode.scala 303:36 337:41]
  wire  _GEN_447 = _T_20 ? _GEN_383 : PRFFreeList_46; // @[decode.scala 303:36 337:41]
  wire  _GEN_448 = _T_20 ? _GEN_384 : PRFFreeList_47; // @[decode.scala 303:36 337:41]
  wire  _GEN_449 = _T_20 ? _GEN_385 : PRFFreeList_48; // @[decode.scala 303:36 337:41]
  wire  _GEN_450 = _T_20 ? _GEN_386 : PRFFreeList_49; // @[decode.scala 303:36 337:41]
  wire  _GEN_451 = _T_20 ? _GEN_387 : PRFFreeList_50; // @[decode.scala 303:36 337:41]
  wire  _GEN_452 = _T_20 ? _GEN_388 : PRFFreeList_51; // @[decode.scala 303:36 337:41]
  wire  _GEN_453 = _T_20 ? _GEN_389 : PRFFreeList_52; // @[decode.scala 303:36 337:41]
  wire  _GEN_454 = _T_20 ? _GEN_390 : PRFFreeList_53; // @[decode.scala 303:36 337:41]
  wire  _GEN_455 = _T_20 ? _GEN_391 : PRFFreeList_54; // @[decode.scala 303:36 337:41]
  wire  _GEN_456 = _T_20 ? _GEN_392 : PRFFreeList_55; // @[decode.scala 303:36 337:41]
  wire  _GEN_457 = _T_20 ? _GEN_393 : PRFFreeList_56; // @[decode.scala 303:36 337:41]
  wire  _GEN_458 = _T_20 ? _GEN_394 : PRFFreeList_57; // @[decode.scala 303:36 337:41]
  wire  _GEN_459 = _T_20 ? _GEN_395 : PRFFreeList_58; // @[decode.scala 303:36 337:41]
  wire  _GEN_460 = _T_20 ? _GEN_396 : PRFFreeList_59; // @[decode.scala 303:36 337:41]
  wire  _GEN_461 = _T_20 ? _GEN_397 : PRFFreeList_60; // @[decode.scala 303:36 337:41]
  wire  _GEN_462 = _T_20 ? _GEN_398 : PRFFreeList_61; // @[decode.scala 303:36 337:41]
  wire  _GEN_463 = _T_20 ? _GEN_399 : PRFFreeList_62; // @[decode.scala 303:36 337:41]
  wire  _GEN_465 = _T_19 ? _GEN_273 : _GEN_401; // @[decode.scala 335:35]
  wire  _GEN_466 = _T_19 ? _GEN_274 : _GEN_402; // @[decode.scala 335:35]
  wire  _GEN_467 = _T_19 ? _GEN_275 : _GEN_403; // @[decode.scala 335:35]
  wire  _GEN_468 = _T_19 ? _GEN_276 : _GEN_404; // @[decode.scala 335:35]
  wire  _GEN_469 = _T_19 ? _GEN_277 : _GEN_405; // @[decode.scala 335:35]
  wire  _GEN_470 = _T_19 ? _GEN_278 : _GEN_406; // @[decode.scala 335:35]
  wire  _GEN_471 = _T_19 ? _GEN_279 : _GEN_407; // @[decode.scala 335:35]
  wire  _GEN_472 = _T_19 ? _GEN_280 : _GEN_408; // @[decode.scala 335:35]
  wire  _GEN_473 = _T_19 ? _GEN_281 : _GEN_409; // @[decode.scala 335:35]
  wire  _GEN_474 = _T_19 ? _GEN_282 : _GEN_410; // @[decode.scala 335:35]
  wire  _GEN_475 = _T_19 ? _GEN_283 : _GEN_411; // @[decode.scala 335:35]
  wire  _GEN_476 = _T_19 ? _GEN_284 : _GEN_412; // @[decode.scala 335:35]
  wire  _GEN_477 = _T_19 ? _GEN_285 : _GEN_413; // @[decode.scala 335:35]
  wire  _GEN_478 = _T_19 ? _GEN_286 : _GEN_414; // @[decode.scala 335:35]
  wire  _GEN_479 = _T_19 ? _GEN_287 : _GEN_415; // @[decode.scala 335:35]
  wire  _GEN_480 = _T_19 ? _GEN_288 : _GEN_416; // @[decode.scala 335:35]
  wire  _GEN_481 = _T_19 ? _GEN_289 : _GEN_417; // @[decode.scala 335:35]
  wire  _GEN_482 = _T_19 ? _GEN_290 : _GEN_418; // @[decode.scala 335:35]
  wire  _GEN_483 = _T_19 ? _GEN_291 : _GEN_419; // @[decode.scala 335:35]
  wire  _GEN_484 = _T_19 ? _GEN_292 : _GEN_420; // @[decode.scala 335:35]
  wire  _GEN_485 = _T_19 ? _GEN_293 : _GEN_421; // @[decode.scala 335:35]
  wire  _GEN_486 = _T_19 ? _GEN_294 : _GEN_422; // @[decode.scala 335:35]
  wire  _GEN_487 = _T_19 ? _GEN_295 : _GEN_423; // @[decode.scala 335:35]
  wire  _GEN_488 = _T_19 ? _GEN_296 : _GEN_424; // @[decode.scala 335:35]
  wire  _GEN_489 = _T_19 ? _GEN_297 : _GEN_425; // @[decode.scala 335:35]
  wire  _GEN_490 = _T_19 ? _GEN_298 : _GEN_426; // @[decode.scala 335:35]
  wire  _GEN_491 = _T_19 ? _GEN_299 : _GEN_427; // @[decode.scala 335:35]
  wire  _GEN_492 = _T_19 ? _GEN_300 : _GEN_428; // @[decode.scala 335:35]
  wire  _GEN_493 = _T_19 ? _GEN_301 : _GEN_429; // @[decode.scala 335:35]
  wire  _GEN_494 = _T_19 ? _GEN_302 : _GEN_430; // @[decode.scala 335:35]
  wire  _GEN_495 = _T_19 ? _GEN_303 : _GEN_431; // @[decode.scala 335:35]
  wire  _GEN_496 = _T_19 ? _GEN_304 : _GEN_432; // @[decode.scala 335:35]
  wire  _GEN_497 = _T_19 ? _GEN_305 : _GEN_433; // @[decode.scala 335:35]
  wire  _GEN_498 = _T_19 ? _GEN_306 : _GEN_434; // @[decode.scala 335:35]
  wire  _GEN_499 = _T_19 ? _GEN_307 : _GEN_435; // @[decode.scala 335:35]
  wire  _GEN_500 = _T_19 ? _GEN_308 : _GEN_436; // @[decode.scala 335:35]
  wire  _GEN_501 = _T_19 ? _GEN_309 : _GEN_437; // @[decode.scala 335:35]
  wire  _GEN_502 = _T_19 ? _GEN_310 : _GEN_438; // @[decode.scala 335:35]
  wire  _GEN_503 = _T_19 ? _GEN_311 : _GEN_439; // @[decode.scala 335:35]
  wire  _GEN_504 = _T_19 ? _GEN_312 : _GEN_440; // @[decode.scala 335:35]
  wire  _GEN_505 = _T_19 ? _GEN_313 : _GEN_441; // @[decode.scala 335:35]
  wire  _GEN_506 = _T_19 ? _GEN_314 : _GEN_442; // @[decode.scala 335:35]
  wire  _GEN_507 = _T_19 ? _GEN_315 : _GEN_443; // @[decode.scala 335:35]
  wire  _GEN_508 = _T_19 ? _GEN_316 : _GEN_444; // @[decode.scala 335:35]
  wire  _GEN_509 = _T_19 ? _GEN_317 : _GEN_445; // @[decode.scala 335:35]
  wire  _GEN_510 = _T_19 ? _GEN_318 : _GEN_446; // @[decode.scala 335:35]
  wire  _GEN_511 = _T_19 ? _GEN_319 : _GEN_447; // @[decode.scala 335:35]
  wire  _GEN_512 = _T_19 ? _GEN_320 : _GEN_448; // @[decode.scala 335:35]
  wire  _GEN_513 = _T_19 ? _GEN_321 : _GEN_449; // @[decode.scala 335:35]
  wire  _GEN_514 = _T_19 ? _GEN_322 : _GEN_450; // @[decode.scala 335:35]
  wire  _GEN_515 = _T_19 ? _GEN_323 : _GEN_451; // @[decode.scala 335:35]
  wire  _GEN_516 = _T_19 ? _GEN_324 : _GEN_452; // @[decode.scala 335:35]
  wire  _GEN_517 = _T_19 ? _GEN_325 : _GEN_453; // @[decode.scala 335:35]
  wire  _GEN_518 = _T_19 ? _GEN_326 : _GEN_454; // @[decode.scala 335:35]
  wire  _GEN_519 = _T_19 ? _GEN_327 : _GEN_455; // @[decode.scala 335:35]
  wire  _GEN_520 = _T_19 ? _GEN_328 : _GEN_456; // @[decode.scala 335:35]
  wire  _GEN_521 = _T_19 ? _GEN_329 : _GEN_457; // @[decode.scala 335:35]
  wire  _GEN_522 = _T_19 ? _GEN_330 : _GEN_458; // @[decode.scala 335:35]
  wire  _GEN_523 = _T_19 ? _GEN_331 : _GEN_459; // @[decode.scala 335:35]
  wire  _GEN_524 = _T_19 ? _GEN_332 : _GEN_460; // @[decode.scala 335:35]
  wire  _GEN_525 = _T_19 ? _GEN_333 : _GEN_461; // @[decode.scala 335:35]
  wire  _GEN_526 = _T_19 ? _GEN_334 : _GEN_462; // @[decode.scala 335:35]
  wire  _GEN_527 = _T_19 ? _GEN_335 : _GEN_463; // @[decode.scala 335:35]
  wire  _GEN_530 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_465 : PRFFreeList_0; // @[decode.scala 303:36 333:60]
  wire  _GEN_531 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_466 : PRFFreeList_1; // @[decode.scala 303:36 333:60]
  wire  _GEN_532 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_467 : PRFFreeList_2; // @[decode.scala 303:36 333:60]
  wire  _GEN_533 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_468 : PRFFreeList_3; // @[decode.scala 303:36 333:60]
  wire  _GEN_534 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_469 : PRFFreeList_4; // @[decode.scala 303:36 333:60]
  wire  _GEN_535 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_470 : PRFFreeList_5; // @[decode.scala 303:36 333:60]
  wire  _GEN_536 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_471 : PRFFreeList_6; // @[decode.scala 303:36 333:60]
  wire  _GEN_537 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_472 : PRFFreeList_7; // @[decode.scala 303:36 333:60]
  wire  _GEN_538 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_473 : PRFFreeList_8; // @[decode.scala 303:36 333:60]
  wire  _GEN_539 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_474 : PRFFreeList_9; // @[decode.scala 303:36 333:60]
  wire  _GEN_540 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_475 : PRFFreeList_10; // @[decode.scala 303:36 333:60]
  wire  _GEN_541 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_476 : PRFFreeList_11; // @[decode.scala 303:36 333:60]
  wire  _GEN_542 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_477 : PRFFreeList_12; // @[decode.scala 303:36 333:60]
  wire  _GEN_543 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_478 : PRFFreeList_13; // @[decode.scala 303:36 333:60]
  wire  _GEN_544 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_479 : PRFFreeList_14; // @[decode.scala 303:36 333:60]
  wire  _GEN_545 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_480 : PRFFreeList_15; // @[decode.scala 303:36 333:60]
  wire  _GEN_546 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_481 : PRFFreeList_16; // @[decode.scala 303:36 333:60]
  wire  _GEN_547 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_482 : PRFFreeList_17; // @[decode.scala 303:36 333:60]
  wire  _GEN_548 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_483 : PRFFreeList_18; // @[decode.scala 303:36 333:60]
  wire  _GEN_549 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_484 : PRFFreeList_19; // @[decode.scala 303:36 333:60]
  wire  _GEN_550 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_485 : PRFFreeList_20; // @[decode.scala 303:36 333:60]
  wire  _GEN_551 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_486 : PRFFreeList_21; // @[decode.scala 303:36 333:60]
  wire  _GEN_552 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_487 : PRFFreeList_22; // @[decode.scala 303:36 333:60]
  wire  _GEN_553 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_488 : PRFFreeList_23; // @[decode.scala 303:36 333:60]
  wire  _GEN_554 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_489 : PRFFreeList_24; // @[decode.scala 303:36 333:60]
  wire  _GEN_555 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_490 : PRFFreeList_25; // @[decode.scala 303:36 333:60]
  wire  _GEN_556 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_491 : PRFFreeList_26; // @[decode.scala 303:36 333:60]
  wire  _GEN_557 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_492 : PRFFreeList_27; // @[decode.scala 303:36 333:60]
  wire  _GEN_558 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_493 : PRFFreeList_28; // @[decode.scala 303:36 333:60]
  wire  _GEN_559 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_494 : PRFFreeList_29; // @[decode.scala 303:36 333:60]
  wire  _GEN_560 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_495 : PRFFreeList_30; // @[decode.scala 303:36 333:60]
  wire  _GEN_561 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_496 : PRFFreeList_31; // @[decode.scala 303:36 333:60]
  wire  _GEN_562 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_497 : PRFFreeList_32; // @[decode.scala 303:36 333:60]
  wire  _GEN_563 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_498 : PRFFreeList_33; // @[decode.scala 303:36 333:60]
  wire  _GEN_564 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_499 : PRFFreeList_34; // @[decode.scala 303:36 333:60]
  wire  _GEN_565 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_500 : PRFFreeList_35; // @[decode.scala 303:36 333:60]
  wire  _GEN_566 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_501 : PRFFreeList_36; // @[decode.scala 303:36 333:60]
  wire  _GEN_567 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_502 : PRFFreeList_37; // @[decode.scala 303:36 333:60]
  wire  _GEN_568 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_503 : PRFFreeList_38; // @[decode.scala 303:36 333:60]
  wire  _GEN_569 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_504 : PRFFreeList_39; // @[decode.scala 303:36 333:60]
  wire  _GEN_570 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_505 : PRFFreeList_40; // @[decode.scala 303:36 333:60]
  wire  _GEN_571 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_506 : PRFFreeList_41; // @[decode.scala 303:36 333:60]
  wire  _GEN_572 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_507 : PRFFreeList_42; // @[decode.scala 303:36 333:60]
  wire  _GEN_573 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_508 : PRFFreeList_43; // @[decode.scala 303:36 333:60]
  wire  _GEN_574 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_509 : PRFFreeList_44; // @[decode.scala 303:36 333:60]
  wire  _GEN_575 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_510 : PRFFreeList_45; // @[decode.scala 303:36 333:60]
  wire  _GEN_576 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_511 : PRFFreeList_46; // @[decode.scala 303:36 333:60]
  wire  _GEN_577 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_512 : PRFFreeList_47; // @[decode.scala 303:36 333:60]
  wire  _GEN_578 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_513 : PRFFreeList_48; // @[decode.scala 303:36 333:60]
  wire  _GEN_579 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_514 : PRFFreeList_49; // @[decode.scala 303:36 333:60]
  wire  _GEN_580 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_515 : PRFFreeList_50; // @[decode.scala 303:36 333:60]
  wire  _GEN_581 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_516 : PRFFreeList_51; // @[decode.scala 303:36 333:60]
  wire  _GEN_582 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_517 : PRFFreeList_52; // @[decode.scala 303:36 333:60]
  wire  _GEN_583 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_518 : PRFFreeList_53; // @[decode.scala 303:36 333:60]
  wire  _GEN_584 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_519 : PRFFreeList_54; // @[decode.scala 303:36 333:60]
  wire  _GEN_585 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_520 : PRFFreeList_55; // @[decode.scala 303:36 333:60]
  wire  _GEN_586 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_521 : PRFFreeList_56; // @[decode.scala 303:36 333:60]
  wire  _GEN_587 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_522 : PRFFreeList_57; // @[decode.scala 303:36 333:60]
  wire  _GEN_588 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_523 : PRFFreeList_58; // @[decode.scala 303:36 333:60]
  wire  _GEN_589 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_524 : PRFFreeList_59; // @[decode.scala 303:36 333:60]
  wire  _GEN_590 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_525 : PRFFreeList_60; // @[decode.scala 303:36 333:60]
  wire  _GEN_591 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_526 : PRFFreeList_61; // @[decode.scala 303:36 333:60]
  wire  _GEN_592 = rs1Addr == freeRegAddr | rs2Addr == freeRegAddr ? _GEN_527 : PRFFreeList_62; // @[decode.scala 303:36 333:60]
  wire  _GEN_658 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h0 == outputBuffer_PRFDest |
    PRFValidList_0 : PRFValidList_0; // @[decode.scala 193:29 342:71]
  wire  _GEN_659 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h1 == outputBuffer_PRFDest |
    PRFValidList_1 : PRFValidList_1; // @[decode.scala 193:29 342:71]
  wire  _GEN_660 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h2 == outputBuffer_PRFDest |
    PRFValidList_2 : PRFValidList_2; // @[decode.scala 193:29 342:71]
  wire  _GEN_661 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h3 == outputBuffer_PRFDest |
    PRFValidList_3 : PRFValidList_3; // @[decode.scala 193:29 342:71]
  wire  _GEN_662 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h4 == outputBuffer_PRFDest |
    PRFValidList_4 : PRFValidList_4; // @[decode.scala 193:29 342:71]
  wire  _GEN_663 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h5 == outputBuffer_PRFDest |
    PRFValidList_5 : PRFValidList_5; // @[decode.scala 193:29 342:71]
  wire  _GEN_664 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h6 == outputBuffer_PRFDest |
    PRFValidList_6 : PRFValidList_6; // @[decode.scala 193:29 342:71]
  wire  _GEN_665 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h7 == outputBuffer_PRFDest |
    PRFValidList_7 : PRFValidList_7; // @[decode.scala 193:29 342:71]
  wire  _GEN_666 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h8 == outputBuffer_PRFDest |
    PRFValidList_8 : PRFValidList_8; // @[decode.scala 193:29 342:71]
  wire  _GEN_667 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h9 == outputBuffer_PRFDest |
    PRFValidList_9 : PRFValidList_9; // @[decode.scala 193:29 342:71]
  wire  _GEN_668 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'ha == outputBuffer_PRFDest |
    PRFValidList_10 : PRFValidList_10; // @[decode.scala 193:29 342:71]
  wire  _GEN_669 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'hb == outputBuffer_PRFDest |
    PRFValidList_11 : PRFValidList_11; // @[decode.scala 193:29 342:71]
  wire  _GEN_670 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'hc == outputBuffer_PRFDest |
    PRFValidList_12 : PRFValidList_12; // @[decode.scala 193:29 342:71]
  wire  _GEN_671 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'hd == outputBuffer_PRFDest |
    PRFValidList_13 : PRFValidList_13; // @[decode.scala 193:29 342:71]
  wire  _GEN_672 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'he == outputBuffer_PRFDest |
    PRFValidList_14 : PRFValidList_14; // @[decode.scala 193:29 342:71]
  wire  _GEN_673 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'hf == outputBuffer_PRFDest |
    PRFValidList_15 : PRFValidList_15; // @[decode.scala 193:29 342:71]
  wire  _GEN_674 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h10 == outputBuffer_PRFDest |
    PRFValidList_16 : PRFValidList_16; // @[decode.scala 193:29 342:71]
  wire  _GEN_675 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h11 == outputBuffer_PRFDest |
    PRFValidList_17 : PRFValidList_17; // @[decode.scala 193:29 342:71]
  wire  _GEN_676 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h12 == outputBuffer_PRFDest |
    PRFValidList_18 : PRFValidList_18; // @[decode.scala 193:29 342:71]
  wire  _GEN_677 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h13 == outputBuffer_PRFDest |
    PRFValidList_19 : PRFValidList_19; // @[decode.scala 193:29 342:71]
  wire  _GEN_678 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h14 == outputBuffer_PRFDest |
    PRFValidList_20 : PRFValidList_20; // @[decode.scala 193:29 342:71]
  wire  _GEN_679 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h15 == outputBuffer_PRFDest |
    PRFValidList_21 : PRFValidList_21; // @[decode.scala 193:29 342:71]
  wire  _GEN_680 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h16 == outputBuffer_PRFDest |
    PRFValidList_22 : PRFValidList_22; // @[decode.scala 193:29 342:71]
  wire  _GEN_681 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h17 == outputBuffer_PRFDest |
    PRFValidList_23 : PRFValidList_23; // @[decode.scala 193:29 342:71]
  wire  _GEN_682 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h18 == outputBuffer_PRFDest |
    PRFValidList_24 : PRFValidList_24; // @[decode.scala 193:29 342:71]
  wire  _GEN_683 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h19 == outputBuffer_PRFDest |
    PRFValidList_25 : PRFValidList_25; // @[decode.scala 193:29 342:71]
  wire  _GEN_684 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h1a == outputBuffer_PRFDest |
    PRFValidList_26 : PRFValidList_26; // @[decode.scala 193:29 342:71]
  wire  _GEN_685 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h1b == outputBuffer_PRFDest |
    PRFValidList_27 : PRFValidList_27; // @[decode.scala 193:29 342:71]
  wire  _GEN_686 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h1c == outputBuffer_PRFDest |
    PRFValidList_28 : PRFValidList_28; // @[decode.scala 193:29 342:71]
  wire  _GEN_687 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h1d == outputBuffer_PRFDest |
    PRFValidList_29 : PRFValidList_29; // @[decode.scala 193:29 342:71]
  wire  _GEN_688 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h1e == outputBuffer_PRFDest |
    PRFValidList_30 : PRFValidList_30; // @[decode.scala 193:29 342:71]
  wire  _GEN_689 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h1f == outputBuffer_PRFDest |
    PRFValidList_31 : PRFValidList_31; // @[decode.scala 193:29 342:71]
  wire  _GEN_690 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h20 == outputBuffer_PRFDest |
    PRFValidList_32 : PRFValidList_32; // @[decode.scala 193:29 342:71]
  wire  _GEN_691 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h21 == outputBuffer_PRFDest |
    PRFValidList_33 : PRFValidList_33; // @[decode.scala 193:29 342:71]
  wire  _GEN_692 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h22 == outputBuffer_PRFDest |
    PRFValidList_34 : PRFValidList_34; // @[decode.scala 193:29 342:71]
  wire  _GEN_693 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h23 == outputBuffer_PRFDest |
    PRFValidList_35 : PRFValidList_35; // @[decode.scala 193:29 342:71]
  wire  _GEN_694 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h24 == outputBuffer_PRFDest |
    PRFValidList_36 : PRFValidList_36; // @[decode.scala 193:29 342:71]
  wire  _GEN_695 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h25 == outputBuffer_PRFDest |
    PRFValidList_37 : PRFValidList_37; // @[decode.scala 193:29 342:71]
  wire  _GEN_696 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h26 == outputBuffer_PRFDest |
    PRFValidList_38 : PRFValidList_38; // @[decode.scala 193:29 342:71]
  wire  _GEN_697 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h27 == outputBuffer_PRFDest |
    PRFValidList_39 : PRFValidList_39; // @[decode.scala 193:29 342:71]
  wire  _GEN_698 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h28 == outputBuffer_PRFDest |
    PRFValidList_40 : PRFValidList_40; // @[decode.scala 193:29 342:71]
  wire  _GEN_699 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h29 == outputBuffer_PRFDest |
    PRFValidList_41 : PRFValidList_41; // @[decode.scala 193:29 342:71]
  wire  _GEN_700 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h2a == outputBuffer_PRFDest |
    PRFValidList_42 : PRFValidList_42; // @[decode.scala 193:29 342:71]
  wire  _GEN_701 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h2b == outputBuffer_PRFDest |
    PRFValidList_43 : PRFValidList_43; // @[decode.scala 193:29 342:71]
  wire  _GEN_702 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h2c == outputBuffer_PRFDest |
    PRFValidList_44 : PRFValidList_44; // @[decode.scala 193:29 342:71]
  wire  _GEN_703 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h2d == outputBuffer_PRFDest |
    PRFValidList_45 : PRFValidList_45; // @[decode.scala 193:29 342:71]
  wire  _GEN_704 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h2e == outputBuffer_PRFDest |
    PRFValidList_46 : PRFValidList_46; // @[decode.scala 193:29 342:71]
  wire  _GEN_705 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h2f == outputBuffer_PRFDest |
    PRFValidList_47 : PRFValidList_47; // @[decode.scala 193:29 342:71]
  wire  _GEN_706 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h30 == outputBuffer_PRFDest |
    PRFValidList_48 : PRFValidList_48; // @[decode.scala 193:29 342:71]
  wire  _GEN_707 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h31 == outputBuffer_PRFDest |
    PRFValidList_49 : PRFValidList_49; // @[decode.scala 193:29 342:71]
  wire  _GEN_708 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h32 == outputBuffer_PRFDest |
    PRFValidList_50 : PRFValidList_50; // @[decode.scala 193:29 342:71]
  wire  _GEN_709 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h33 == outputBuffer_PRFDest |
    PRFValidList_51 : PRFValidList_51; // @[decode.scala 193:29 342:71]
  wire  _GEN_710 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h34 == outputBuffer_PRFDest |
    PRFValidList_52 : PRFValidList_52; // @[decode.scala 193:29 342:71]
  wire  _GEN_711 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h35 == outputBuffer_PRFDest |
    PRFValidList_53 : PRFValidList_53; // @[decode.scala 193:29 342:71]
  wire  _GEN_712 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h36 == outputBuffer_PRFDest |
    PRFValidList_54 : PRFValidList_54; // @[decode.scala 193:29 342:71]
  wire  _GEN_713 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h37 == outputBuffer_PRFDest |
    PRFValidList_55 : PRFValidList_55; // @[decode.scala 193:29 342:71]
  wire  _GEN_714 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h38 == outputBuffer_PRFDest |
    PRFValidList_56 : PRFValidList_56; // @[decode.scala 193:29 342:71]
  wire  _GEN_715 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h39 == outputBuffer_PRFDest |
    PRFValidList_57 : PRFValidList_57; // @[decode.scala 193:29 342:71]
  wire  _GEN_716 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h3a == outputBuffer_PRFDest |
    PRFValidList_58 : PRFValidList_58; // @[decode.scala 193:29 342:71]
  wire  _GEN_717 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h3b == outputBuffer_PRFDest |
    PRFValidList_59 : PRFValidList_59; // @[decode.scala 193:29 342:71]
  wire  _GEN_718 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h3c == outputBuffer_PRFDest |
    PRFValidList_60 : PRFValidList_60; // @[decode.scala 193:29 342:71]
  wire  _GEN_719 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h3d == outputBuffer_PRFDest |
    PRFValidList_61 : PRFValidList_61; // @[decode.scala 193:29 342:71]
  wire  _GEN_720 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h3e == outputBuffer_PRFDest |
    PRFValidList_62 : PRFValidList_62; // @[decode.scala 193:29 342:71]
  wire  _GEN_721 = jumpAddrWrite_fired & outputBuffer_instruction[11:7] != 5'h0 ? 6'h3f == outputBuffer_PRFDest |
    PRFValidList_63 : PRFValidList_63; // @[decode.scala 193:29 342:71]
  wire  _GEN_722 = 6'h0 == freeRegAddr ? 1'h0 : _GEN_530; // @[decode.scala 346:{33,33}]
  wire  _GEN_723 = 6'h1 == freeRegAddr ? 1'h0 : _GEN_531; // @[decode.scala 346:{33,33}]
  wire  _GEN_724 = 6'h2 == freeRegAddr ? 1'h0 : _GEN_532; // @[decode.scala 346:{33,33}]
  wire  _GEN_725 = 6'h3 == freeRegAddr ? 1'h0 : _GEN_533; // @[decode.scala 346:{33,33}]
  wire  _GEN_726 = 6'h4 == freeRegAddr ? 1'h0 : _GEN_534; // @[decode.scala 346:{33,33}]
  wire  _GEN_727 = 6'h5 == freeRegAddr ? 1'h0 : _GEN_535; // @[decode.scala 346:{33,33}]
  wire  _GEN_728 = 6'h6 == freeRegAddr ? 1'h0 : _GEN_536; // @[decode.scala 346:{33,33}]
  wire  _GEN_729 = 6'h7 == freeRegAddr ? 1'h0 : _GEN_537; // @[decode.scala 346:{33,33}]
  wire  _GEN_730 = 6'h8 == freeRegAddr ? 1'h0 : _GEN_538; // @[decode.scala 346:{33,33}]
  wire  _GEN_731 = 6'h9 == freeRegAddr ? 1'h0 : _GEN_539; // @[decode.scala 346:{33,33}]
  wire  _GEN_732 = 6'ha == freeRegAddr ? 1'h0 : _GEN_540; // @[decode.scala 346:{33,33}]
  wire  _GEN_733 = 6'hb == freeRegAddr ? 1'h0 : _GEN_541; // @[decode.scala 346:{33,33}]
  wire  _GEN_734 = 6'hc == freeRegAddr ? 1'h0 : _GEN_542; // @[decode.scala 346:{33,33}]
  wire  _GEN_735 = 6'hd == freeRegAddr ? 1'h0 : _GEN_543; // @[decode.scala 346:{33,33}]
  wire  _GEN_736 = 6'he == freeRegAddr ? 1'h0 : _GEN_544; // @[decode.scala 346:{33,33}]
  wire  _GEN_737 = 6'hf == freeRegAddr ? 1'h0 : _GEN_545; // @[decode.scala 346:{33,33}]
  wire  _GEN_738 = 6'h10 == freeRegAddr ? 1'h0 : _GEN_546; // @[decode.scala 346:{33,33}]
  wire  _GEN_739 = 6'h11 == freeRegAddr ? 1'h0 : _GEN_547; // @[decode.scala 346:{33,33}]
  wire  _GEN_740 = 6'h12 == freeRegAddr ? 1'h0 : _GEN_548; // @[decode.scala 346:{33,33}]
  wire  _GEN_741 = 6'h13 == freeRegAddr ? 1'h0 : _GEN_549; // @[decode.scala 346:{33,33}]
  wire  _GEN_742 = 6'h14 == freeRegAddr ? 1'h0 : _GEN_550; // @[decode.scala 346:{33,33}]
  wire  _GEN_743 = 6'h15 == freeRegAddr ? 1'h0 : _GEN_551; // @[decode.scala 346:{33,33}]
  wire  _GEN_744 = 6'h16 == freeRegAddr ? 1'h0 : _GEN_552; // @[decode.scala 346:{33,33}]
  wire  _GEN_745 = 6'h17 == freeRegAddr ? 1'h0 : _GEN_553; // @[decode.scala 346:{33,33}]
  wire  _GEN_746 = 6'h18 == freeRegAddr ? 1'h0 : _GEN_554; // @[decode.scala 346:{33,33}]
  wire  _GEN_747 = 6'h19 == freeRegAddr ? 1'h0 : _GEN_555; // @[decode.scala 346:{33,33}]
  wire  _GEN_748 = 6'h1a == freeRegAddr ? 1'h0 : _GEN_556; // @[decode.scala 346:{33,33}]
  wire  _GEN_749 = 6'h1b == freeRegAddr ? 1'h0 : _GEN_557; // @[decode.scala 346:{33,33}]
  wire  _GEN_750 = 6'h1c == freeRegAddr ? 1'h0 : _GEN_558; // @[decode.scala 346:{33,33}]
  wire  _GEN_751 = 6'h1d == freeRegAddr ? 1'h0 : _GEN_559; // @[decode.scala 346:{33,33}]
  wire  _GEN_752 = 6'h1e == freeRegAddr ? 1'h0 : _GEN_560; // @[decode.scala 346:{33,33}]
  wire  _GEN_753 = 6'h1f == freeRegAddr ? 1'h0 : _GEN_561; // @[decode.scala 346:{33,33}]
  wire  _GEN_754 = 6'h20 == freeRegAddr ? 1'h0 : _GEN_562; // @[decode.scala 346:{33,33}]
  wire  _GEN_755 = 6'h21 == freeRegAddr ? 1'h0 : _GEN_563; // @[decode.scala 346:{33,33}]
  wire  _GEN_756 = 6'h22 == freeRegAddr ? 1'h0 : _GEN_564; // @[decode.scala 346:{33,33}]
  wire  _GEN_757 = 6'h23 == freeRegAddr ? 1'h0 : _GEN_565; // @[decode.scala 346:{33,33}]
  wire  _GEN_758 = 6'h24 == freeRegAddr ? 1'h0 : _GEN_566; // @[decode.scala 346:{33,33}]
  wire  _GEN_759 = 6'h25 == freeRegAddr ? 1'h0 : _GEN_567; // @[decode.scala 346:{33,33}]
  wire  _GEN_760 = 6'h26 == freeRegAddr ? 1'h0 : _GEN_568; // @[decode.scala 346:{33,33}]
  wire  _GEN_761 = 6'h27 == freeRegAddr ? 1'h0 : _GEN_569; // @[decode.scala 346:{33,33}]
  wire  _GEN_762 = 6'h28 == freeRegAddr ? 1'h0 : _GEN_570; // @[decode.scala 346:{33,33}]
  wire  _GEN_763 = 6'h29 == freeRegAddr ? 1'h0 : _GEN_571; // @[decode.scala 346:{33,33}]
  wire  _GEN_764 = 6'h2a == freeRegAddr ? 1'h0 : _GEN_572; // @[decode.scala 346:{33,33}]
  wire  _GEN_765 = 6'h2b == freeRegAddr ? 1'h0 : _GEN_573; // @[decode.scala 346:{33,33}]
  wire  _GEN_766 = 6'h2c == freeRegAddr ? 1'h0 : _GEN_574; // @[decode.scala 346:{33,33}]
  wire  _GEN_767 = 6'h2d == freeRegAddr ? 1'h0 : _GEN_575; // @[decode.scala 346:{33,33}]
  wire  _GEN_768 = 6'h2e == freeRegAddr ? 1'h0 : _GEN_576; // @[decode.scala 346:{33,33}]
  wire  _GEN_769 = 6'h2f == freeRegAddr ? 1'h0 : _GEN_577; // @[decode.scala 346:{33,33}]
  wire  _GEN_770 = 6'h30 == freeRegAddr ? 1'h0 : _GEN_578; // @[decode.scala 346:{33,33}]
  wire  _GEN_771 = 6'h31 == freeRegAddr ? 1'h0 : _GEN_579; // @[decode.scala 346:{33,33}]
  wire  _GEN_772 = 6'h32 == freeRegAddr ? 1'h0 : _GEN_580; // @[decode.scala 346:{33,33}]
  wire  _GEN_773 = 6'h33 == freeRegAddr ? 1'h0 : _GEN_581; // @[decode.scala 346:{33,33}]
  wire  _GEN_774 = 6'h34 == freeRegAddr ? 1'h0 : _GEN_582; // @[decode.scala 346:{33,33}]
  wire  _GEN_775 = 6'h35 == freeRegAddr ? 1'h0 : _GEN_583; // @[decode.scala 346:{33,33}]
  wire  _GEN_776 = 6'h36 == freeRegAddr ? 1'h0 : _GEN_584; // @[decode.scala 346:{33,33}]
  wire  _GEN_777 = 6'h37 == freeRegAddr ? 1'h0 : _GEN_585; // @[decode.scala 346:{33,33}]
  wire  _GEN_778 = 6'h38 == freeRegAddr ? 1'h0 : _GEN_586; // @[decode.scala 346:{33,33}]
  wire  _GEN_779 = 6'h39 == freeRegAddr ? 1'h0 : _GEN_587; // @[decode.scala 346:{33,33}]
  wire  _GEN_780 = 6'h3a == freeRegAddr ? 1'h0 : _GEN_588; // @[decode.scala 346:{33,33}]
  wire  _GEN_781 = 6'h3b == freeRegAddr ? 1'h0 : _GEN_589; // @[decode.scala 346:{33,33}]
  wire  _GEN_782 = 6'h3c == freeRegAddr ? 1'h0 : _GEN_590; // @[decode.scala 346:{33,33}]
  wire  _GEN_783 = 6'h3d == freeRegAddr ? 1'h0 : _GEN_591; // @[decode.scala 346:{33,33}]
  wire  _GEN_784 = 6'h3e == freeRegAddr ? 1'h0 : _GEN_592; // @[decode.scala 346:{33,33}]
  wire  _GEN_786 = 6'h0 == freeRegAddr ? 1'h0 : _GEN_658; // @[decode.scala 347:{33,33}]
  wire  _GEN_787 = 6'h1 == freeRegAddr ? 1'h0 : _GEN_659; // @[decode.scala 347:{33,33}]
  wire  _GEN_788 = 6'h2 == freeRegAddr ? 1'h0 : _GEN_660; // @[decode.scala 347:{33,33}]
  wire  _GEN_789 = 6'h3 == freeRegAddr ? 1'h0 : _GEN_661; // @[decode.scala 347:{33,33}]
  wire  _GEN_790 = 6'h4 == freeRegAddr ? 1'h0 : _GEN_662; // @[decode.scala 347:{33,33}]
  wire  _GEN_791 = 6'h5 == freeRegAddr ? 1'h0 : _GEN_663; // @[decode.scala 347:{33,33}]
  wire  _GEN_792 = 6'h6 == freeRegAddr ? 1'h0 : _GEN_664; // @[decode.scala 347:{33,33}]
  wire  _GEN_793 = 6'h7 == freeRegAddr ? 1'h0 : _GEN_665; // @[decode.scala 347:{33,33}]
  wire  _GEN_794 = 6'h8 == freeRegAddr ? 1'h0 : _GEN_666; // @[decode.scala 347:{33,33}]
  wire  _GEN_795 = 6'h9 == freeRegAddr ? 1'h0 : _GEN_667; // @[decode.scala 347:{33,33}]
  wire  _GEN_796 = 6'ha == freeRegAddr ? 1'h0 : _GEN_668; // @[decode.scala 347:{33,33}]
  wire  _GEN_797 = 6'hb == freeRegAddr ? 1'h0 : _GEN_669; // @[decode.scala 347:{33,33}]
  wire  _GEN_798 = 6'hc == freeRegAddr ? 1'h0 : _GEN_670; // @[decode.scala 347:{33,33}]
  wire  _GEN_799 = 6'hd == freeRegAddr ? 1'h0 : _GEN_671; // @[decode.scala 347:{33,33}]
  wire  _GEN_800 = 6'he == freeRegAddr ? 1'h0 : _GEN_672; // @[decode.scala 347:{33,33}]
  wire  _GEN_801 = 6'hf == freeRegAddr ? 1'h0 : _GEN_673; // @[decode.scala 347:{33,33}]
  wire  _GEN_802 = 6'h10 == freeRegAddr ? 1'h0 : _GEN_674; // @[decode.scala 347:{33,33}]
  wire  _GEN_803 = 6'h11 == freeRegAddr ? 1'h0 : _GEN_675; // @[decode.scala 347:{33,33}]
  wire  _GEN_804 = 6'h12 == freeRegAddr ? 1'h0 : _GEN_676; // @[decode.scala 347:{33,33}]
  wire  _GEN_805 = 6'h13 == freeRegAddr ? 1'h0 : _GEN_677; // @[decode.scala 347:{33,33}]
  wire  _GEN_806 = 6'h14 == freeRegAddr ? 1'h0 : _GEN_678; // @[decode.scala 347:{33,33}]
  wire  _GEN_807 = 6'h15 == freeRegAddr ? 1'h0 : _GEN_679; // @[decode.scala 347:{33,33}]
  wire  _GEN_808 = 6'h16 == freeRegAddr ? 1'h0 : _GEN_680; // @[decode.scala 347:{33,33}]
  wire  _GEN_809 = 6'h17 == freeRegAddr ? 1'h0 : _GEN_681; // @[decode.scala 347:{33,33}]
  wire  _GEN_810 = 6'h18 == freeRegAddr ? 1'h0 : _GEN_682; // @[decode.scala 347:{33,33}]
  wire  _GEN_811 = 6'h19 == freeRegAddr ? 1'h0 : _GEN_683; // @[decode.scala 347:{33,33}]
  wire  _GEN_812 = 6'h1a == freeRegAddr ? 1'h0 : _GEN_684; // @[decode.scala 347:{33,33}]
  wire  _GEN_813 = 6'h1b == freeRegAddr ? 1'h0 : _GEN_685; // @[decode.scala 347:{33,33}]
  wire  _GEN_814 = 6'h1c == freeRegAddr ? 1'h0 : _GEN_686; // @[decode.scala 347:{33,33}]
  wire  _GEN_815 = 6'h1d == freeRegAddr ? 1'h0 : _GEN_687; // @[decode.scala 347:{33,33}]
  wire  _GEN_816 = 6'h1e == freeRegAddr ? 1'h0 : _GEN_688; // @[decode.scala 347:{33,33}]
  wire  _GEN_817 = 6'h1f == freeRegAddr ? 1'h0 : _GEN_689; // @[decode.scala 347:{33,33}]
  wire  _GEN_818 = 6'h20 == freeRegAddr ? 1'h0 : _GEN_690; // @[decode.scala 347:{33,33}]
  wire  _GEN_819 = 6'h21 == freeRegAddr ? 1'h0 : _GEN_691; // @[decode.scala 347:{33,33}]
  wire  _GEN_820 = 6'h22 == freeRegAddr ? 1'h0 : _GEN_692; // @[decode.scala 347:{33,33}]
  wire  _GEN_821 = 6'h23 == freeRegAddr ? 1'h0 : _GEN_693; // @[decode.scala 347:{33,33}]
  wire  _GEN_822 = 6'h24 == freeRegAddr ? 1'h0 : _GEN_694; // @[decode.scala 347:{33,33}]
  wire  _GEN_823 = 6'h25 == freeRegAddr ? 1'h0 : _GEN_695; // @[decode.scala 347:{33,33}]
  wire  _GEN_824 = 6'h26 == freeRegAddr ? 1'h0 : _GEN_696; // @[decode.scala 347:{33,33}]
  wire  _GEN_825 = 6'h27 == freeRegAddr ? 1'h0 : _GEN_697; // @[decode.scala 347:{33,33}]
  wire  _GEN_826 = 6'h28 == freeRegAddr ? 1'h0 : _GEN_698; // @[decode.scala 347:{33,33}]
  wire  _GEN_827 = 6'h29 == freeRegAddr ? 1'h0 : _GEN_699; // @[decode.scala 347:{33,33}]
  wire  _GEN_828 = 6'h2a == freeRegAddr ? 1'h0 : _GEN_700; // @[decode.scala 347:{33,33}]
  wire  _GEN_829 = 6'h2b == freeRegAddr ? 1'h0 : _GEN_701; // @[decode.scala 347:{33,33}]
  wire  _GEN_830 = 6'h2c == freeRegAddr ? 1'h0 : _GEN_702; // @[decode.scala 347:{33,33}]
  wire  _GEN_831 = 6'h2d == freeRegAddr ? 1'h0 : _GEN_703; // @[decode.scala 347:{33,33}]
  wire  _GEN_832 = 6'h2e == freeRegAddr ? 1'h0 : _GEN_704; // @[decode.scala 347:{33,33}]
  wire  _GEN_833 = 6'h2f == freeRegAddr ? 1'h0 : _GEN_705; // @[decode.scala 347:{33,33}]
  wire  _GEN_834 = 6'h30 == freeRegAddr ? 1'h0 : _GEN_706; // @[decode.scala 347:{33,33}]
  wire  _GEN_835 = 6'h31 == freeRegAddr ? 1'h0 : _GEN_707; // @[decode.scala 347:{33,33}]
  wire  _GEN_836 = 6'h32 == freeRegAddr ? 1'h0 : _GEN_708; // @[decode.scala 347:{33,33}]
  wire  _GEN_837 = 6'h33 == freeRegAddr ? 1'h0 : _GEN_709; // @[decode.scala 347:{33,33}]
  wire  _GEN_838 = 6'h34 == freeRegAddr ? 1'h0 : _GEN_710; // @[decode.scala 347:{33,33}]
  wire  _GEN_839 = 6'h35 == freeRegAddr ? 1'h0 : _GEN_711; // @[decode.scala 347:{33,33}]
  wire  _GEN_840 = 6'h36 == freeRegAddr ? 1'h0 : _GEN_712; // @[decode.scala 347:{33,33}]
  wire  _GEN_841 = 6'h37 == freeRegAddr ? 1'h0 : _GEN_713; // @[decode.scala 347:{33,33}]
  wire  _GEN_842 = 6'h38 == freeRegAddr ? 1'h0 : _GEN_714; // @[decode.scala 347:{33,33}]
  wire  _GEN_843 = 6'h39 == freeRegAddr ? 1'h0 : _GEN_715; // @[decode.scala 347:{33,33}]
  wire  _GEN_844 = 6'h3a == freeRegAddr ? 1'h0 : _GEN_716; // @[decode.scala 347:{33,33}]
  wire  _GEN_845 = 6'h3b == freeRegAddr ? 1'h0 : _GEN_717; // @[decode.scala 347:{33,33}]
  wire  _GEN_846 = 6'h3c == freeRegAddr ? 1'h0 : _GEN_718; // @[decode.scala 347:{33,33}]
  wire  _GEN_847 = 6'h3d == freeRegAddr ? 1'h0 : _GEN_719; // @[decode.scala 347:{33,33}]
  wire  _GEN_848 = 6'h3e == freeRegAddr ? 1'h0 : _GEN_720; // @[decode.scala 347:{33,33}]
  wire  _GEN_849 = 6'h3f == freeRegAddr ? 1'h0 : _GEN_721; // @[decode.scala 347:{33,33}]
  wire [5:0] _GEN_850 = 5'h0 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_0; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_851 = 5'h1 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_1; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_852 = 5'h2 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_2; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_853 = 5'h3 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_3; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_854 = 5'h4 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_4; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_855 = 5'h5 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_5; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_856 = 5'h6 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_6; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_857 = 5'h7 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_7; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_858 = 5'h8 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_8; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_859 = 5'h9 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_9; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_860 = 5'ha == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_10; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_861 = 5'hb == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_11; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_862 = 5'hc == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_12; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_863 = 5'hd == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_13; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_864 = 5'he == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_14; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_865 = 5'hf == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_15; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_866 = 5'h10 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_16; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_867 = 5'h11 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_17; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_868 = 5'h12 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_18; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_869 = 5'h13 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_19; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_870 = 5'h14 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_20; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_871 = 5'h15 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_21; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_872 = 5'h16 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_22; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_873 = 5'h17 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_23; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_874 = 5'h18 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_24; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_875 = 5'h19 == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_25; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_876 = 5'h1a == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_26; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_877 = 5'h1b == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_27; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_878 = 5'h1c == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_28; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_879 = 5'h1d == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_29; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_880 = 5'h1e == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_30; // @[decode.scala 348:{33,33} 301:36]
  wire [5:0] _GEN_881 = 5'h1f == inputBuffer_instruction[11:7] ? freeRegAddr : frontEndRegMap_31; // @[decode.scala 348:{33,33} 301:36]
  wire  _GEN_882 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_722 : _GEN_530; // @[decode.scala 345:55]
  wire  _GEN_883 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_723 : _GEN_531; // @[decode.scala 345:55]
  wire  _GEN_884 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_724 : _GEN_532; // @[decode.scala 345:55]
  wire  _GEN_885 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_725 : _GEN_533; // @[decode.scala 345:55]
  wire  _GEN_886 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_726 : _GEN_534; // @[decode.scala 345:55]
  wire  _GEN_887 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_727 : _GEN_535; // @[decode.scala 345:55]
  wire  _GEN_888 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_728 : _GEN_536; // @[decode.scala 345:55]
  wire  _GEN_889 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_729 : _GEN_537; // @[decode.scala 345:55]
  wire  _GEN_890 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_730 : _GEN_538; // @[decode.scala 345:55]
  wire  _GEN_891 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_731 : _GEN_539; // @[decode.scala 345:55]
  wire  _GEN_892 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_732 : _GEN_540; // @[decode.scala 345:55]
  wire  _GEN_893 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_733 : _GEN_541; // @[decode.scala 345:55]
  wire  _GEN_894 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_734 : _GEN_542; // @[decode.scala 345:55]
  wire  _GEN_895 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_735 : _GEN_543; // @[decode.scala 345:55]
  wire  _GEN_896 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_736 : _GEN_544; // @[decode.scala 345:55]
  wire  _GEN_897 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_737 : _GEN_545; // @[decode.scala 345:55]
  wire  _GEN_898 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_738 : _GEN_546; // @[decode.scala 345:55]
  wire  _GEN_899 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_739 : _GEN_547; // @[decode.scala 345:55]
  wire  _GEN_900 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_740 : _GEN_548; // @[decode.scala 345:55]
  wire  _GEN_901 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_741 : _GEN_549; // @[decode.scala 345:55]
  wire  _GEN_902 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_742 : _GEN_550; // @[decode.scala 345:55]
  wire  _GEN_903 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_743 : _GEN_551; // @[decode.scala 345:55]
  wire  _GEN_904 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_744 : _GEN_552; // @[decode.scala 345:55]
  wire  _GEN_905 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_745 : _GEN_553; // @[decode.scala 345:55]
  wire  _GEN_906 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_746 : _GEN_554; // @[decode.scala 345:55]
  wire  _GEN_907 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_747 : _GEN_555; // @[decode.scala 345:55]
  wire  _GEN_908 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_748 : _GEN_556; // @[decode.scala 345:55]
  wire  _GEN_909 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_749 : _GEN_557; // @[decode.scala 345:55]
  wire  _GEN_910 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_750 : _GEN_558; // @[decode.scala 345:55]
  wire  _GEN_911 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_751 : _GEN_559; // @[decode.scala 345:55]
  wire  _GEN_912 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_752 : _GEN_560; // @[decode.scala 345:55]
  wire  _GEN_913 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_753 : _GEN_561; // @[decode.scala 345:55]
  wire  _GEN_914 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_754 : _GEN_562; // @[decode.scala 345:55]
  wire  _GEN_915 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_755 : _GEN_563; // @[decode.scala 345:55]
  wire  _GEN_916 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_756 : _GEN_564; // @[decode.scala 345:55]
  wire  _GEN_917 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_757 : _GEN_565; // @[decode.scala 345:55]
  wire  _GEN_918 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_758 : _GEN_566; // @[decode.scala 345:55]
  wire  _GEN_919 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_759 : _GEN_567; // @[decode.scala 345:55]
  wire  _GEN_920 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_760 : _GEN_568; // @[decode.scala 345:55]
  wire  _GEN_921 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_761 : _GEN_569; // @[decode.scala 345:55]
  wire  _GEN_922 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_762 : _GEN_570; // @[decode.scala 345:55]
  wire  _GEN_923 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_763 : _GEN_571; // @[decode.scala 345:55]
  wire  _GEN_924 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_764 : _GEN_572; // @[decode.scala 345:55]
  wire  _GEN_925 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_765 : _GEN_573; // @[decode.scala 345:55]
  wire  _GEN_926 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_766 : _GEN_574; // @[decode.scala 345:55]
  wire  _GEN_927 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_767 : _GEN_575; // @[decode.scala 345:55]
  wire  _GEN_928 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_768 : _GEN_576; // @[decode.scala 345:55]
  wire  _GEN_929 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_769 : _GEN_577; // @[decode.scala 345:55]
  wire  _GEN_930 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_770 : _GEN_578; // @[decode.scala 345:55]
  wire  _GEN_931 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_771 : _GEN_579; // @[decode.scala 345:55]
  wire  _GEN_932 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_772 : _GEN_580; // @[decode.scala 345:55]
  wire  _GEN_933 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_773 : _GEN_581; // @[decode.scala 345:55]
  wire  _GEN_934 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_774 : _GEN_582; // @[decode.scala 345:55]
  wire  _GEN_935 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_775 : _GEN_583; // @[decode.scala 345:55]
  wire  _GEN_936 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_776 : _GEN_584; // @[decode.scala 345:55]
  wire  _GEN_937 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_777 : _GEN_585; // @[decode.scala 345:55]
  wire  _GEN_938 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_778 : _GEN_586; // @[decode.scala 345:55]
  wire  _GEN_939 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_779 : _GEN_587; // @[decode.scala 345:55]
  wire  _GEN_940 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_780 : _GEN_588; // @[decode.scala 345:55]
  wire  _GEN_941 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_781 : _GEN_589; // @[decode.scala 345:55]
  wire  _GEN_942 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_782 : _GEN_590; // @[decode.scala 345:55]
  wire  _GEN_943 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_783 : _GEN_591; // @[decode.scala 345:55]
  wire  _GEN_944 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_784 : _GEN_592; // @[decode.scala 345:55]
  wire  _GEN_946 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_786 : _GEN_658; // @[decode.scala 345:55]
  wire  _GEN_947 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_787 : _GEN_659; // @[decode.scala 345:55]
  wire  _GEN_948 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_788 : _GEN_660; // @[decode.scala 345:55]
  wire  _GEN_949 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_789 : _GEN_661; // @[decode.scala 345:55]
  wire  _GEN_950 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_790 : _GEN_662; // @[decode.scala 345:55]
  wire  _GEN_951 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_791 : _GEN_663; // @[decode.scala 345:55]
  wire  _GEN_952 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_792 : _GEN_664; // @[decode.scala 345:55]
  wire  _GEN_953 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_793 : _GEN_665; // @[decode.scala 345:55]
  wire  _GEN_954 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_794 : _GEN_666; // @[decode.scala 345:55]
  wire  _GEN_955 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_795 : _GEN_667; // @[decode.scala 345:55]
  wire  _GEN_956 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_796 : _GEN_668; // @[decode.scala 345:55]
  wire  _GEN_957 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_797 : _GEN_669; // @[decode.scala 345:55]
  wire  _GEN_958 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_798 : _GEN_670; // @[decode.scala 345:55]
  wire  _GEN_959 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_799 : _GEN_671; // @[decode.scala 345:55]
  wire  _GEN_960 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_800 : _GEN_672; // @[decode.scala 345:55]
  wire  _GEN_961 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_801 : _GEN_673; // @[decode.scala 345:55]
  wire  _GEN_962 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_802 : _GEN_674; // @[decode.scala 345:55]
  wire  _GEN_963 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_803 : _GEN_675; // @[decode.scala 345:55]
  wire  _GEN_964 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_804 : _GEN_676; // @[decode.scala 345:55]
  wire  _GEN_965 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_805 : _GEN_677; // @[decode.scala 345:55]
  wire  _GEN_966 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_806 : _GEN_678; // @[decode.scala 345:55]
  wire  _GEN_967 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_807 : _GEN_679; // @[decode.scala 345:55]
  wire  _GEN_968 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_808 : _GEN_680; // @[decode.scala 345:55]
  wire  _GEN_969 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_809 : _GEN_681; // @[decode.scala 345:55]
  wire  _GEN_970 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_810 : _GEN_682; // @[decode.scala 345:55]
  wire  _GEN_971 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_811 : _GEN_683; // @[decode.scala 345:55]
  wire  _GEN_972 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_812 : _GEN_684; // @[decode.scala 345:55]
  wire  _GEN_973 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_813 : _GEN_685; // @[decode.scala 345:55]
  wire  _GEN_974 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_814 : _GEN_686; // @[decode.scala 345:55]
  wire  _GEN_975 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_815 : _GEN_687; // @[decode.scala 345:55]
  wire  _GEN_976 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_816 : _GEN_688; // @[decode.scala 345:55]
  wire  _GEN_977 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_817 : _GEN_689; // @[decode.scala 345:55]
  wire  _GEN_978 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_818 : _GEN_690; // @[decode.scala 345:55]
  wire  _GEN_979 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_819 : _GEN_691; // @[decode.scala 345:55]
  wire  _GEN_980 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_820 : _GEN_692; // @[decode.scala 345:55]
  wire  _GEN_981 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_821 : _GEN_693; // @[decode.scala 345:55]
  wire  _GEN_982 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_822 : _GEN_694; // @[decode.scala 345:55]
  wire  _GEN_983 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_823 : _GEN_695; // @[decode.scala 345:55]
  wire  _GEN_984 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_824 : _GEN_696; // @[decode.scala 345:55]
  wire  _GEN_985 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_825 : _GEN_697; // @[decode.scala 345:55]
  wire  _GEN_986 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_826 : _GEN_698; // @[decode.scala 345:55]
  wire  _GEN_987 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_827 : _GEN_699; // @[decode.scala 345:55]
  wire  _GEN_988 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_828 : _GEN_700; // @[decode.scala 345:55]
  wire  _GEN_989 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_829 : _GEN_701; // @[decode.scala 345:55]
  wire  _GEN_990 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_830 : _GEN_702; // @[decode.scala 345:55]
  wire  _GEN_991 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_831 : _GEN_703; // @[decode.scala 345:55]
  wire  _GEN_992 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_832 : _GEN_704; // @[decode.scala 345:55]
  wire  _GEN_993 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_833 : _GEN_705; // @[decode.scala 345:55]
  wire  _GEN_994 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_834 : _GEN_706; // @[decode.scala 345:55]
  wire  _GEN_995 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_835 : _GEN_707; // @[decode.scala 345:55]
  wire  _GEN_996 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_836 : _GEN_708; // @[decode.scala 345:55]
  wire  _GEN_997 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_837 : _GEN_709; // @[decode.scala 345:55]
  wire  _GEN_998 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_838 : _GEN_710; // @[decode.scala 345:55]
  wire  _GEN_999 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_839 : _GEN_711; // @[decode.scala 345:55]
  wire  _GEN_1000 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_840 : _GEN_712; // @[decode.scala 345:55]
  wire  _GEN_1001 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_841 : _GEN_713; // @[decode.scala 345:55]
  wire  _GEN_1002 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_842 : _GEN_714; // @[decode.scala 345:55]
  wire  _GEN_1003 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_843 : _GEN_715; // @[decode.scala 345:55]
  wire  _GEN_1004 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_844 : _GEN_716; // @[decode.scala 345:55]
  wire  _GEN_1005 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_845 : _GEN_717; // @[decode.scala 345:55]
  wire  _GEN_1006 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_846 : _GEN_718; // @[decode.scala 345:55]
  wire  _GEN_1007 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_847 : _GEN_719; // @[decode.scala 345:55]
  wire  _GEN_1008 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_848 : _GEN_720; // @[decode.scala 345:55]
  wire  _GEN_1009 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_849 : _GEN_721; // @[decode.scala 345:55]
  wire [5:0] _GEN_1010 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_850 : frontEndRegMap_0; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1011 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_851 : frontEndRegMap_1; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1012 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_852 : frontEndRegMap_2; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1013 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_853 : frontEndRegMap_3; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1014 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_854 : frontEndRegMap_4; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1015 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_855 : frontEndRegMap_5; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1016 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_856 : frontEndRegMap_6; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1017 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_857 : frontEndRegMap_7; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1018 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_858 : frontEndRegMap_8; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1019 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_859 : frontEndRegMap_9; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1020 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_860 : frontEndRegMap_10; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1021 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_861 : frontEndRegMap_11; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1022 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_862 : frontEndRegMap_12; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1023 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_863 : frontEndRegMap_13; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1024 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_864 : frontEndRegMap_14; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1025 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_865 : frontEndRegMap_15; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1026 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_866 : frontEndRegMap_16; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1027 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_867 : frontEndRegMap_17; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1028 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_868 : frontEndRegMap_18; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1029 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_869 : frontEndRegMap_19; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1030 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_870 : frontEndRegMap_20; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1031 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_871 : frontEndRegMap_21; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1032 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_872 : frontEndRegMap_22; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1033 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_873 : frontEndRegMap_23; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1034 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_874 : frontEndRegMap_24; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1035 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_875 : frontEndRegMap_25; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1036 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_876 : frontEndRegMap_26; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1037 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_877 : frontEndRegMap_27; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1038 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_878 : frontEndRegMap_28; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1039 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_879 : frontEndRegMap_29; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1040 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_880 : frontEndRegMap_30; // @[decode.scala 301:36 345:55]
  wire [5:0] _GEN_1041 = ~branchEvalIn_fired | branchEvalIn_passFail ? _GEN_881 : frontEndRegMap_31; // @[decode.scala 301:36 345:55]
  wire  _GEN_1042 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_882 : _GEN_530; // @[decode.scala 344:149]
  wire  _GEN_1043 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_883 : _GEN_531; // @[decode.scala 344:149]
  wire  _GEN_1044 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_884 : _GEN_532; // @[decode.scala 344:149]
  wire  _GEN_1045 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_885 : _GEN_533; // @[decode.scala 344:149]
  wire  _GEN_1046 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_886 : _GEN_534; // @[decode.scala 344:149]
  wire  _GEN_1047 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_887 : _GEN_535; // @[decode.scala 344:149]
  wire  _GEN_1048 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_888 : _GEN_536; // @[decode.scala 344:149]
  wire  _GEN_1049 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_889 : _GEN_537; // @[decode.scala 344:149]
  wire  _GEN_1050 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_890 : _GEN_538; // @[decode.scala 344:149]
  wire  _GEN_1051 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_891 : _GEN_539; // @[decode.scala 344:149]
  wire  _GEN_1052 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_892 : _GEN_540; // @[decode.scala 344:149]
  wire  _GEN_1053 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_893 : _GEN_541; // @[decode.scala 344:149]
  wire  _GEN_1054 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_894 : _GEN_542; // @[decode.scala 344:149]
  wire  _GEN_1055 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_895 : _GEN_543; // @[decode.scala 344:149]
  wire  _GEN_1056 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_896 : _GEN_544; // @[decode.scala 344:149]
  wire  _GEN_1057 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_897 : _GEN_545; // @[decode.scala 344:149]
  wire  _GEN_1058 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_898 : _GEN_546; // @[decode.scala 344:149]
  wire  _GEN_1059 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_899 : _GEN_547; // @[decode.scala 344:149]
  wire  _GEN_1060 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_900 : _GEN_548; // @[decode.scala 344:149]
  wire  _GEN_1061 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_901 : _GEN_549; // @[decode.scala 344:149]
  wire  _GEN_1062 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_902 : _GEN_550; // @[decode.scala 344:149]
  wire  _GEN_1063 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_903 : _GEN_551; // @[decode.scala 344:149]
  wire  _GEN_1064 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_904 : _GEN_552; // @[decode.scala 344:149]
  wire  _GEN_1065 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_905 : _GEN_553; // @[decode.scala 344:149]
  wire  _GEN_1066 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_906 : _GEN_554; // @[decode.scala 344:149]
  wire  _GEN_1067 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_907 : _GEN_555; // @[decode.scala 344:149]
  wire  _GEN_1068 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_908 : _GEN_556; // @[decode.scala 344:149]
  wire  _GEN_1069 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_909 : _GEN_557; // @[decode.scala 344:149]
  wire  _GEN_1070 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_910 : _GEN_558; // @[decode.scala 344:149]
  wire  _GEN_1071 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_911 : _GEN_559; // @[decode.scala 344:149]
  wire  _GEN_1072 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_912 : _GEN_560; // @[decode.scala 344:149]
  wire  _GEN_1073 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_913 : _GEN_561; // @[decode.scala 344:149]
  wire  _GEN_1074 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_914 : _GEN_562; // @[decode.scala 344:149]
  wire  _GEN_1075 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_915 : _GEN_563; // @[decode.scala 344:149]
  wire  _GEN_1076 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_916 : _GEN_564; // @[decode.scala 344:149]
  wire  _GEN_1077 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_917 : _GEN_565; // @[decode.scala 344:149]
  wire  _GEN_1078 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_918 : _GEN_566; // @[decode.scala 344:149]
  wire  _GEN_1079 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_919 : _GEN_567; // @[decode.scala 344:149]
  wire  _GEN_1080 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_920 : _GEN_568; // @[decode.scala 344:149]
  wire  _GEN_1081 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_921 : _GEN_569; // @[decode.scala 344:149]
  wire  _GEN_1082 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_922 : _GEN_570; // @[decode.scala 344:149]
  wire  _GEN_1083 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_923 : _GEN_571; // @[decode.scala 344:149]
  wire  _GEN_1084 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_924 : _GEN_572; // @[decode.scala 344:149]
  wire  _GEN_1085 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_925 : _GEN_573; // @[decode.scala 344:149]
  wire  _GEN_1086 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_926 : _GEN_574; // @[decode.scala 344:149]
  wire  _GEN_1087 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_927 : _GEN_575; // @[decode.scala 344:149]
  wire  _GEN_1088 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_928 : _GEN_576; // @[decode.scala 344:149]
  wire  _GEN_1089 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_929 : _GEN_577; // @[decode.scala 344:149]
  wire  _GEN_1090 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_930 : _GEN_578; // @[decode.scala 344:149]
  wire  _GEN_1091 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_931 : _GEN_579; // @[decode.scala 344:149]
  wire  _GEN_1092 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_932 : _GEN_580; // @[decode.scala 344:149]
  wire  _GEN_1093 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_933 : _GEN_581; // @[decode.scala 344:149]
  wire  _GEN_1094 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_934 : _GEN_582; // @[decode.scala 344:149]
  wire  _GEN_1095 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_935 : _GEN_583; // @[decode.scala 344:149]
  wire  _GEN_1096 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_936 : _GEN_584; // @[decode.scala 344:149]
  wire  _GEN_1097 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_937 : _GEN_585; // @[decode.scala 344:149]
  wire  _GEN_1098 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_938 : _GEN_586; // @[decode.scala 344:149]
  wire  _GEN_1099 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_939 : _GEN_587; // @[decode.scala 344:149]
  wire  _GEN_1100 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_940 : _GEN_588; // @[decode.scala 344:149]
  wire  _GEN_1101 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_941 : _GEN_589; // @[decode.scala 344:149]
  wire  _GEN_1102 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_942 : _GEN_590; // @[decode.scala 344:149]
  wire  _GEN_1103 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_943 : _GEN_591; // @[decode.scala 344:149]
  wire  _GEN_1104 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_944 : _GEN_592; // @[decode.scala 344:149]
  wire  _GEN_1106 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_946 : _GEN_658; // @[decode.scala 344:149]
  wire  _GEN_1107 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_947 : _GEN_659; // @[decode.scala 344:149]
  wire  _GEN_1108 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_948 : _GEN_660; // @[decode.scala 344:149]
  wire  _GEN_1109 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_949 : _GEN_661; // @[decode.scala 344:149]
  wire  _GEN_1110 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_950 : _GEN_662; // @[decode.scala 344:149]
  wire  _GEN_1111 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_951 : _GEN_663; // @[decode.scala 344:149]
  wire  _GEN_1112 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_952 : _GEN_664; // @[decode.scala 344:149]
  wire  _GEN_1113 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_953 : _GEN_665; // @[decode.scala 344:149]
  wire  _GEN_1114 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_954 : _GEN_666; // @[decode.scala 344:149]
  wire  _GEN_1115 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_955 : _GEN_667; // @[decode.scala 344:149]
  wire  _GEN_1116 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_956 : _GEN_668; // @[decode.scala 344:149]
  wire  _GEN_1117 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_957 : _GEN_669; // @[decode.scala 344:149]
  wire  _GEN_1118 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_958 : _GEN_670; // @[decode.scala 344:149]
  wire  _GEN_1119 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_959 : _GEN_671; // @[decode.scala 344:149]
  wire  _GEN_1120 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_960 : _GEN_672; // @[decode.scala 344:149]
  wire  _GEN_1121 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_961 : _GEN_673; // @[decode.scala 344:149]
  wire  _GEN_1122 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_962 : _GEN_674; // @[decode.scala 344:149]
  wire  _GEN_1123 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_963 : _GEN_675; // @[decode.scala 344:149]
  wire  _GEN_1124 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_964 : _GEN_676; // @[decode.scala 344:149]
  wire  _GEN_1125 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_965 : _GEN_677; // @[decode.scala 344:149]
  wire  _GEN_1126 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_966 : _GEN_678; // @[decode.scala 344:149]
  wire  _GEN_1127 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_967 : _GEN_679; // @[decode.scala 344:149]
  wire  _GEN_1128 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_968 : _GEN_680; // @[decode.scala 344:149]
  wire  _GEN_1129 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_969 : _GEN_681; // @[decode.scala 344:149]
  wire  _GEN_1130 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_970 : _GEN_682; // @[decode.scala 344:149]
  wire  _GEN_1131 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_971 : _GEN_683; // @[decode.scala 344:149]
  wire  _GEN_1132 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_972 : _GEN_684; // @[decode.scala 344:149]
  wire  _GEN_1133 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_973 : _GEN_685; // @[decode.scala 344:149]
  wire  _GEN_1134 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_974 : _GEN_686; // @[decode.scala 344:149]
  wire  _GEN_1135 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_975 : _GEN_687; // @[decode.scala 344:149]
  wire  _GEN_1136 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_976 : _GEN_688; // @[decode.scala 344:149]
  wire  _GEN_1137 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_977 : _GEN_689; // @[decode.scala 344:149]
  wire  _GEN_1138 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_978 : _GEN_690; // @[decode.scala 344:149]
  wire  _GEN_1139 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_979 : _GEN_691; // @[decode.scala 344:149]
  wire  _GEN_1140 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_980 : _GEN_692; // @[decode.scala 344:149]
  wire  _GEN_1141 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_981 : _GEN_693; // @[decode.scala 344:149]
  wire  _GEN_1142 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_982 : _GEN_694; // @[decode.scala 344:149]
  wire  _GEN_1143 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_983 : _GEN_695; // @[decode.scala 344:149]
  wire  _GEN_1144 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_984 : _GEN_696; // @[decode.scala 344:149]
  wire  _GEN_1145 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_985 : _GEN_697; // @[decode.scala 344:149]
  wire  _GEN_1146 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_986 : _GEN_698; // @[decode.scala 344:149]
  wire  _GEN_1147 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_987 : _GEN_699; // @[decode.scala 344:149]
  wire  _GEN_1148 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_988 : _GEN_700; // @[decode.scala 344:149]
  wire  _GEN_1149 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_989 : _GEN_701; // @[decode.scala 344:149]
  wire  _GEN_1150 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_990 : _GEN_702; // @[decode.scala 344:149]
  wire  _GEN_1151 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_991 : _GEN_703; // @[decode.scala 344:149]
  wire  _GEN_1152 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_992 : _GEN_704; // @[decode.scala 344:149]
  wire  _GEN_1153 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_993 : _GEN_705; // @[decode.scala 344:149]
  wire  _GEN_1154 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_994 : _GEN_706; // @[decode.scala 344:149]
  wire  _GEN_1155 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_995 : _GEN_707; // @[decode.scala 344:149]
  wire  _GEN_1156 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_996 : _GEN_708; // @[decode.scala 344:149]
  wire  _GEN_1157 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_997 : _GEN_709; // @[decode.scala 344:149]
  wire  _GEN_1158 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_998 : _GEN_710; // @[decode.scala 344:149]
  wire  _GEN_1159 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_999 : _GEN_711; // @[decode.scala 344:149]
  wire  _GEN_1160 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1000 : _GEN_712; // @[decode.scala 344:149]
  wire  _GEN_1161 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1001 : _GEN_713; // @[decode.scala 344:149]
  wire  _GEN_1162 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1002 : _GEN_714; // @[decode.scala 344:149]
  wire  _GEN_1163 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1003 : _GEN_715; // @[decode.scala 344:149]
  wire  _GEN_1164 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1004 : _GEN_716; // @[decode.scala 344:149]
  wire  _GEN_1165 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1005 : _GEN_717; // @[decode.scala 344:149]
  wire  _GEN_1166 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1006 : _GEN_718; // @[decode.scala 344:149]
  wire  _GEN_1167 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1007 : _GEN_719; // @[decode.scala 344:149]
  wire  _GEN_1168 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1008 : _GEN_720; // @[decode.scala 344:149]
  wire  _GEN_1169 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1009 : _GEN_721; // @[decode.scala 344:149]
  wire [5:0] _GEN_1170 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1010 : frontEndRegMap_0; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1171 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1011 : frontEndRegMap_1; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1172 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1012 : frontEndRegMap_2; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1173 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1013 : frontEndRegMap_3; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1174 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1014 : frontEndRegMap_4; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1175 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1015 : frontEndRegMap_5; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1176 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1016 : frontEndRegMap_6; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1177 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1017 : frontEndRegMap_7; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1178 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1018 : frontEndRegMap_8; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1179 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1019 : frontEndRegMap_9; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1180 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1020 : frontEndRegMap_10; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1181 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1021 : frontEndRegMap_11; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1182 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1022 : frontEndRegMap_12; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1183 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1023 : frontEndRegMap_13; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1184 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1024 : frontEndRegMap_14; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1185 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1025 : frontEndRegMap_15; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1186 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1026 : frontEndRegMap_16; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1187 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1027 : frontEndRegMap_17; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1188 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1028 : frontEndRegMap_18; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1189 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1029 : frontEndRegMap_19; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1190 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1030 : frontEndRegMap_20; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1191 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1031 : frontEndRegMap_21; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1192 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1032 : frontEndRegMap_22; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1193 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1033 : frontEndRegMap_23; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1194 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1034 : frontEndRegMap_24; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1195 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1035 : frontEndRegMap_25; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1196 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1036 : frontEndRegMap_26; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1197 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1037 : frontEndRegMap_27; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1198 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1038 : frontEndRegMap_28; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1199 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1039 : frontEndRegMap_29; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1200 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1040 : frontEndRegMap_30; // @[decode.scala 344:149 301:36]
  wire [5:0] _GEN_1201 = _T_3 & (insType_insType == 3'h1 | insType_insType == 3'h0 | insType_insType == 3'h4 |
    insType_insType == 3'h5) & inputBuffer_instruction[11:7] != 5'h0 ? _GEN_1041 : frontEndRegMap_31; // @[decode.scala 344:149 301:36]
  wire [2:0] _branchTracker_T_1 = branchTracker - 3'h1; // @[decode.scala 353:36]
  wire [3:0] _T_41 = ~branchEvalIn_branchMask; // @[decode.scala 354:75]
  wire [3:0] _T_42 = _toExec_branchMask_T & _T_41; // @[decode.scala 354:72]
  wire  _GEN_1203 = _T_424 ? 1'h0 : _T_42[0]; // @[decode.scala 354:29 356:34 359:34]
  wire  _GEN_1204 = _T_424 ? 1'h0 : _T_42[1]; // @[decode.scala 354:29 356:34 360:34]
  wire  _GEN_1205 = _T_424 ? 1'h0 : _T_42[2]; // @[decode.scala 354:29 356:34 361:34]
  wire  _GEN_1206 = _T_424 ? 1'h0 : _T_42[3]; // @[decode.scala 354:29 356:34 362:34]
  wire [63:0] _GEN_1207 = _T_424 ? branchEvalIn_targetPC : expectedPC; // @[decode.scala 356:34 363:18 183:27]
  wire  _GEN_1240 = _T_424 ? reservedFreeList1_0 | PRFFreeList_0 : _GEN_1042; // @[decode.scala 356:34 366:22]
  wire  _GEN_1241 = _T_424 ? reservedFreeList1_1 | PRFFreeList_1 : _GEN_1043; // @[decode.scala 356:34 366:22]
  wire  _GEN_1242 = _T_424 ? reservedFreeList1_2 | PRFFreeList_2 : _GEN_1044; // @[decode.scala 356:34 366:22]
  wire  _GEN_1243 = _T_424 ? reservedFreeList1_3 | PRFFreeList_3 : _GEN_1045; // @[decode.scala 356:34 366:22]
  wire  _GEN_1244 = _T_424 ? reservedFreeList1_4 | PRFFreeList_4 : _GEN_1046; // @[decode.scala 356:34 366:22]
  wire  _GEN_1245 = _T_424 ? reservedFreeList1_5 | PRFFreeList_5 : _GEN_1047; // @[decode.scala 356:34 366:22]
  wire  _GEN_1246 = _T_424 ? reservedFreeList1_6 | PRFFreeList_6 : _GEN_1048; // @[decode.scala 356:34 366:22]
  wire  _GEN_1247 = _T_424 ? reservedFreeList1_7 | PRFFreeList_7 : _GEN_1049; // @[decode.scala 356:34 366:22]
  wire  _GEN_1248 = _T_424 ? reservedFreeList1_8 | PRFFreeList_8 : _GEN_1050; // @[decode.scala 356:34 366:22]
  wire  _GEN_1249 = _T_424 ? reservedFreeList1_9 | PRFFreeList_9 : _GEN_1051; // @[decode.scala 356:34 366:22]
  wire  _GEN_1250 = _T_424 ? reservedFreeList1_10 | PRFFreeList_10 : _GEN_1052; // @[decode.scala 356:34 366:22]
  wire  _GEN_1251 = _T_424 ? reservedFreeList1_11 | PRFFreeList_11 : _GEN_1053; // @[decode.scala 356:34 366:22]
  wire  _GEN_1252 = _T_424 ? reservedFreeList1_12 | PRFFreeList_12 : _GEN_1054; // @[decode.scala 356:34 366:22]
  wire  _GEN_1253 = _T_424 ? reservedFreeList1_13 | PRFFreeList_13 : _GEN_1055; // @[decode.scala 356:34 366:22]
  wire  _GEN_1254 = _T_424 ? reservedFreeList1_14 | PRFFreeList_14 : _GEN_1056; // @[decode.scala 356:34 366:22]
  wire  _GEN_1255 = _T_424 ? reservedFreeList1_15 | PRFFreeList_15 : _GEN_1057; // @[decode.scala 356:34 366:22]
  wire  _GEN_1256 = _T_424 ? reservedFreeList1_16 | PRFFreeList_16 : _GEN_1058; // @[decode.scala 356:34 366:22]
  wire  _GEN_1257 = _T_424 ? reservedFreeList1_17 | PRFFreeList_17 : _GEN_1059; // @[decode.scala 356:34 366:22]
  wire  _GEN_1258 = _T_424 ? reservedFreeList1_18 | PRFFreeList_18 : _GEN_1060; // @[decode.scala 356:34 366:22]
  wire  _GEN_1259 = _T_424 ? reservedFreeList1_19 | PRFFreeList_19 : _GEN_1061; // @[decode.scala 356:34 366:22]
  wire  _GEN_1260 = _T_424 ? reservedFreeList1_20 | PRFFreeList_20 : _GEN_1062; // @[decode.scala 356:34 366:22]
  wire  _GEN_1261 = _T_424 ? reservedFreeList1_21 | PRFFreeList_21 : _GEN_1063; // @[decode.scala 356:34 366:22]
  wire  _GEN_1262 = _T_424 ? reservedFreeList1_22 | PRFFreeList_22 : _GEN_1064; // @[decode.scala 356:34 366:22]
  wire  _GEN_1263 = _T_424 ? reservedFreeList1_23 | PRFFreeList_23 : _GEN_1065; // @[decode.scala 356:34 366:22]
  wire  _GEN_1264 = _T_424 ? reservedFreeList1_24 | PRFFreeList_24 : _GEN_1066; // @[decode.scala 356:34 366:22]
  wire  _GEN_1265 = _T_424 ? reservedFreeList1_25 | PRFFreeList_25 : _GEN_1067; // @[decode.scala 356:34 366:22]
  wire  _GEN_1266 = _T_424 ? reservedFreeList1_26 | PRFFreeList_26 : _GEN_1068; // @[decode.scala 356:34 366:22]
  wire  _GEN_1267 = _T_424 ? reservedFreeList1_27 | PRFFreeList_27 : _GEN_1069; // @[decode.scala 356:34 366:22]
  wire  _GEN_1268 = _T_424 ? reservedFreeList1_28 | PRFFreeList_28 : _GEN_1070; // @[decode.scala 356:34 366:22]
  wire  _GEN_1269 = _T_424 ? reservedFreeList1_29 | PRFFreeList_29 : _GEN_1071; // @[decode.scala 356:34 366:22]
  wire  _GEN_1270 = _T_424 ? reservedFreeList1_30 | PRFFreeList_30 : _GEN_1072; // @[decode.scala 356:34 366:22]
  wire  _GEN_1271 = _T_424 ? reservedFreeList1_31 | PRFFreeList_31 : _GEN_1073; // @[decode.scala 356:34 366:22]
  wire  _GEN_1272 = _T_424 ? reservedFreeList1_32 | PRFFreeList_32 : _GEN_1074; // @[decode.scala 356:34 366:22]
  wire  _GEN_1273 = _T_424 ? reservedFreeList1_33 | PRFFreeList_33 : _GEN_1075; // @[decode.scala 356:34 366:22]
  wire  _GEN_1274 = _T_424 ? reservedFreeList1_34 | PRFFreeList_34 : _GEN_1076; // @[decode.scala 356:34 366:22]
  wire  _GEN_1275 = _T_424 ? reservedFreeList1_35 | PRFFreeList_35 : _GEN_1077; // @[decode.scala 356:34 366:22]
  wire  _GEN_1276 = _T_424 ? reservedFreeList1_36 | PRFFreeList_36 : _GEN_1078; // @[decode.scala 356:34 366:22]
  wire  _GEN_1277 = _T_424 ? reservedFreeList1_37 | PRFFreeList_37 : _GEN_1079; // @[decode.scala 356:34 366:22]
  wire  _GEN_1278 = _T_424 ? reservedFreeList1_38 | PRFFreeList_38 : _GEN_1080; // @[decode.scala 356:34 366:22]
  wire  _GEN_1279 = _T_424 ? reservedFreeList1_39 | PRFFreeList_39 : _GEN_1081; // @[decode.scala 356:34 366:22]
  wire  _GEN_1280 = _T_424 ? reservedFreeList1_40 | PRFFreeList_40 : _GEN_1082; // @[decode.scala 356:34 366:22]
  wire  _GEN_1281 = _T_424 ? reservedFreeList1_41 | PRFFreeList_41 : _GEN_1083; // @[decode.scala 356:34 366:22]
  wire  _GEN_1282 = _T_424 ? reservedFreeList1_42 | PRFFreeList_42 : _GEN_1084; // @[decode.scala 356:34 366:22]
  wire  _GEN_1283 = _T_424 ? reservedFreeList1_43 | PRFFreeList_43 : _GEN_1085; // @[decode.scala 356:34 366:22]
  wire  _GEN_1284 = _T_424 ? reservedFreeList1_44 | PRFFreeList_44 : _GEN_1086; // @[decode.scala 356:34 366:22]
  wire  _GEN_1285 = _T_424 ? reservedFreeList1_45 | PRFFreeList_45 : _GEN_1087; // @[decode.scala 356:34 366:22]
  wire  _GEN_1286 = _T_424 ? reservedFreeList1_46 | PRFFreeList_46 : _GEN_1088; // @[decode.scala 356:34 366:22]
  wire  _GEN_1287 = _T_424 ? reservedFreeList1_47 | PRFFreeList_47 : _GEN_1089; // @[decode.scala 356:34 366:22]
  wire  _GEN_1288 = _T_424 ? reservedFreeList1_48 | PRFFreeList_48 : _GEN_1090; // @[decode.scala 356:34 366:22]
  wire  _GEN_1289 = _T_424 ? reservedFreeList1_49 | PRFFreeList_49 : _GEN_1091; // @[decode.scala 356:34 366:22]
  wire  _GEN_1290 = _T_424 ? reservedFreeList1_50 | PRFFreeList_50 : _GEN_1092; // @[decode.scala 356:34 366:22]
  wire  _GEN_1291 = _T_424 ? reservedFreeList1_51 | PRFFreeList_51 : _GEN_1093; // @[decode.scala 356:34 366:22]
  wire  _GEN_1292 = _T_424 ? reservedFreeList1_52 | PRFFreeList_52 : _GEN_1094; // @[decode.scala 356:34 366:22]
  wire  _GEN_1293 = _T_424 ? reservedFreeList1_53 | PRFFreeList_53 : _GEN_1095; // @[decode.scala 356:34 366:22]
  wire  _GEN_1294 = _T_424 ? reservedFreeList1_54 | PRFFreeList_54 : _GEN_1096; // @[decode.scala 356:34 366:22]
  wire  _GEN_1295 = _T_424 ? reservedFreeList1_55 | PRFFreeList_55 : _GEN_1097; // @[decode.scala 356:34 366:22]
  wire  _GEN_1296 = _T_424 ? reservedFreeList1_56 | PRFFreeList_56 : _GEN_1098; // @[decode.scala 356:34 366:22]
  wire  _GEN_1297 = _T_424 ? reservedFreeList1_57 | PRFFreeList_57 : _GEN_1099; // @[decode.scala 356:34 366:22]
  wire  _GEN_1298 = _T_424 ? reservedFreeList1_58 | PRFFreeList_58 : _GEN_1100; // @[decode.scala 356:34 366:22]
  wire  _GEN_1299 = _T_424 ? reservedFreeList1_59 | PRFFreeList_59 : _GEN_1101; // @[decode.scala 356:34 366:22]
  wire  _GEN_1300 = _T_424 ? reservedFreeList1_60 | PRFFreeList_60 : _GEN_1102; // @[decode.scala 356:34 366:22]
  wire  _GEN_1301 = _T_424 ? reservedFreeList1_61 | PRFFreeList_61 : _GEN_1103; // @[decode.scala 356:34 366:22]
  wire  _GEN_1302 = _T_424 ? reservedFreeList1_62 | PRFFreeList_62 : _GEN_1104; // @[decode.scala 356:34 366:22]
  wire  _GEN_1304 = _T_424 ? reservedValidList1_0 | PRFValidList_0 : _GEN_1106; // @[decode.scala 356:34 367:22]
  wire  _GEN_1305 = _T_424 ? reservedValidList1_1 | PRFValidList_1 : _GEN_1107; // @[decode.scala 356:34 367:22]
  wire  _GEN_1306 = _T_424 ? reservedValidList1_2 | PRFValidList_2 : _GEN_1108; // @[decode.scala 356:34 367:22]
  wire  _GEN_1307 = _T_424 ? reservedValidList1_3 | PRFValidList_3 : _GEN_1109; // @[decode.scala 356:34 367:22]
  wire  _GEN_1308 = _T_424 ? reservedValidList1_4 | PRFValidList_4 : _GEN_1110; // @[decode.scala 356:34 367:22]
  wire  _GEN_1309 = _T_424 ? reservedValidList1_5 | PRFValidList_5 : _GEN_1111; // @[decode.scala 356:34 367:22]
  wire  _GEN_1310 = _T_424 ? reservedValidList1_6 | PRFValidList_6 : _GEN_1112; // @[decode.scala 356:34 367:22]
  wire  _GEN_1311 = _T_424 ? reservedValidList1_7 | PRFValidList_7 : _GEN_1113; // @[decode.scala 356:34 367:22]
  wire  _GEN_1312 = _T_424 ? reservedValidList1_8 | PRFValidList_8 : _GEN_1114; // @[decode.scala 356:34 367:22]
  wire  _GEN_1313 = _T_424 ? reservedValidList1_9 | PRFValidList_9 : _GEN_1115; // @[decode.scala 356:34 367:22]
  wire  _GEN_1314 = _T_424 ? reservedValidList1_10 | PRFValidList_10 : _GEN_1116; // @[decode.scala 356:34 367:22]
  wire  _GEN_1315 = _T_424 ? reservedValidList1_11 | PRFValidList_11 : _GEN_1117; // @[decode.scala 356:34 367:22]
  wire  _GEN_1316 = _T_424 ? reservedValidList1_12 | PRFValidList_12 : _GEN_1118; // @[decode.scala 356:34 367:22]
  wire  _GEN_1317 = _T_424 ? reservedValidList1_13 | PRFValidList_13 : _GEN_1119; // @[decode.scala 356:34 367:22]
  wire  _GEN_1318 = _T_424 ? reservedValidList1_14 | PRFValidList_14 : _GEN_1120; // @[decode.scala 356:34 367:22]
  wire  _GEN_1319 = _T_424 ? reservedValidList1_15 | PRFValidList_15 : _GEN_1121; // @[decode.scala 356:34 367:22]
  wire  _GEN_1320 = _T_424 ? reservedValidList1_16 | PRFValidList_16 : _GEN_1122; // @[decode.scala 356:34 367:22]
  wire  _GEN_1321 = _T_424 ? reservedValidList1_17 | PRFValidList_17 : _GEN_1123; // @[decode.scala 356:34 367:22]
  wire  _GEN_1322 = _T_424 ? reservedValidList1_18 | PRFValidList_18 : _GEN_1124; // @[decode.scala 356:34 367:22]
  wire  _GEN_1323 = _T_424 ? reservedValidList1_19 | PRFValidList_19 : _GEN_1125; // @[decode.scala 356:34 367:22]
  wire  _GEN_1324 = _T_424 ? reservedValidList1_20 | PRFValidList_20 : _GEN_1126; // @[decode.scala 356:34 367:22]
  wire  _GEN_1325 = _T_424 ? reservedValidList1_21 | PRFValidList_21 : _GEN_1127; // @[decode.scala 356:34 367:22]
  wire  _GEN_1326 = _T_424 ? reservedValidList1_22 | PRFValidList_22 : _GEN_1128; // @[decode.scala 356:34 367:22]
  wire  _GEN_1327 = _T_424 ? reservedValidList1_23 | PRFValidList_23 : _GEN_1129; // @[decode.scala 356:34 367:22]
  wire  _GEN_1328 = _T_424 ? reservedValidList1_24 | PRFValidList_24 : _GEN_1130; // @[decode.scala 356:34 367:22]
  wire  _GEN_1329 = _T_424 ? reservedValidList1_25 | PRFValidList_25 : _GEN_1131; // @[decode.scala 356:34 367:22]
  wire  _GEN_1330 = _T_424 ? reservedValidList1_26 | PRFValidList_26 : _GEN_1132; // @[decode.scala 356:34 367:22]
  wire  _GEN_1331 = _T_424 ? reservedValidList1_27 | PRFValidList_27 : _GEN_1133; // @[decode.scala 356:34 367:22]
  wire  _GEN_1332 = _T_424 ? reservedValidList1_28 | PRFValidList_28 : _GEN_1134; // @[decode.scala 356:34 367:22]
  wire  _GEN_1333 = _T_424 ? reservedValidList1_29 | PRFValidList_29 : _GEN_1135; // @[decode.scala 356:34 367:22]
  wire  _GEN_1334 = _T_424 ? reservedValidList1_30 | PRFValidList_30 : _GEN_1136; // @[decode.scala 356:34 367:22]
  wire  _GEN_1335 = _T_424 ? reservedValidList1_31 | PRFValidList_31 : _GEN_1137; // @[decode.scala 356:34 367:22]
  wire  _GEN_1336 = _T_424 ? reservedValidList1_32 | PRFValidList_32 : _GEN_1138; // @[decode.scala 356:34 367:22]
  wire  _GEN_1337 = _T_424 ? reservedValidList1_33 | PRFValidList_33 : _GEN_1139; // @[decode.scala 356:34 367:22]
  wire  _GEN_1338 = _T_424 ? reservedValidList1_34 | PRFValidList_34 : _GEN_1140; // @[decode.scala 356:34 367:22]
  wire  _GEN_1339 = _T_424 ? reservedValidList1_35 | PRFValidList_35 : _GEN_1141; // @[decode.scala 356:34 367:22]
  wire  _GEN_1340 = _T_424 ? reservedValidList1_36 | PRFValidList_36 : _GEN_1142; // @[decode.scala 356:34 367:22]
  wire  _GEN_1341 = _T_424 ? reservedValidList1_37 | PRFValidList_37 : _GEN_1143; // @[decode.scala 356:34 367:22]
  wire  _GEN_1342 = _T_424 ? reservedValidList1_38 | PRFValidList_38 : _GEN_1144; // @[decode.scala 356:34 367:22]
  wire  _GEN_1343 = _T_424 ? reservedValidList1_39 | PRFValidList_39 : _GEN_1145; // @[decode.scala 356:34 367:22]
  wire  _GEN_1344 = _T_424 ? reservedValidList1_40 | PRFValidList_40 : _GEN_1146; // @[decode.scala 356:34 367:22]
  wire  _GEN_1345 = _T_424 ? reservedValidList1_41 | PRFValidList_41 : _GEN_1147; // @[decode.scala 356:34 367:22]
  wire  _GEN_1346 = _T_424 ? reservedValidList1_42 | PRFValidList_42 : _GEN_1148; // @[decode.scala 356:34 367:22]
  wire  _GEN_1347 = _T_424 ? reservedValidList1_43 | PRFValidList_43 : _GEN_1149; // @[decode.scala 356:34 367:22]
  wire  _GEN_1348 = _T_424 ? reservedValidList1_44 | PRFValidList_44 : _GEN_1150; // @[decode.scala 356:34 367:22]
  wire  _GEN_1349 = _T_424 ? reservedValidList1_45 | PRFValidList_45 : _GEN_1151; // @[decode.scala 356:34 367:22]
  wire  _GEN_1350 = _T_424 ? reservedValidList1_46 | PRFValidList_46 : _GEN_1152; // @[decode.scala 356:34 367:22]
  wire  _GEN_1351 = _T_424 ? reservedValidList1_47 | PRFValidList_47 : _GEN_1153; // @[decode.scala 356:34 367:22]
  wire  _GEN_1352 = _T_424 ? reservedValidList1_48 | PRFValidList_48 : _GEN_1154; // @[decode.scala 356:34 367:22]
  wire  _GEN_1353 = _T_424 ? reservedValidList1_49 | PRFValidList_49 : _GEN_1155; // @[decode.scala 356:34 367:22]
  wire  _GEN_1354 = _T_424 ? reservedValidList1_50 | PRFValidList_50 : _GEN_1156; // @[decode.scala 356:34 367:22]
  wire  _GEN_1355 = _T_424 ? reservedValidList1_51 | PRFValidList_51 : _GEN_1157; // @[decode.scala 356:34 367:22]
  wire  _GEN_1356 = _T_424 ? reservedValidList1_52 | PRFValidList_52 : _GEN_1158; // @[decode.scala 356:34 367:22]
  wire  _GEN_1357 = _T_424 ? reservedValidList1_53 | PRFValidList_53 : _GEN_1159; // @[decode.scala 356:34 367:22]
  wire  _GEN_1358 = _T_424 ? reservedValidList1_54 | PRFValidList_54 : _GEN_1160; // @[decode.scala 356:34 367:22]
  wire  _GEN_1359 = _T_424 ? reservedValidList1_55 | PRFValidList_55 : _GEN_1161; // @[decode.scala 356:34 367:22]
  wire  _GEN_1360 = _T_424 ? reservedValidList1_56 | PRFValidList_56 : _GEN_1162; // @[decode.scala 356:34 367:22]
  wire  _GEN_1361 = _T_424 ? reservedValidList1_57 | PRFValidList_57 : _GEN_1163; // @[decode.scala 356:34 367:22]
  wire  _GEN_1362 = _T_424 ? reservedValidList1_58 | PRFValidList_58 : _GEN_1164; // @[decode.scala 356:34 367:22]
  wire  _GEN_1363 = _T_424 ? reservedValidList1_59 | PRFValidList_59 : _GEN_1165; // @[decode.scala 356:34 367:22]
  wire  _GEN_1364 = _T_424 ? reservedValidList1_60 | PRFValidList_60 : _GEN_1166; // @[decode.scala 356:34 367:22]
  wire  _GEN_1365 = _T_424 ? reservedValidList1_61 | PRFValidList_61 : _GEN_1167; // @[decode.scala 356:34 367:22]
  wire  _GEN_1366 = _T_424 ? reservedValidList1_62 | PRFValidList_62 : _GEN_1168; // @[decode.scala 356:34 367:22]
  wire  _GEN_1367 = _T_424 ? reservedValidList1_63 | PRFValidList_63 : _GEN_1169; // @[decode.scala 356:34 367:22]
  wire [2:0] _GEN_1368 = _T_424 ? 3'h0 : _branchTracker_T_1; // @[decode.scala 353:19 356:34 369:21]
  wire [5:0] _GEN_1369 = _T_424 ? reservedRegMap1_0 : reservedRegMap2_0; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1370 = _T_424 ? reservedRegMap1_1 : reservedRegMap2_1; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1371 = _T_424 ? reservedRegMap1_2 : reservedRegMap2_2; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1372 = _T_424 ? reservedRegMap1_3 : reservedRegMap2_3; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1373 = _T_424 ? reservedRegMap1_4 : reservedRegMap2_4; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1374 = _T_424 ? reservedRegMap1_5 : reservedRegMap2_5; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1375 = _T_424 ? reservedRegMap1_6 : reservedRegMap2_6; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1376 = _T_424 ? reservedRegMap1_7 : reservedRegMap2_7; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1377 = _T_424 ? reservedRegMap1_8 : reservedRegMap2_8; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1378 = _T_424 ? reservedRegMap1_9 : reservedRegMap2_9; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1379 = _T_424 ? reservedRegMap1_10 : reservedRegMap2_10; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1380 = _T_424 ? reservedRegMap1_11 : reservedRegMap2_11; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1381 = _T_424 ? reservedRegMap1_12 : reservedRegMap2_12; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1382 = _T_424 ? reservedRegMap1_13 : reservedRegMap2_13; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1383 = _T_424 ? reservedRegMap1_14 : reservedRegMap2_14; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1384 = _T_424 ? reservedRegMap1_15 : reservedRegMap2_15; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1385 = _T_424 ? reservedRegMap1_16 : reservedRegMap2_16; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1386 = _T_424 ? reservedRegMap1_17 : reservedRegMap2_17; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1387 = _T_424 ? reservedRegMap1_18 : reservedRegMap2_18; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1388 = _T_424 ? reservedRegMap1_19 : reservedRegMap2_19; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1389 = _T_424 ? reservedRegMap1_20 : reservedRegMap2_20; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1390 = _T_424 ? reservedRegMap1_21 : reservedRegMap2_21; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1391 = _T_424 ? reservedRegMap1_22 : reservedRegMap2_22; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1392 = _T_424 ? reservedRegMap1_23 : reservedRegMap2_23; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1393 = _T_424 ? reservedRegMap1_24 : reservedRegMap2_24; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1394 = _T_424 ? reservedRegMap1_25 : reservedRegMap2_25; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1395 = _T_424 ? reservedRegMap1_26 : reservedRegMap2_26; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1396 = _T_424 ? reservedRegMap1_27 : reservedRegMap2_27; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1397 = _T_424 ? reservedRegMap1_28 : reservedRegMap2_28; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1398 = _T_424 ? reservedRegMap1_29 : reservedRegMap2_29; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1399 = _T_424 ? reservedRegMap1_30 : reservedRegMap2_30; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1400 = _T_424 ? reservedRegMap1_31 : reservedRegMap2_31; // @[decode.scala 310:28 356:34 371:23]
  wire [5:0] _GEN_1401 = _T_424 ? reservedRegMap2_0 : reservedRegMap3_0; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1402 = _T_424 ? reservedRegMap2_1 : reservedRegMap3_1; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1403 = _T_424 ? reservedRegMap2_2 : reservedRegMap3_2; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1404 = _T_424 ? reservedRegMap2_3 : reservedRegMap3_3; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1405 = _T_424 ? reservedRegMap2_4 : reservedRegMap3_4; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1406 = _T_424 ? reservedRegMap2_5 : reservedRegMap3_5; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1407 = _T_424 ? reservedRegMap2_6 : reservedRegMap3_6; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1408 = _T_424 ? reservedRegMap2_7 : reservedRegMap3_7; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1409 = _T_424 ? reservedRegMap2_8 : reservedRegMap3_8; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1410 = _T_424 ? reservedRegMap2_9 : reservedRegMap3_9; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1411 = _T_424 ? reservedRegMap2_10 : reservedRegMap3_10; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1412 = _T_424 ? reservedRegMap2_11 : reservedRegMap3_11; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1413 = _T_424 ? reservedRegMap2_12 : reservedRegMap3_12; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1414 = _T_424 ? reservedRegMap2_13 : reservedRegMap3_13; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1415 = _T_424 ? reservedRegMap2_14 : reservedRegMap3_14; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1416 = _T_424 ? reservedRegMap2_15 : reservedRegMap3_15; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1417 = _T_424 ? reservedRegMap2_16 : reservedRegMap3_16; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1418 = _T_424 ? reservedRegMap2_17 : reservedRegMap3_17; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1419 = _T_424 ? reservedRegMap2_18 : reservedRegMap3_18; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1420 = _T_424 ? reservedRegMap2_19 : reservedRegMap3_19; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1421 = _T_424 ? reservedRegMap2_20 : reservedRegMap3_20; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1422 = _T_424 ? reservedRegMap2_21 : reservedRegMap3_21; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1423 = _T_424 ? reservedRegMap2_22 : reservedRegMap3_22; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1424 = _T_424 ? reservedRegMap2_23 : reservedRegMap3_23; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1425 = _T_424 ? reservedRegMap2_24 : reservedRegMap3_24; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1426 = _T_424 ? reservedRegMap2_25 : reservedRegMap3_25; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1427 = _T_424 ? reservedRegMap2_26 : reservedRegMap3_26; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1428 = _T_424 ? reservedRegMap2_27 : reservedRegMap3_27; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1429 = _T_424 ? reservedRegMap2_28 : reservedRegMap3_28; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1430 = _T_424 ? reservedRegMap2_29 : reservedRegMap3_29; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1431 = _T_424 ? reservedRegMap2_30 : reservedRegMap3_30; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1432 = _T_424 ? reservedRegMap2_31 : reservedRegMap3_31; // @[decode.scala 311:28 356:34 372:23]
  wire [5:0] _GEN_1433 = _T_424 ? reservedRegMap3_0 : reservedRegMap4_0; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1434 = _T_424 ? reservedRegMap3_1 : reservedRegMap4_1; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1435 = _T_424 ? reservedRegMap3_2 : reservedRegMap4_2; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1436 = _T_424 ? reservedRegMap3_3 : reservedRegMap4_3; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1437 = _T_424 ? reservedRegMap3_4 : reservedRegMap4_4; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1438 = _T_424 ? reservedRegMap3_5 : reservedRegMap4_5; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1439 = _T_424 ? reservedRegMap3_6 : reservedRegMap4_6; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1440 = _T_424 ? reservedRegMap3_7 : reservedRegMap4_7; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1441 = _T_424 ? reservedRegMap3_8 : reservedRegMap4_8; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1442 = _T_424 ? reservedRegMap3_9 : reservedRegMap4_9; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1443 = _T_424 ? reservedRegMap3_10 : reservedRegMap4_10; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1444 = _T_424 ? reservedRegMap3_11 : reservedRegMap4_11; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1445 = _T_424 ? reservedRegMap3_12 : reservedRegMap4_12; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1446 = _T_424 ? reservedRegMap3_13 : reservedRegMap4_13; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1447 = _T_424 ? reservedRegMap3_14 : reservedRegMap4_14; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1448 = _T_424 ? reservedRegMap3_15 : reservedRegMap4_15; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1449 = _T_424 ? reservedRegMap3_16 : reservedRegMap4_16; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1450 = _T_424 ? reservedRegMap3_17 : reservedRegMap4_17; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1451 = _T_424 ? reservedRegMap3_18 : reservedRegMap4_18; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1452 = _T_424 ? reservedRegMap3_19 : reservedRegMap4_19; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1453 = _T_424 ? reservedRegMap3_20 : reservedRegMap4_20; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1454 = _T_424 ? reservedRegMap3_21 : reservedRegMap4_21; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1455 = _T_424 ? reservedRegMap3_22 : reservedRegMap4_22; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1456 = _T_424 ? reservedRegMap3_23 : reservedRegMap4_23; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1457 = _T_424 ? reservedRegMap3_24 : reservedRegMap4_24; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1458 = _T_424 ? reservedRegMap3_25 : reservedRegMap4_25; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1459 = _T_424 ? reservedRegMap3_26 : reservedRegMap4_26; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1460 = _T_424 ? reservedRegMap3_27 : reservedRegMap4_27; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1461 = _T_424 ? reservedRegMap3_28 : reservedRegMap4_28; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1462 = _T_424 ? reservedRegMap3_29 : reservedRegMap4_29; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1463 = _T_424 ? reservedRegMap3_30 : reservedRegMap4_30; // @[decode.scala 312:28 356:34 373:23]
  wire [5:0] _GEN_1464 = _T_424 ? reservedRegMap3_31 : reservedRegMap4_31; // @[decode.scala 312:28 356:34 373:23]
  wire  _GEN_1465 = _T_424 ? reservedFreeList1_0 : reservedFreeList2_0; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1466 = _T_424 ? reservedFreeList1_1 : reservedFreeList2_1; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1467 = _T_424 ? reservedFreeList1_2 : reservedFreeList2_2; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1468 = _T_424 ? reservedFreeList1_3 : reservedFreeList2_3; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1469 = _T_424 ? reservedFreeList1_4 : reservedFreeList2_4; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1470 = _T_424 ? reservedFreeList1_5 : reservedFreeList2_5; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1471 = _T_424 ? reservedFreeList1_6 : reservedFreeList2_6; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1472 = _T_424 ? reservedFreeList1_7 : reservedFreeList2_7; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1473 = _T_424 ? reservedFreeList1_8 : reservedFreeList2_8; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1474 = _T_424 ? reservedFreeList1_9 : reservedFreeList2_9; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1475 = _T_424 ? reservedFreeList1_10 : reservedFreeList2_10; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1476 = _T_424 ? reservedFreeList1_11 : reservedFreeList2_11; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1477 = _T_424 ? reservedFreeList1_12 : reservedFreeList2_12; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1478 = _T_424 ? reservedFreeList1_13 : reservedFreeList2_13; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1479 = _T_424 ? reservedFreeList1_14 : reservedFreeList2_14; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1480 = _T_424 ? reservedFreeList1_15 : reservedFreeList2_15; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1481 = _T_424 ? reservedFreeList1_16 : reservedFreeList2_16; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1482 = _T_424 ? reservedFreeList1_17 : reservedFreeList2_17; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1483 = _T_424 ? reservedFreeList1_18 : reservedFreeList2_18; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1484 = _T_424 ? reservedFreeList1_19 : reservedFreeList2_19; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1485 = _T_424 ? reservedFreeList1_20 : reservedFreeList2_20; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1486 = _T_424 ? reservedFreeList1_21 : reservedFreeList2_21; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1487 = _T_424 ? reservedFreeList1_22 : reservedFreeList2_22; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1488 = _T_424 ? reservedFreeList1_23 : reservedFreeList2_23; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1489 = _T_424 ? reservedFreeList1_24 : reservedFreeList2_24; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1490 = _T_424 ? reservedFreeList1_25 : reservedFreeList2_25; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1491 = _T_424 ? reservedFreeList1_26 : reservedFreeList2_26; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1492 = _T_424 ? reservedFreeList1_27 : reservedFreeList2_27; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1493 = _T_424 ? reservedFreeList1_28 : reservedFreeList2_28; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1494 = _T_424 ? reservedFreeList1_29 : reservedFreeList2_29; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1495 = _T_424 ? reservedFreeList1_30 : reservedFreeList2_30; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1496 = _T_424 ? reservedFreeList1_31 : reservedFreeList2_31; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1497 = _T_424 ? reservedFreeList1_32 : reservedFreeList2_32; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1498 = _T_424 ? reservedFreeList1_33 : reservedFreeList2_33; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1499 = _T_424 ? reservedFreeList1_34 : reservedFreeList2_34; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1500 = _T_424 ? reservedFreeList1_35 : reservedFreeList2_35; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1501 = _T_424 ? reservedFreeList1_36 : reservedFreeList2_36; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1502 = _T_424 ? reservedFreeList1_37 : reservedFreeList2_37; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1503 = _T_424 ? reservedFreeList1_38 : reservedFreeList2_38; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1504 = _T_424 ? reservedFreeList1_39 : reservedFreeList2_39; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1505 = _T_424 ? reservedFreeList1_40 : reservedFreeList2_40; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1506 = _T_424 ? reservedFreeList1_41 : reservedFreeList2_41; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1507 = _T_424 ? reservedFreeList1_42 : reservedFreeList2_42; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1508 = _T_424 ? reservedFreeList1_43 : reservedFreeList2_43; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1509 = _T_424 ? reservedFreeList1_44 : reservedFreeList2_44; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1510 = _T_424 ? reservedFreeList1_45 : reservedFreeList2_45; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1511 = _T_424 ? reservedFreeList1_46 : reservedFreeList2_46; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1512 = _T_424 ? reservedFreeList1_47 : reservedFreeList2_47; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1513 = _T_424 ? reservedFreeList1_48 : reservedFreeList2_48; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1514 = _T_424 ? reservedFreeList1_49 : reservedFreeList2_49; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1515 = _T_424 ? reservedFreeList1_50 : reservedFreeList2_50; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1516 = _T_424 ? reservedFreeList1_51 : reservedFreeList2_51; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1517 = _T_424 ? reservedFreeList1_52 : reservedFreeList2_52; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1518 = _T_424 ? reservedFreeList1_53 : reservedFreeList2_53; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1519 = _T_424 ? reservedFreeList1_54 : reservedFreeList2_54; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1520 = _T_424 ? reservedFreeList1_55 : reservedFreeList2_55; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1521 = _T_424 ? reservedFreeList1_56 : reservedFreeList2_56; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1522 = _T_424 ? reservedFreeList1_57 : reservedFreeList2_57; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1523 = _T_424 ? reservedFreeList1_58 : reservedFreeList2_58; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1524 = _T_424 ? reservedFreeList1_59 : reservedFreeList2_59; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1525 = _T_424 ? reservedFreeList1_60 : reservedFreeList2_60; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1526 = _T_424 ? reservedFreeList1_61 : reservedFreeList2_61; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1527 = _T_424 ? reservedFreeList1_62 : reservedFreeList2_62; // @[decode.scala 315:30 356:34 375:25]
  wire  _GEN_1529 = _T_424 ? reservedFreeList2_0 : reservedFreeList3_0; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1530 = _T_424 ? reservedFreeList2_1 : reservedFreeList3_1; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1531 = _T_424 ? reservedFreeList2_2 : reservedFreeList3_2; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1532 = _T_424 ? reservedFreeList2_3 : reservedFreeList3_3; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1533 = _T_424 ? reservedFreeList2_4 : reservedFreeList3_4; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1534 = _T_424 ? reservedFreeList2_5 : reservedFreeList3_5; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1535 = _T_424 ? reservedFreeList2_6 : reservedFreeList3_6; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1536 = _T_424 ? reservedFreeList2_7 : reservedFreeList3_7; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1537 = _T_424 ? reservedFreeList2_8 : reservedFreeList3_8; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1538 = _T_424 ? reservedFreeList2_9 : reservedFreeList3_9; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1539 = _T_424 ? reservedFreeList2_10 : reservedFreeList3_10; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1540 = _T_424 ? reservedFreeList2_11 : reservedFreeList3_11; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1541 = _T_424 ? reservedFreeList2_12 : reservedFreeList3_12; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1542 = _T_424 ? reservedFreeList2_13 : reservedFreeList3_13; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1543 = _T_424 ? reservedFreeList2_14 : reservedFreeList3_14; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1544 = _T_424 ? reservedFreeList2_15 : reservedFreeList3_15; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1545 = _T_424 ? reservedFreeList2_16 : reservedFreeList3_16; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1546 = _T_424 ? reservedFreeList2_17 : reservedFreeList3_17; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1547 = _T_424 ? reservedFreeList2_18 : reservedFreeList3_18; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1548 = _T_424 ? reservedFreeList2_19 : reservedFreeList3_19; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1549 = _T_424 ? reservedFreeList2_20 : reservedFreeList3_20; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1550 = _T_424 ? reservedFreeList2_21 : reservedFreeList3_21; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1551 = _T_424 ? reservedFreeList2_22 : reservedFreeList3_22; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1552 = _T_424 ? reservedFreeList2_23 : reservedFreeList3_23; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1553 = _T_424 ? reservedFreeList2_24 : reservedFreeList3_24; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1554 = _T_424 ? reservedFreeList2_25 : reservedFreeList3_25; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1555 = _T_424 ? reservedFreeList2_26 : reservedFreeList3_26; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1556 = _T_424 ? reservedFreeList2_27 : reservedFreeList3_27; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1557 = _T_424 ? reservedFreeList2_28 : reservedFreeList3_28; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1558 = _T_424 ? reservedFreeList2_29 : reservedFreeList3_29; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1559 = _T_424 ? reservedFreeList2_30 : reservedFreeList3_30; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1560 = _T_424 ? reservedFreeList2_31 : reservedFreeList3_31; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1561 = _T_424 ? reservedFreeList2_32 : reservedFreeList3_32; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1562 = _T_424 ? reservedFreeList2_33 : reservedFreeList3_33; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1563 = _T_424 ? reservedFreeList2_34 : reservedFreeList3_34; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1564 = _T_424 ? reservedFreeList2_35 : reservedFreeList3_35; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1565 = _T_424 ? reservedFreeList2_36 : reservedFreeList3_36; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1566 = _T_424 ? reservedFreeList2_37 : reservedFreeList3_37; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1567 = _T_424 ? reservedFreeList2_38 : reservedFreeList3_38; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1568 = _T_424 ? reservedFreeList2_39 : reservedFreeList3_39; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1569 = _T_424 ? reservedFreeList2_40 : reservedFreeList3_40; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1570 = _T_424 ? reservedFreeList2_41 : reservedFreeList3_41; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1571 = _T_424 ? reservedFreeList2_42 : reservedFreeList3_42; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1572 = _T_424 ? reservedFreeList2_43 : reservedFreeList3_43; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1573 = _T_424 ? reservedFreeList2_44 : reservedFreeList3_44; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1574 = _T_424 ? reservedFreeList2_45 : reservedFreeList3_45; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1575 = _T_424 ? reservedFreeList2_46 : reservedFreeList3_46; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1576 = _T_424 ? reservedFreeList2_47 : reservedFreeList3_47; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1577 = _T_424 ? reservedFreeList2_48 : reservedFreeList3_48; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1578 = _T_424 ? reservedFreeList2_49 : reservedFreeList3_49; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1579 = _T_424 ? reservedFreeList2_50 : reservedFreeList3_50; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1580 = _T_424 ? reservedFreeList2_51 : reservedFreeList3_51; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1581 = _T_424 ? reservedFreeList2_52 : reservedFreeList3_52; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1582 = _T_424 ? reservedFreeList2_53 : reservedFreeList3_53; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1583 = _T_424 ? reservedFreeList2_54 : reservedFreeList3_54; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1584 = _T_424 ? reservedFreeList2_55 : reservedFreeList3_55; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1585 = _T_424 ? reservedFreeList2_56 : reservedFreeList3_56; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1586 = _T_424 ? reservedFreeList2_57 : reservedFreeList3_57; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1587 = _T_424 ? reservedFreeList2_58 : reservedFreeList3_58; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1588 = _T_424 ? reservedFreeList2_59 : reservedFreeList3_59; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1589 = _T_424 ? reservedFreeList2_60 : reservedFreeList3_60; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1590 = _T_424 ? reservedFreeList2_61 : reservedFreeList3_61; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1591 = _T_424 ? reservedFreeList2_62 : reservedFreeList3_62; // @[decode.scala 316:30 356:34 376:25]
  wire  _GEN_1593 = _T_424 ? reservedFreeList3_0 : reservedFreeList4_0; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1594 = _T_424 ? reservedFreeList3_1 : reservedFreeList4_1; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1595 = _T_424 ? reservedFreeList3_2 : reservedFreeList4_2; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1596 = _T_424 ? reservedFreeList3_3 : reservedFreeList4_3; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1597 = _T_424 ? reservedFreeList3_4 : reservedFreeList4_4; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1598 = _T_424 ? reservedFreeList3_5 : reservedFreeList4_5; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1599 = _T_424 ? reservedFreeList3_6 : reservedFreeList4_6; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1600 = _T_424 ? reservedFreeList3_7 : reservedFreeList4_7; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1601 = _T_424 ? reservedFreeList3_8 : reservedFreeList4_8; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1602 = _T_424 ? reservedFreeList3_9 : reservedFreeList4_9; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1603 = _T_424 ? reservedFreeList3_10 : reservedFreeList4_10; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1604 = _T_424 ? reservedFreeList3_11 : reservedFreeList4_11; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1605 = _T_424 ? reservedFreeList3_12 : reservedFreeList4_12; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1606 = _T_424 ? reservedFreeList3_13 : reservedFreeList4_13; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1607 = _T_424 ? reservedFreeList3_14 : reservedFreeList4_14; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1608 = _T_424 ? reservedFreeList3_15 : reservedFreeList4_15; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1609 = _T_424 ? reservedFreeList3_16 : reservedFreeList4_16; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1610 = _T_424 ? reservedFreeList3_17 : reservedFreeList4_17; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1611 = _T_424 ? reservedFreeList3_18 : reservedFreeList4_18; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1612 = _T_424 ? reservedFreeList3_19 : reservedFreeList4_19; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1613 = _T_424 ? reservedFreeList3_20 : reservedFreeList4_20; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1614 = _T_424 ? reservedFreeList3_21 : reservedFreeList4_21; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1615 = _T_424 ? reservedFreeList3_22 : reservedFreeList4_22; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1616 = _T_424 ? reservedFreeList3_23 : reservedFreeList4_23; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1617 = _T_424 ? reservedFreeList3_24 : reservedFreeList4_24; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1618 = _T_424 ? reservedFreeList3_25 : reservedFreeList4_25; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1619 = _T_424 ? reservedFreeList3_26 : reservedFreeList4_26; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1620 = _T_424 ? reservedFreeList3_27 : reservedFreeList4_27; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1621 = _T_424 ? reservedFreeList3_28 : reservedFreeList4_28; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1622 = _T_424 ? reservedFreeList3_29 : reservedFreeList4_29; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1623 = _T_424 ? reservedFreeList3_30 : reservedFreeList4_30; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1624 = _T_424 ? reservedFreeList3_31 : reservedFreeList4_31; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1625 = _T_424 ? reservedFreeList3_32 : reservedFreeList4_32; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1626 = _T_424 ? reservedFreeList3_33 : reservedFreeList4_33; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1627 = _T_424 ? reservedFreeList3_34 : reservedFreeList4_34; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1628 = _T_424 ? reservedFreeList3_35 : reservedFreeList4_35; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1629 = _T_424 ? reservedFreeList3_36 : reservedFreeList4_36; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1630 = _T_424 ? reservedFreeList3_37 : reservedFreeList4_37; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1631 = _T_424 ? reservedFreeList3_38 : reservedFreeList4_38; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1632 = _T_424 ? reservedFreeList3_39 : reservedFreeList4_39; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1633 = _T_424 ? reservedFreeList3_40 : reservedFreeList4_40; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1634 = _T_424 ? reservedFreeList3_41 : reservedFreeList4_41; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1635 = _T_424 ? reservedFreeList3_42 : reservedFreeList4_42; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1636 = _T_424 ? reservedFreeList3_43 : reservedFreeList4_43; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1637 = _T_424 ? reservedFreeList3_44 : reservedFreeList4_44; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1638 = _T_424 ? reservedFreeList3_45 : reservedFreeList4_45; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1639 = _T_424 ? reservedFreeList3_46 : reservedFreeList4_46; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1640 = _T_424 ? reservedFreeList3_47 : reservedFreeList4_47; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1641 = _T_424 ? reservedFreeList3_48 : reservedFreeList4_48; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1642 = _T_424 ? reservedFreeList3_49 : reservedFreeList4_49; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1643 = _T_424 ? reservedFreeList3_50 : reservedFreeList4_50; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1644 = _T_424 ? reservedFreeList3_51 : reservedFreeList4_51; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1645 = _T_424 ? reservedFreeList3_52 : reservedFreeList4_52; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1646 = _T_424 ? reservedFreeList3_53 : reservedFreeList4_53; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1647 = _T_424 ? reservedFreeList3_54 : reservedFreeList4_54; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1648 = _T_424 ? reservedFreeList3_55 : reservedFreeList4_55; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1649 = _T_424 ? reservedFreeList3_56 : reservedFreeList4_56; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1650 = _T_424 ? reservedFreeList3_57 : reservedFreeList4_57; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1651 = _T_424 ? reservedFreeList3_58 : reservedFreeList4_58; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1652 = _T_424 ? reservedFreeList3_59 : reservedFreeList4_59; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1653 = _T_424 ? reservedFreeList3_60 : reservedFreeList4_60; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1654 = _T_424 ? reservedFreeList3_61 : reservedFreeList4_61; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1655 = _T_424 ? reservedFreeList3_62 : reservedFreeList4_62; // @[decode.scala 317:30 356:34 377:25]
  wire  _GEN_1657 = _T_424 ? reservedValidList1_0 : reservedValidList2_0; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1658 = _T_424 ? reservedValidList1_1 : reservedValidList2_1; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1659 = _T_424 ? reservedValidList1_2 : reservedValidList2_2; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1660 = _T_424 ? reservedValidList1_3 : reservedValidList2_3; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1661 = _T_424 ? reservedValidList1_4 : reservedValidList2_4; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1662 = _T_424 ? reservedValidList1_5 : reservedValidList2_5; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1663 = _T_424 ? reservedValidList1_6 : reservedValidList2_6; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1664 = _T_424 ? reservedValidList1_7 : reservedValidList2_7; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1665 = _T_424 ? reservedValidList1_8 : reservedValidList2_8; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1666 = _T_424 ? reservedValidList1_9 : reservedValidList2_9; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1667 = _T_424 ? reservedValidList1_10 : reservedValidList2_10; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1668 = _T_424 ? reservedValidList1_11 : reservedValidList2_11; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1669 = _T_424 ? reservedValidList1_12 : reservedValidList2_12; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1670 = _T_424 ? reservedValidList1_13 : reservedValidList2_13; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1671 = _T_424 ? reservedValidList1_14 : reservedValidList2_14; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1672 = _T_424 ? reservedValidList1_15 : reservedValidList2_15; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1673 = _T_424 ? reservedValidList1_16 : reservedValidList2_16; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1674 = _T_424 ? reservedValidList1_17 : reservedValidList2_17; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1675 = _T_424 ? reservedValidList1_18 : reservedValidList2_18; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1676 = _T_424 ? reservedValidList1_19 : reservedValidList2_19; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1677 = _T_424 ? reservedValidList1_20 : reservedValidList2_20; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1678 = _T_424 ? reservedValidList1_21 : reservedValidList2_21; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1679 = _T_424 ? reservedValidList1_22 : reservedValidList2_22; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1680 = _T_424 ? reservedValidList1_23 : reservedValidList2_23; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1681 = _T_424 ? reservedValidList1_24 : reservedValidList2_24; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1682 = _T_424 ? reservedValidList1_25 : reservedValidList2_25; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1683 = _T_424 ? reservedValidList1_26 : reservedValidList2_26; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1684 = _T_424 ? reservedValidList1_27 : reservedValidList2_27; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1685 = _T_424 ? reservedValidList1_28 : reservedValidList2_28; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1686 = _T_424 ? reservedValidList1_29 : reservedValidList2_29; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1687 = _T_424 ? reservedValidList1_30 : reservedValidList2_30; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1688 = _T_424 ? reservedValidList1_31 : reservedValidList2_31; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1689 = _T_424 ? reservedValidList1_32 : reservedValidList2_32; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1690 = _T_424 ? reservedValidList1_33 : reservedValidList2_33; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1691 = _T_424 ? reservedValidList1_34 : reservedValidList2_34; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1692 = _T_424 ? reservedValidList1_35 : reservedValidList2_35; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1693 = _T_424 ? reservedValidList1_36 : reservedValidList2_36; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1694 = _T_424 ? reservedValidList1_37 : reservedValidList2_37; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1695 = _T_424 ? reservedValidList1_38 : reservedValidList2_38; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1696 = _T_424 ? reservedValidList1_39 : reservedValidList2_39; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1697 = _T_424 ? reservedValidList1_40 : reservedValidList2_40; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1698 = _T_424 ? reservedValidList1_41 : reservedValidList2_41; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1699 = _T_424 ? reservedValidList1_42 : reservedValidList2_42; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1700 = _T_424 ? reservedValidList1_43 : reservedValidList2_43; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1701 = _T_424 ? reservedValidList1_44 : reservedValidList2_44; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1702 = _T_424 ? reservedValidList1_45 : reservedValidList2_45; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1703 = _T_424 ? reservedValidList1_46 : reservedValidList2_46; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1704 = _T_424 ? reservedValidList1_47 : reservedValidList2_47; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1705 = _T_424 ? reservedValidList1_48 : reservedValidList2_48; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1706 = _T_424 ? reservedValidList1_49 : reservedValidList2_49; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1707 = _T_424 ? reservedValidList1_50 : reservedValidList2_50; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1708 = _T_424 ? reservedValidList1_51 : reservedValidList2_51; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1709 = _T_424 ? reservedValidList1_52 : reservedValidList2_52; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1710 = _T_424 ? reservedValidList1_53 : reservedValidList2_53; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1711 = _T_424 ? reservedValidList1_54 : reservedValidList2_54; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1712 = _T_424 ? reservedValidList1_55 : reservedValidList2_55; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1713 = _T_424 ? reservedValidList1_56 : reservedValidList2_56; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1714 = _T_424 ? reservedValidList1_57 : reservedValidList2_57; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1715 = _T_424 ? reservedValidList1_58 : reservedValidList2_58; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1716 = _T_424 ? reservedValidList1_59 : reservedValidList2_59; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1717 = _T_424 ? reservedValidList1_60 : reservedValidList2_60; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1718 = _T_424 ? reservedValidList1_61 : reservedValidList2_61; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1719 = _T_424 ? reservedValidList1_62 : reservedValidList2_62; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1720 = _T_424 ? reservedValidList1_63 : reservedValidList2_63; // @[decode.scala 320:31 356:34 379:26]
  wire  _GEN_1721 = _T_424 ? reservedValidList2_0 : reservedValidList3_0; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1722 = _T_424 ? reservedValidList2_1 : reservedValidList3_1; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1723 = _T_424 ? reservedValidList2_2 : reservedValidList3_2; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1724 = _T_424 ? reservedValidList2_3 : reservedValidList3_3; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1725 = _T_424 ? reservedValidList2_4 : reservedValidList3_4; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1726 = _T_424 ? reservedValidList2_5 : reservedValidList3_5; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1727 = _T_424 ? reservedValidList2_6 : reservedValidList3_6; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1728 = _T_424 ? reservedValidList2_7 : reservedValidList3_7; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1729 = _T_424 ? reservedValidList2_8 : reservedValidList3_8; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1730 = _T_424 ? reservedValidList2_9 : reservedValidList3_9; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1731 = _T_424 ? reservedValidList2_10 : reservedValidList3_10; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1732 = _T_424 ? reservedValidList2_11 : reservedValidList3_11; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1733 = _T_424 ? reservedValidList2_12 : reservedValidList3_12; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1734 = _T_424 ? reservedValidList2_13 : reservedValidList3_13; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1735 = _T_424 ? reservedValidList2_14 : reservedValidList3_14; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1736 = _T_424 ? reservedValidList2_15 : reservedValidList3_15; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1737 = _T_424 ? reservedValidList2_16 : reservedValidList3_16; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1738 = _T_424 ? reservedValidList2_17 : reservedValidList3_17; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1739 = _T_424 ? reservedValidList2_18 : reservedValidList3_18; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1740 = _T_424 ? reservedValidList2_19 : reservedValidList3_19; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1741 = _T_424 ? reservedValidList2_20 : reservedValidList3_20; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1742 = _T_424 ? reservedValidList2_21 : reservedValidList3_21; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1743 = _T_424 ? reservedValidList2_22 : reservedValidList3_22; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1744 = _T_424 ? reservedValidList2_23 : reservedValidList3_23; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1745 = _T_424 ? reservedValidList2_24 : reservedValidList3_24; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1746 = _T_424 ? reservedValidList2_25 : reservedValidList3_25; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1747 = _T_424 ? reservedValidList2_26 : reservedValidList3_26; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1748 = _T_424 ? reservedValidList2_27 : reservedValidList3_27; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1749 = _T_424 ? reservedValidList2_28 : reservedValidList3_28; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1750 = _T_424 ? reservedValidList2_29 : reservedValidList3_29; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1751 = _T_424 ? reservedValidList2_30 : reservedValidList3_30; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1752 = _T_424 ? reservedValidList2_31 : reservedValidList3_31; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1753 = _T_424 ? reservedValidList2_32 : reservedValidList3_32; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1754 = _T_424 ? reservedValidList2_33 : reservedValidList3_33; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1755 = _T_424 ? reservedValidList2_34 : reservedValidList3_34; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1756 = _T_424 ? reservedValidList2_35 : reservedValidList3_35; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1757 = _T_424 ? reservedValidList2_36 : reservedValidList3_36; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1758 = _T_424 ? reservedValidList2_37 : reservedValidList3_37; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1759 = _T_424 ? reservedValidList2_38 : reservedValidList3_38; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1760 = _T_424 ? reservedValidList2_39 : reservedValidList3_39; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1761 = _T_424 ? reservedValidList2_40 : reservedValidList3_40; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1762 = _T_424 ? reservedValidList2_41 : reservedValidList3_41; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1763 = _T_424 ? reservedValidList2_42 : reservedValidList3_42; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1764 = _T_424 ? reservedValidList2_43 : reservedValidList3_43; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1765 = _T_424 ? reservedValidList2_44 : reservedValidList3_44; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1766 = _T_424 ? reservedValidList2_45 : reservedValidList3_45; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1767 = _T_424 ? reservedValidList2_46 : reservedValidList3_46; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1768 = _T_424 ? reservedValidList2_47 : reservedValidList3_47; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1769 = _T_424 ? reservedValidList2_48 : reservedValidList3_48; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1770 = _T_424 ? reservedValidList2_49 : reservedValidList3_49; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1771 = _T_424 ? reservedValidList2_50 : reservedValidList3_50; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1772 = _T_424 ? reservedValidList2_51 : reservedValidList3_51; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1773 = _T_424 ? reservedValidList2_52 : reservedValidList3_52; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1774 = _T_424 ? reservedValidList2_53 : reservedValidList3_53; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1775 = _T_424 ? reservedValidList2_54 : reservedValidList3_54; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1776 = _T_424 ? reservedValidList2_55 : reservedValidList3_55; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1777 = _T_424 ? reservedValidList2_56 : reservedValidList3_56; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1778 = _T_424 ? reservedValidList2_57 : reservedValidList3_57; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1779 = _T_424 ? reservedValidList2_58 : reservedValidList3_58; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1780 = _T_424 ? reservedValidList2_59 : reservedValidList3_59; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1781 = _T_424 ? reservedValidList2_60 : reservedValidList3_60; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1782 = _T_424 ? reservedValidList2_61 : reservedValidList3_61; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1783 = _T_424 ? reservedValidList2_62 : reservedValidList3_62; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1784 = _T_424 ? reservedValidList2_63 : reservedValidList3_63; // @[decode.scala 321:31 356:34 380:26]
  wire  _GEN_1785 = _T_424 ? reservedValidList3_0 : reservedValidList4_0; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1786 = _T_424 ? reservedValidList3_1 : reservedValidList4_1; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1787 = _T_424 ? reservedValidList3_2 : reservedValidList4_2; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1788 = _T_424 ? reservedValidList3_3 : reservedValidList4_3; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1789 = _T_424 ? reservedValidList3_4 : reservedValidList4_4; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1790 = _T_424 ? reservedValidList3_5 : reservedValidList4_5; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1791 = _T_424 ? reservedValidList3_6 : reservedValidList4_6; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1792 = _T_424 ? reservedValidList3_7 : reservedValidList4_7; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1793 = _T_424 ? reservedValidList3_8 : reservedValidList4_8; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1794 = _T_424 ? reservedValidList3_9 : reservedValidList4_9; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1795 = _T_424 ? reservedValidList3_10 : reservedValidList4_10; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1796 = _T_424 ? reservedValidList3_11 : reservedValidList4_11; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1797 = _T_424 ? reservedValidList3_12 : reservedValidList4_12; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1798 = _T_424 ? reservedValidList3_13 : reservedValidList4_13; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1799 = _T_424 ? reservedValidList3_14 : reservedValidList4_14; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1800 = _T_424 ? reservedValidList3_15 : reservedValidList4_15; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1801 = _T_424 ? reservedValidList3_16 : reservedValidList4_16; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1802 = _T_424 ? reservedValidList3_17 : reservedValidList4_17; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1803 = _T_424 ? reservedValidList3_18 : reservedValidList4_18; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1804 = _T_424 ? reservedValidList3_19 : reservedValidList4_19; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1805 = _T_424 ? reservedValidList3_20 : reservedValidList4_20; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1806 = _T_424 ? reservedValidList3_21 : reservedValidList4_21; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1807 = _T_424 ? reservedValidList3_22 : reservedValidList4_22; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1808 = _T_424 ? reservedValidList3_23 : reservedValidList4_23; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1809 = _T_424 ? reservedValidList3_24 : reservedValidList4_24; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1810 = _T_424 ? reservedValidList3_25 : reservedValidList4_25; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1811 = _T_424 ? reservedValidList3_26 : reservedValidList4_26; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1812 = _T_424 ? reservedValidList3_27 : reservedValidList4_27; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1813 = _T_424 ? reservedValidList3_28 : reservedValidList4_28; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1814 = _T_424 ? reservedValidList3_29 : reservedValidList4_29; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1815 = _T_424 ? reservedValidList3_30 : reservedValidList4_30; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1816 = _T_424 ? reservedValidList3_31 : reservedValidList4_31; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1817 = _T_424 ? reservedValidList3_32 : reservedValidList4_32; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1818 = _T_424 ? reservedValidList3_33 : reservedValidList4_33; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1819 = _T_424 ? reservedValidList3_34 : reservedValidList4_34; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1820 = _T_424 ? reservedValidList3_35 : reservedValidList4_35; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1821 = _T_424 ? reservedValidList3_36 : reservedValidList4_36; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1822 = _T_424 ? reservedValidList3_37 : reservedValidList4_37; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1823 = _T_424 ? reservedValidList3_38 : reservedValidList4_38; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1824 = _T_424 ? reservedValidList3_39 : reservedValidList4_39; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1825 = _T_424 ? reservedValidList3_40 : reservedValidList4_40; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1826 = _T_424 ? reservedValidList3_41 : reservedValidList4_41; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1827 = _T_424 ? reservedValidList3_42 : reservedValidList4_42; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1828 = _T_424 ? reservedValidList3_43 : reservedValidList4_43; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1829 = _T_424 ? reservedValidList3_44 : reservedValidList4_44; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1830 = _T_424 ? reservedValidList3_45 : reservedValidList4_45; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1831 = _T_424 ? reservedValidList3_46 : reservedValidList4_46; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1832 = _T_424 ? reservedValidList3_47 : reservedValidList4_47; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1833 = _T_424 ? reservedValidList3_48 : reservedValidList4_48; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1834 = _T_424 ? reservedValidList3_49 : reservedValidList4_49; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1835 = _T_424 ? reservedValidList3_50 : reservedValidList4_50; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1836 = _T_424 ? reservedValidList3_51 : reservedValidList4_51; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1837 = _T_424 ? reservedValidList3_52 : reservedValidList4_52; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1838 = _T_424 ? reservedValidList3_53 : reservedValidList4_53; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1839 = _T_424 ? reservedValidList3_54 : reservedValidList4_54; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1840 = _T_424 ? reservedValidList3_55 : reservedValidList4_55; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1841 = _T_424 ? reservedValidList3_56 : reservedValidList4_56; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1842 = _T_424 ? reservedValidList3_57 : reservedValidList4_57; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1843 = _T_424 ? reservedValidList3_58 : reservedValidList4_58; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1844 = _T_424 ? reservedValidList3_59 : reservedValidList4_59; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1845 = _T_424 ? reservedValidList3_60 : reservedValidList4_60; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1846 = _T_424 ? reservedValidList3_61 : reservedValidList4_61; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1847 = _T_424 ? reservedValidList3_62 : reservedValidList4_62; // @[decode.scala 322:31 356:34 381:26]
  wire  _GEN_1848 = _T_424 ? reservedValidList3_63 : reservedValidList4_63; // @[decode.scala 322:31 356:34 381:26]
  wire [2:0] _GEN_1849 = branchEvalIn_fired ? _GEN_1368 : branchTracker; // @[decode.scala 352:28 173:30]
  wire  _GEN_1850 = branchEvalIn_fired ? _GEN_1203 : branchBuffer_branchMask_0; // @[decode.scala 352:28 138:29]
  wire  _GEN_1851 = branchEvalIn_fired ? _GEN_1204 : branchBuffer_branchMask_1; // @[decode.scala 352:28 138:29]
  wire  _GEN_1852 = branchEvalIn_fired ? _GEN_1205 : branchBuffer_branchMask_2; // @[decode.scala 352:28 138:29]
  wire  _GEN_1853 = branchEvalIn_fired ? _GEN_1206 : branchBuffer_branchMask_3; // @[decode.scala 352:28 138:29]
  wire [63:0] _GEN_1855 = branchEvalIn_fired ? _GEN_1207 : expectedPC; // @[decode.scala 183:27 352:28]
  wire  _GEN_1888 = branchEvalIn_fired ? _GEN_1240 : _GEN_1042; // @[decode.scala 352:28]
  wire  _GEN_1889 = branchEvalIn_fired ? _GEN_1241 : _GEN_1043; // @[decode.scala 352:28]
  wire  _GEN_1890 = branchEvalIn_fired ? _GEN_1242 : _GEN_1044; // @[decode.scala 352:28]
  wire  _GEN_1891 = branchEvalIn_fired ? _GEN_1243 : _GEN_1045; // @[decode.scala 352:28]
  wire  _GEN_1892 = branchEvalIn_fired ? _GEN_1244 : _GEN_1046; // @[decode.scala 352:28]
  wire  _GEN_1893 = branchEvalIn_fired ? _GEN_1245 : _GEN_1047; // @[decode.scala 352:28]
  wire  _GEN_1894 = branchEvalIn_fired ? _GEN_1246 : _GEN_1048; // @[decode.scala 352:28]
  wire  _GEN_1895 = branchEvalIn_fired ? _GEN_1247 : _GEN_1049; // @[decode.scala 352:28]
  wire  _GEN_1896 = branchEvalIn_fired ? _GEN_1248 : _GEN_1050; // @[decode.scala 352:28]
  wire  _GEN_1897 = branchEvalIn_fired ? _GEN_1249 : _GEN_1051; // @[decode.scala 352:28]
  wire  _GEN_1898 = branchEvalIn_fired ? _GEN_1250 : _GEN_1052; // @[decode.scala 352:28]
  wire  _GEN_1899 = branchEvalIn_fired ? _GEN_1251 : _GEN_1053; // @[decode.scala 352:28]
  wire  _GEN_1900 = branchEvalIn_fired ? _GEN_1252 : _GEN_1054; // @[decode.scala 352:28]
  wire  _GEN_1901 = branchEvalIn_fired ? _GEN_1253 : _GEN_1055; // @[decode.scala 352:28]
  wire  _GEN_1902 = branchEvalIn_fired ? _GEN_1254 : _GEN_1056; // @[decode.scala 352:28]
  wire  _GEN_1903 = branchEvalIn_fired ? _GEN_1255 : _GEN_1057; // @[decode.scala 352:28]
  wire  _GEN_1904 = branchEvalIn_fired ? _GEN_1256 : _GEN_1058; // @[decode.scala 352:28]
  wire  _GEN_1905 = branchEvalIn_fired ? _GEN_1257 : _GEN_1059; // @[decode.scala 352:28]
  wire  _GEN_1906 = branchEvalIn_fired ? _GEN_1258 : _GEN_1060; // @[decode.scala 352:28]
  wire  _GEN_1907 = branchEvalIn_fired ? _GEN_1259 : _GEN_1061; // @[decode.scala 352:28]
  wire  _GEN_1908 = branchEvalIn_fired ? _GEN_1260 : _GEN_1062; // @[decode.scala 352:28]
  wire  _GEN_1909 = branchEvalIn_fired ? _GEN_1261 : _GEN_1063; // @[decode.scala 352:28]
  wire  _GEN_1910 = branchEvalIn_fired ? _GEN_1262 : _GEN_1064; // @[decode.scala 352:28]
  wire  _GEN_1911 = branchEvalIn_fired ? _GEN_1263 : _GEN_1065; // @[decode.scala 352:28]
  wire  _GEN_1912 = branchEvalIn_fired ? _GEN_1264 : _GEN_1066; // @[decode.scala 352:28]
  wire  _GEN_1913 = branchEvalIn_fired ? _GEN_1265 : _GEN_1067; // @[decode.scala 352:28]
  wire  _GEN_1914 = branchEvalIn_fired ? _GEN_1266 : _GEN_1068; // @[decode.scala 352:28]
  wire  _GEN_1915 = branchEvalIn_fired ? _GEN_1267 : _GEN_1069; // @[decode.scala 352:28]
  wire  _GEN_1916 = branchEvalIn_fired ? _GEN_1268 : _GEN_1070; // @[decode.scala 352:28]
  wire  _GEN_1917 = branchEvalIn_fired ? _GEN_1269 : _GEN_1071; // @[decode.scala 352:28]
  wire  _GEN_1918 = branchEvalIn_fired ? _GEN_1270 : _GEN_1072; // @[decode.scala 352:28]
  wire  _GEN_1919 = branchEvalIn_fired ? _GEN_1271 : _GEN_1073; // @[decode.scala 352:28]
  wire  _GEN_1920 = branchEvalIn_fired ? _GEN_1272 : _GEN_1074; // @[decode.scala 352:28]
  wire  _GEN_1921 = branchEvalIn_fired ? _GEN_1273 : _GEN_1075; // @[decode.scala 352:28]
  wire  _GEN_1922 = branchEvalIn_fired ? _GEN_1274 : _GEN_1076; // @[decode.scala 352:28]
  wire  _GEN_1923 = branchEvalIn_fired ? _GEN_1275 : _GEN_1077; // @[decode.scala 352:28]
  wire  _GEN_1924 = branchEvalIn_fired ? _GEN_1276 : _GEN_1078; // @[decode.scala 352:28]
  wire  _GEN_1925 = branchEvalIn_fired ? _GEN_1277 : _GEN_1079; // @[decode.scala 352:28]
  wire  _GEN_1926 = branchEvalIn_fired ? _GEN_1278 : _GEN_1080; // @[decode.scala 352:28]
  wire  _GEN_1927 = branchEvalIn_fired ? _GEN_1279 : _GEN_1081; // @[decode.scala 352:28]
  wire  _GEN_1928 = branchEvalIn_fired ? _GEN_1280 : _GEN_1082; // @[decode.scala 352:28]
  wire  _GEN_1929 = branchEvalIn_fired ? _GEN_1281 : _GEN_1083; // @[decode.scala 352:28]
  wire  _GEN_1930 = branchEvalIn_fired ? _GEN_1282 : _GEN_1084; // @[decode.scala 352:28]
  wire  _GEN_1931 = branchEvalIn_fired ? _GEN_1283 : _GEN_1085; // @[decode.scala 352:28]
  wire  _GEN_1932 = branchEvalIn_fired ? _GEN_1284 : _GEN_1086; // @[decode.scala 352:28]
  wire  _GEN_1933 = branchEvalIn_fired ? _GEN_1285 : _GEN_1087; // @[decode.scala 352:28]
  wire  _GEN_1934 = branchEvalIn_fired ? _GEN_1286 : _GEN_1088; // @[decode.scala 352:28]
  wire  _GEN_1935 = branchEvalIn_fired ? _GEN_1287 : _GEN_1089; // @[decode.scala 352:28]
  wire  _GEN_1936 = branchEvalIn_fired ? _GEN_1288 : _GEN_1090; // @[decode.scala 352:28]
  wire  _GEN_1937 = branchEvalIn_fired ? _GEN_1289 : _GEN_1091; // @[decode.scala 352:28]
  wire  _GEN_1938 = branchEvalIn_fired ? _GEN_1290 : _GEN_1092; // @[decode.scala 352:28]
  wire  _GEN_1939 = branchEvalIn_fired ? _GEN_1291 : _GEN_1093; // @[decode.scala 352:28]
  wire  _GEN_1940 = branchEvalIn_fired ? _GEN_1292 : _GEN_1094; // @[decode.scala 352:28]
  wire  _GEN_1941 = branchEvalIn_fired ? _GEN_1293 : _GEN_1095; // @[decode.scala 352:28]
  wire  _GEN_1942 = branchEvalIn_fired ? _GEN_1294 : _GEN_1096; // @[decode.scala 352:28]
  wire  _GEN_1943 = branchEvalIn_fired ? _GEN_1295 : _GEN_1097; // @[decode.scala 352:28]
  wire  _GEN_1944 = branchEvalIn_fired ? _GEN_1296 : _GEN_1098; // @[decode.scala 352:28]
  wire  _GEN_1945 = branchEvalIn_fired ? _GEN_1297 : _GEN_1099; // @[decode.scala 352:28]
  wire  _GEN_1946 = branchEvalIn_fired ? _GEN_1298 : _GEN_1100; // @[decode.scala 352:28]
  wire  _GEN_1947 = branchEvalIn_fired ? _GEN_1299 : _GEN_1101; // @[decode.scala 352:28]
  wire  _GEN_1948 = branchEvalIn_fired ? _GEN_1300 : _GEN_1102; // @[decode.scala 352:28]
  wire  _GEN_1949 = branchEvalIn_fired ? _GEN_1301 : _GEN_1103; // @[decode.scala 352:28]
  wire  _GEN_1950 = branchEvalIn_fired ? _GEN_1302 : _GEN_1104; // @[decode.scala 352:28]
  wire  _GEN_1952 = branchEvalIn_fired ? _GEN_1304 : _GEN_1106; // @[decode.scala 352:28]
  wire  _GEN_1953 = branchEvalIn_fired ? _GEN_1305 : _GEN_1107; // @[decode.scala 352:28]
  wire  _GEN_1954 = branchEvalIn_fired ? _GEN_1306 : _GEN_1108; // @[decode.scala 352:28]
  wire  _GEN_1955 = branchEvalIn_fired ? _GEN_1307 : _GEN_1109; // @[decode.scala 352:28]
  wire  _GEN_1956 = branchEvalIn_fired ? _GEN_1308 : _GEN_1110; // @[decode.scala 352:28]
  wire  _GEN_1957 = branchEvalIn_fired ? _GEN_1309 : _GEN_1111; // @[decode.scala 352:28]
  wire  _GEN_1958 = branchEvalIn_fired ? _GEN_1310 : _GEN_1112; // @[decode.scala 352:28]
  wire  _GEN_1959 = branchEvalIn_fired ? _GEN_1311 : _GEN_1113; // @[decode.scala 352:28]
  wire  _GEN_1960 = branchEvalIn_fired ? _GEN_1312 : _GEN_1114; // @[decode.scala 352:28]
  wire  _GEN_1961 = branchEvalIn_fired ? _GEN_1313 : _GEN_1115; // @[decode.scala 352:28]
  wire  _GEN_1962 = branchEvalIn_fired ? _GEN_1314 : _GEN_1116; // @[decode.scala 352:28]
  wire  _GEN_1963 = branchEvalIn_fired ? _GEN_1315 : _GEN_1117; // @[decode.scala 352:28]
  wire  _GEN_1964 = branchEvalIn_fired ? _GEN_1316 : _GEN_1118; // @[decode.scala 352:28]
  wire  _GEN_1965 = branchEvalIn_fired ? _GEN_1317 : _GEN_1119; // @[decode.scala 352:28]
  wire  _GEN_1966 = branchEvalIn_fired ? _GEN_1318 : _GEN_1120; // @[decode.scala 352:28]
  wire  _GEN_1967 = branchEvalIn_fired ? _GEN_1319 : _GEN_1121; // @[decode.scala 352:28]
  wire  _GEN_1968 = branchEvalIn_fired ? _GEN_1320 : _GEN_1122; // @[decode.scala 352:28]
  wire  _GEN_1969 = branchEvalIn_fired ? _GEN_1321 : _GEN_1123; // @[decode.scala 352:28]
  wire  _GEN_1970 = branchEvalIn_fired ? _GEN_1322 : _GEN_1124; // @[decode.scala 352:28]
  wire  _GEN_1971 = branchEvalIn_fired ? _GEN_1323 : _GEN_1125; // @[decode.scala 352:28]
  wire  _GEN_1972 = branchEvalIn_fired ? _GEN_1324 : _GEN_1126; // @[decode.scala 352:28]
  wire  _GEN_1973 = branchEvalIn_fired ? _GEN_1325 : _GEN_1127; // @[decode.scala 352:28]
  wire  _GEN_1974 = branchEvalIn_fired ? _GEN_1326 : _GEN_1128; // @[decode.scala 352:28]
  wire  _GEN_1975 = branchEvalIn_fired ? _GEN_1327 : _GEN_1129; // @[decode.scala 352:28]
  wire  _GEN_1976 = branchEvalIn_fired ? _GEN_1328 : _GEN_1130; // @[decode.scala 352:28]
  wire  _GEN_1977 = branchEvalIn_fired ? _GEN_1329 : _GEN_1131; // @[decode.scala 352:28]
  wire  _GEN_1978 = branchEvalIn_fired ? _GEN_1330 : _GEN_1132; // @[decode.scala 352:28]
  wire  _GEN_1979 = branchEvalIn_fired ? _GEN_1331 : _GEN_1133; // @[decode.scala 352:28]
  wire  _GEN_1980 = branchEvalIn_fired ? _GEN_1332 : _GEN_1134; // @[decode.scala 352:28]
  wire  _GEN_1981 = branchEvalIn_fired ? _GEN_1333 : _GEN_1135; // @[decode.scala 352:28]
  wire  _GEN_1982 = branchEvalIn_fired ? _GEN_1334 : _GEN_1136; // @[decode.scala 352:28]
  wire  _GEN_1983 = branchEvalIn_fired ? _GEN_1335 : _GEN_1137; // @[decode.scala 352:28]
  wire  _GEN_1984 = branchEvalIn_fired ? _GEN_1336 : _GEN_1138; // @[decode.scala 352:28]
  wire  _GEN_1985 = branchEvalIn_fired ? _GEN_1337 : _GEN_1139; // @[decode.scala 352:28]
  wire  _GEN_1986 = branchEvalIn_fired ? _GEN_1338 : _GEN_1140; // @[decode.scala 352:28]
  wire  _GEN_1987 = branchEvalIn_fired ? _GEN_1339 : _GEN_1141; // @[decode.scala 352:28]
  wire  _GEN_1988 = branchEvalIn_fired ? _GEN_1340 : _GEN_1142; // @[decode.scala 352:28]
  wire  _GEN_1989 = branchEvalIn_fired ? _GEN_1341 : _GEN_1143; // @[decode.scala 352:28]
  wire  _GEN_1990 = branchEvalIn_fired ? _GEN_1342 : _GEN_1144; // @[decode.scala 352:28]
  wire  _GEN_1991 = branchEvalIn_fired ? _GEN_1343 : _GEN_1145; // @[decode.scala 352:28]
  wire  _GEN_1992 = branchEvalIn_fired ? _GEN_1344 : _GEN_1146; // @[decode.scala 352:28]
  wire  _GEN_1993 = branchEvalIn_fired ? _GEN_1345 : _GEN_1147; // @[decode.scala 352:28]
  wire  _GEN_1994 = branchEvalIn_fired ? _GEN_1346 : _GEN_1148; // @[decode.scala 352:28]
  wire  _GEN_1995 = branchEvalIn_fired ? _GEN_1347 : _GEN_1149; // @[decode.scala 352:28]
  wire  _GEN_1996 = branchEvalIn_fired ? _GEN_1348 : _GEN_1150; // @[decode.scala 352:28]
  wire  _GEN_1997 = branchEvalIn_fired ? _GEN_1349 : _GEN_1151; // @[decode.scala 352:28]
  wire  _GEN_1998 = branchEvalIn_fired ? _GEN_1350 : _GEN_1152; // @[decode.scala 352:28]
  wire  _GEN_1999 = branchEvalIn_fired ? _GEN_1351 : _GEN_1153; // @[decode.scala 352:28]
  wire  _GEN_2000 = branchEvalIn_fired ? _GEN_1352 : _GEN_1154; // @[decode.scala 352:28]
  wire  _GEN_2001 = branchEvalIn_fired ? _GEN_1353 : _GEN_1155; // @[decode.scala 352:28]
  wire  _GEN_2002 = branchEvalIn_fired ? _GEN_1354 : _GEN_1156; // @[decode.scala 352:28]
  wire  _GEN_2003 = branchEvalIn_fired ? _GEN_1355 : _GEN_1157; // @[decode.scala 352:28]
  wire  _GEN_2004 = branchEvalIn_fired ? _GEN_1356 : _GEN_1158; // @[decode.scala 352:28]
  wire  _GEN_2005 = branchEvalIn_fired ? _GEN_1357 : _GEN_1159; // @[decode.scala 352:28]
  wire  _GEN_2006 = branchEvalIn_fired ? _GEN_1358 : _GEN_1160; // @[decode.scala 352:28]
  wire  _GEN_2007 = branchEvalIn_fired ? _GEN_1359 : _GEN_1161; // @[decode.scala 352:28]
  wire  _GEN_2008 = branchEvalIn_fired ? _GEN_1360 : _GEN_1162; // @[decode.scala 352:28]
  wire  _GEN_2009 = branchEvalIn_fired ? _GEN_1361 : _GEN_1163; // @[decode.scala 352:28]
  wire  _GEN_2010 = branchEvalIn_fired ? _GEN_1362 : _GEN_1164; // @[decode.scala 352:28]
  wire  _GEN_2011 = branchEvalIn_fired ? _GEN_1363 : _GEN_1165; // @[decode.scala 352:28]
  wire  _GEN_2012 = branchEvalIn_fired ? _GEN_1364 : _GEN_1166; // @[decode.scala 352:28]
  wire  _GEN_2013 = branchEvalIn_fired ? _GEN_1365 : _GEN_1167; // @[decode.scala 352:28]
  wire  _GEN_2014 = branchEvalIn_fired ? _GEN_1366 : _GEN_1168; // @[decode.scala 352:28]
  wire  _GEN_2015 = branchEvalIn_fired ? _GEN_1367 : _GEN_1169; // @[decode.scala 352:28]
  wire [5:0] _GEN_2016 = branchEvalIn_fired ? _GEN_1369 : reservedRegMap1_0; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2017 = branchEvalIn_fired ? _GEN_1370 : reservedRegMap1_1; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2018 = branchEvalIn_fired ? _GEN_1371 : reservedRegMap1_2; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2019 = branchEvalIn_fired ? _GEN_1372 : reservedRegMap1_3; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2020 = branchEvalIn_fired ? _GEN_1373 : reservedRegMap1_4; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2021 = branchEvalIn_fired ? _GEN_1374 : reservedRegMap1_5; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2022 = branchEvalIn_fired ? _GEN_1375 : reservedRegMap1_6; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2023 = branchEvalIn_fired ? _GEN_1376 : reservedRegMap1_7; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2024 = branchEvalIn_fired ? _GEN_1377 : reservedRegMap1_8; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2025 = branchEvalIn_fired ? _GEN_1378 : reservedRegMap1_9; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2026 = branchEvalIn_fired ? _GEN_1379 : reservedRegMap1_10; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2027 = branchEvalIn_fired ? _GEN_1380 : reservedRegMap1_11; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2028 = branchEvalIn_fired ? _GEN_1381 : reservedRegMap1_12; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2029 = branchEvalIn_fired ? _GEN_1382 : reservedRegMap1_13; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2030 = branchEvalIn_fired ? _GEN_1383 : reservedRegMap1_14; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2031 = branchEvalIn_fired ? _GEN_1384 : reservedRegMap1_15; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2032 = branchEvalIn_fired ? _GEN_1385 : reservedRegMap1_16; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2033 = branchEvalIn_fired ? _GEN_1386 : reservedRegMap1_17; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2034 = branchEvalIn_fired ? _GEN_1387 : reservedRegMap1_18; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2035 = branchEvalIn_fired ? _GEN_1388 : reservedRegMap1_19; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2036 = branchEvalIn_fired ? _GEN_1389 : reservedRegMap1_20; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2037 = branchEvalIn_fired ? _GEN_1390 : reservedRegMap1_21; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2038 = branchEvalIn_fired ? _GEN_1391 : reservedRegMap1_22; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2039 = branchEvalIn_fired ? _GEN_1392 : reservedRegMap1_23; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2040 = branchEvalIn_fired ? _GEN_1393 : reservedRegMap1_24; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2041 = branchEvalIn_fired ? _GEN_1394 : reservedRegMap1_25; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2042 = branchEvalIn_fired ? _GEN_1395 : reservedRegMap1_26; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2043 = branchEvalIn_fired ? _GEN_1396 : reservedRegMap1_27; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2044 = branchEvalIn_fired ? _GEN_1397 : reservedRegMap1_28; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2045 = branchEvalIn_fired ? _GEN_1398 : reservedRegMap1_29; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2046 = branchEvalIn_fired ? _GEN_1399 : reservedRegMap1_30; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2047 = branchEvalIn_fired ? _GEN_1400 : reservedRegMap1_31; // @[decode.scala 310:28 352:28]
  wire [5:0] _GEN_2048 = branchEvalIn_fired ? _GEN_1401 : reservedRegMap2_0; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2049 = branchEvalIn_fired ? _GEN_1402 : reservedRegMap2_1; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2050 = branchEvalIn_fired ? _GEN_1403 : reservedRegMap2_2; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2051 = branchEvalIn_fired ? _GEN_1404 : reservedRegMap2_3; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2052 = branchEvalIn_fired ? _GEN_1405 : reservedRegMap2_4; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2053 = branchEvalIn_fired ? _GEN_1406 : reservedRegMap2_5; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2054 = branchEvalIn_fired ? _GEN_1407 : reservedRegMap2_6; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2055 = branchEvalIn_fired ? _GEN_1408 : reservedRegMap2_7; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2056 = branchEvalIn_fired ? _GEN_1409 : reservedRegMap2_8; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2057 = branchEvalIn_fired ? _GEN_1410 : reservedRegMap2_9; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2058 = branchEvalIn_fired ? _GEN_1411 : reservedRegMap2_10; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2059 = branchEvalIn_fired ? _GEN_1412 : reservedRegMap2_11; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2060 = branchEvalIn_fired ? _GEN_1413 : reservedRegMap2_12; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2061 = branchEvalIn_fired ? _GEN_1414 : reservedRegMap2_13; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2062 = branchEvalIn_fired ? _GEN_1415 : reservedRegMap2_14; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2063 = branchEvalIn_fired ? _GEN_1416 : reservedRegMap2_15; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2064 = branchEvalIn_fired ? _GEN_1417 : reservedRegMap2_16; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2065 = branchEvalIn_fired ? _GEN_1418 : reservedRegMap2_17; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2066 = branchEvalIn_fired ? _GEN_1419 : reservedRegMap2_18; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2067 = branchEvalIn_fired ? _GEN_1420 : reservedRegMap2_19; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2068 = branchEvalIn_fired ? _GEN_1421 : reservedRegMap2_20; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2069 = branchEvalIn_fired ? _GEN_1422 : reservedRegMap2_21; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2070 = branchEvalIn_fired ? _GEN_1423 : reservedRegMap2_22; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2071 = branchEvalIn_fired ? _GEN_1424 : reservedRegMap2_23; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2072 = branchEvalIn_fired ? _GEN_1425 : reservedRegMap2_24; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2073 = branchEvalIn_fired ? _GEN_1426 : reservedRegMap2_25; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2074 = branchEvalIn_fired ? _GEN_1427 : reservedRegMap2_26; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2075 = branchEvalIn_fired ? _GEN_1428 : reservedRegMap2_27; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2076 = branchEvalIn_fired ? _GEN_1429 : reservedRegMap2_28; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2077 = branchEvalIn_fired ? _GEN_1430 : reservedRegMap2_29; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2078 = branchEvalIn_fired ? _GEN_1431 : reservedRegMap2_30; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2079 = branchEvalIn_fired ? _GEN_1432 : reservedRegMap2_31; // @[decode.scala 311:28 352:28]
  wire [5:0] _GEN_2080 = branchEvalIn_fired ? _GEN_1433 : reservedRegMap3_0; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2081 = branchEvalIn_fired ? _GEN_1434 : reservedRegMap3_1; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2082 = branchEvalIn_fired ? _GEN_1435 : reservedRegMap3_2; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2083 = branchEvalIn_fired ? _GEN_1436 : reservedRegMap3_3; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2084 = branchEvalIn_fired ? _GEN_1437 : reservedRegMap3_4; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2085 = branchEvalIn_fired ? _GEN_1438 : reservedRegMap3_5; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2086 = branchEvalIn_fired ? _GEN_1439 : reservedRegMap3_6; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2087 = branchEvalIn_fired ? _GEN_1440 : reservedRegMap3_7; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2088 = branchEvalIn_fired ? _GEN_1441 : reservedRegMap3_8; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2089 = branchEvalIn_fired ? _GEN_1442 : reservedRegMap3_9; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2090 = branchEvalIn_fired ? _GEN_1443 : reservedRegMap3_10; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2091 = branchEvalIn_fired ? _GEN_1444 : reservedRegMap3_11; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2092 = branchEvalIn_fired ? _GEN_1445 : reservedRegMap3_12; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2093 = branchEvalIn_fired ? _GEN_1446 : reservedRegMap3_13; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2094 = branchEvalIn_fired ? _GEN_1447 : reservedRegMap3_14; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2095 = branchEvalIn_fired ? _GEN_1448 : reservedRegMap3_15; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2096 = branchEvalIn_fired ? _GEN_1449 : reservedRegMap3_16; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2097 = branchEvalIn_fired ? _GEN_1450 : reservedRegMap3_17; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2098 = branchEvalIn_fired ? _GEN_1451 : reservedRegMap3_18; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2099 = branchEvalIn_fired ? _GEN_1452 : reservedRegMap3_19; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2100 = branchEvalIn_fired ? _GEN_1453 : reservedRegMap3_20; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2101 = branchEvalIn_fired ? _GEN_1454 : reservedRegMap3_21; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2102 = branchEvalIn_fired ? _GEN_1455 : reservedRegMap3_22; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2103 = branchEvalIn_fired ? _GEN_1456 : reservedRegMap3_23; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2104 = branchEvalIn_fired ? _GEN_1457 : reservedRegMap3_24; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2105 = branchEvalIn_fired ? _GEN_1458 : reservedRegMap3_25; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2106 = branchEvalIn_fired ? _GEN_1459 : reservedRegMap3_26; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2107 = branchEvalIn_fired ? _GEN_1460 : reservedRegMap3_27; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2108 = branchEvalIn_fired ? _GEN_1461 : reservedRegMap3_28; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2109 = branchEvalIn_fired ? _GEN_1462 : reservedRegMap3_29; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2110 = branchEvalIn_fired ? _GEN_1463 : reservedRegMap3_30; // @[decode.scala 312:28 352:28]
  wire [5:0] _GEN_2111 = branchEvalIn_fired ? _GEN_1464 : reservedRegMap3_31; // @[decode.scala 312:28 352:28]
  wire  _GEN_2112 = branchEvalIn_fired ? _GEN_1465 : reservedFreeList1_0; // @[decode.scala 352:28 315:30]
  wire  _GEN_2113 = branchEvalIn_fired ? _GEN_1466 : reservedFreeList1_1; // @[decode.scala 352:28 315:30]
  wire  _GEN_2114 = branchEvalIn_fired ? _GEN_1467 : reservedFreeList1_2; // @[decode.scala 352:28 315:30]
  wire  _GEN_2115 = branchEvalIn_fired ? _GEN_1468 : reservedFreeList1_3; // @[decode.scala 352:28 315:30]
  wire  _GEN_2116 = branchEvalIn_fired ? _GEN_1469 : reservedFreeList1_4; // @[decode.scala 352:28 315:30]
  wire  _GEN_2117 = branchEvalIn_fired ? _GEN_1470 : reservedFreeList1_5; // @[decode.scala 352:28 315:30]
  wire  _GEN_2118 = branchEvalIn_fired ? _GEN_1471 : reservedFreeList1_6; // @[decode.scala 352:28 315:30]
  wire  _GEN_2119 = branchEvalIn_fired ? _GEN_1472 : reservedFreeList1_7; // @[decode.scala 352:28 315:30]
  wire  _GEN_2120 = branchEvalIn_fired ? _GEN_1473 : reservedFreeList1_8; // @[decode.scala 352:28 315:30]
  wire  _GEN_2121 = branchEvalIn_fired ? _GEN_1474 : reservedFreeList1_9; // @[decode.scala 352:28 315:30]
  wire  _GEN_2122 = branchEvalIn_fired ? _GEN_1475 : reservedFreeList1_10; // @[decode.scala 352:28 315:30]
  wire  _GEN_2123 = branchEvalIn_fired ? _GEN_1476 : reservedFreeList1_11; // @[decode.scala 352:28 315:30]
  wire  _GEN_2124 = branchEvalIn_fired ? _GEN_1477 : reservedFreeList1_12; // @[decode.scala 352:28 315:30]
  wire  _GEN_2125 = branchEvalIn_fired ? _GEN_1478 : reservedFreeList1_13; // @[decode.scala 352:28 315:30]
  wire  _GEN_2126 = branchEvalIn_fired ? _GEN_1479 : reservedFreeList1_14; // @[decode.scala 352:28 315:30]
  wire  _GEN_2127 = branchEvalIn_fired ? _GEN_1480 : reservedFreeList1_15; // @[decode.scala 352:28 315:30]
  wire  _GEN_2128 = branchEvalIn_fired ? _GEN_1481 : reservedFreeList1_16; // @[decode.scala 352:28 315:30]
  wire  _GEN_2129 = branchEvalIn_fired ? _GEN_1482 : reservedFreeList1_17; // @[decode.scala 352:28 315:30]
  wire  _GEN_2130 = branchEvalIn_fired ? _GEN_1483 : reservedFreeList1_18; // @[decode.scala 352:28 315:30]
  wire  _GEN_2131 = branchEvalIn_fired ? _GEN_1484 : reservedFreeList1_19; // @[decode.scala 352:28 315:30]
  wire  _GEN_2132 = branchEvalIn_fired ? _GEN_1485 : reservedFreeList1_20; // @[decode.scala 352:28 315:30]
  wire  _GEN_2133 = branchEvalIn_fired ? _GEN_1486 : reservedFreeList1_21; // @[decode.scala 352:28 315:30]
  wire  _GEN_2134 = branchEvalIn_fired ? _GEN_1487 : reservedFreeList1_22; // @[decode.scala 352:28 315:30]
  wire  _GEN_2135 = branchEvalIn_fired ? _GEN_1488 : reservedFreeList1_23; // @[decode.scala 352:28 315:30]
  wire  _GEN_2136 = branchEvalIn_fired ? _GEN_1489 : reservedFreeList1_24; // @[decode.scala 352:28 315:30]
  wire  _GEN_2137 = branchEvalIn_fired ? _GEN_1490 : reservedFreeList1_25; // @[decode.scala 352:28 315:30]
  wire  _GEN_2138 = branchEvalIn_fired ? _GEN_1491 : reservedFreeList1_26; // @[decode.scala 352:28 315:30]
  wire  _GEN_2139 = branchEvalIn_fired ? _GEN_1492 : reservedFreeList1_27; // @[decode.scala 352:28 315:30]
  wire  _GEN_2140 = branchEvalIn_fired ? _GEN_1493 : reservedFreeList1_28; // @[decode.scala 352:28 315:30]
  wire  _GEN_2141 = branchEvalIn_fired ? _GEN_1494 : reservedFreeList1_29; // @[decode.scala 352:28 315:30]
  wire  _GEN_2142 = branchEvalIn_fired ? _GEN_1495 : reservedFreeList1_30; // @[decode.scala 352:28 315:30]
  wire  _GEN_2143 = branchEvalIn_fired ? _GEN_1496 : reservedFreeList1_31; // @[decode.scala 352:28 315:30]
  wire  _GEN_2144 = branchEvalIn_fired ? _GEN_1497 : reservedFreeList1_32; // @[decode.scala 352:28 315:30]
  wire  _GEN_2145 = branchEvalIn_fired ? _GEN_1498 : reservedFreeList1_33; // @[decode.scala 352:28 315:30]
  wire  _GEN_2146 = branchEvalIn_fired ? _GEN_1499 : reservedFreeList1_34; // @[decode.scala 352:28 315:30]
  wire  _GEN_2147 = branchEvalIn_fired ? _GEN_1500 : reservedFreeList1_35; // @[decode.scala 352:28 315:30]
  wire  _GEN_2148 = branchEvalIn_fired ? _GEN_1501 : reservedFreeList1_36; // @[decode.scala 352:28 315:30]
  wire  _GEN_2149 = branchEvalIn_fired ? _GEN_1502 : reservedFreeList1_37; // @[decode.scala 352:28 315:30]
  wire  _GEN_2150 = branchEvalIn_fired ? _GEN_1503 : reservedFreeList1_38; // @[decode.scala 352:28 315:30]
  wire  _GEN_2151 = branchEvalIn_fired ? _GEN_1504 : reservedFreeList1_39; // @[decode.scala 352:28 315:30]
  wire  _GEN_2152 = branchEvalIn_fired ? _GEN_1505 : reservedFreeList1_40; // @[decode.scala 352:28 315:30]
  wire  _GEN_2153 = branchEvalIn_fired ? _GEN_1506 : reservedFreeList1_41; // @[decode.scala 352:28 315:30]
  wire  _GEN_2154 = branchEvalIn_fired ? _GEN_1507 : reservedFreeList1_42; // @[decode.scala 352:28 315:30]
  wire  _GEN_2155 = branchEvalIn_fired ? _GEN_1508 : reservedFreeList1_43; // @[decode.scala 352:28 315:30]
  wire  _GEN_2156 = branchEvalIn_fired ? _GEN_1509 : reservedFreeList1_44; // @[decode.scala 352:28 315:30]
  wire  _GEN_2157 = branchEvalIn_fired ? _GEN_1510 : reservedFreeList1_45; // @[decode.scala 352:28 315:30]
  wire  _GEN_2158 = branchEvalIn_fired ? _GEN_1511 : reservedFreeList1_46; // @[decode.scala 352:28 315:30]
  wire  _GEN_2159 = branchEvalIn_fired ? _GEN_1512 : reservedFreeList1_47; // @[decode.scala 352:28 315:30]
  wire  _GEN_2160 = branchEvalIn_fired ? _GEN_1513 : reservedFreeList1_48; // @[decode.scala 352:28 315:30]
  wire  _GEN_2161 = branchEvalIn_fired ? _GEN_1514 : reservedFreeList1_49; // @[decode.scala 352:28 315:30]
  wire  _GEN_2162 = branchEvalIn_fired ? _GEN_1515 : reservedFreeList1_50; // @[decode.scala 352:28 315:30]
  wire  _GEN_2163 = branchEvalIn_fired ? _GEN_1516 : reservedFreeList1_51; // @[decode.scala 352:28 315:30]
  wire  _GEN_2164 = branchEvalIn_fired ? _GEN_1517 : reservedFreeList1_52; // @[decode.scala 352:28 315:30]
  wire  _GEN_2165 = branchEvalIn_fired ? _GEN_1518 : reservedFreeList1_53; // @[decode.scala 352:28 315:30]
  wire  _GEN_2166 = branchEvalIn_fired ? _GEN_1519 : reservedFreeList1_54; // @[decode.scala 352:28 315:30]
  wire  _GEN_2167 = branchEvalIn_fired ? _GEN_1520 : reservedFreeList1_55; // @[decode.scala 352:28 315:30]
  wire  _GEN_2168 = branchEvalIn_fired ? _GEN_1521 : reservedFreeList1_56; // @[decode.scala 352:28 315:30]
  wire  _GEN_2169 = branchEvalIn_fired ? _GEN_1522 : reservedFreeList1_57; // @[decode.scala 352:28 315:30]
  wire  _GEN_2170 = branchEvalIn_fired ? _GEN_1523 : reservedFreeList1_58; // @[decode.scala 352:28 315:30]
  wire  _GEN_2171 = branchEvalIn_fired ? _GEN_1524 : reservedFreeList1_59; // @[decode.scala 352:28 315:30]
  wire  _GEN_2172 = branchEvalIn_fired ? _GEN_1525 : reservedFreeList1_60; // @[decode.scala 352:28 315:30]
  wire  _GEN_2173 = branchEvalIn_fired ? _GEN_1526 : reservedFreeList1_61; // @[decode.scala 352:28 315:30]
  wire  _GEN_2174 = branchEvalIn_fired ? _GEN_1527 : reservedFreeList1_62; // @[decode.scala 352:28 315:30]
  wire  _GEN_2176 = branchEvalIn_fired ? _GEN_1529 : reservedFreeList2_0; // @[decode.scala 352:28 316:30]
  wire  _GEN_2177 = branchEvalIn_fired ? _GEN_1530 : reservedFreeList2_1; // @[decode.scala 352:28 316:30]
  wire  _GEN_2178 = branchEvalIn_fired ? _GEN_1531 : reservedFreeList2_2; // @[decode.scala 352:28 316:30]
  wire  _GEN_2179 = branchEvalIn_fired ? _GEN_1532 : reservedFreeList2_3; // @[decode.scala 352:28 316:30]
  wire  _GEN_2180 = branchEvalIn_fired ? _GEN_1533 : reservedFreeList2_4; // @[decode.scala 352:28 316:30]
  wire  _GEN_2181 = branchEvalIn_fired ? _GEN_1534 : reservedFreeList2_5; // @[decode.scala 352:28 316:30]
  wire  _GEN_2182 = branchEvalIn_fired ? _GEN_1535 : reservedFreeList2_6; // @[decode.scala 352:28 316:30]
  wire  _GEN_2183 = branchEvalIn_fired ? _GEN_1536 : reservedFreeList2_7; // @[decode.scala 352:28 316:30]
  wire  _GEN_2184 = branchEvalIn_fired ? _GEN_1537 : reservedFreeList2_8; // @[decode.scala 352:28 316:30]
  wire  _GEN_2185 = branchEvalIn_fired ? _GEN_1538 : reservedFreeList2_9; // @[decode.scala 352:28 316:30]
  wire  _GEN_2186 = branchEvalIn_fired ? _GEN_1539 : reservedFreeList2_10; // @[decode.scala 352:28 316:30]
  wire  _GEN_2187 = branchEvalIn_fired ? _GEN_1540 : reservedFreeList2_11; // @[decode.scala 352:28 316:30]
  wire  _GEN_2188 = branchEvalIn_fired ? _GEN_1541 : reservedFreeList2_12; // @[decode.scala 352:28 316:30]
  wire  _GEN_2189 = branchEvalIn_fired ? _GEN_1542 : reservedFreeList2_13; // @[decode.scala 352:28 316:30]
  wire  _GEN_2190 = branchEvalIn_fired ? _GEN_1543 : reservedFreeList2_14; // @[decode.scala 352:28 316:30]
  wire  _GEN_2191 = branchEvalIn_fired ? _GEN_1544 : reservedFreeList2_15; // @[decode.scala 352:28 316:30]
  wire  _GEN_2192 = branchEvalIn_fired ? _GEN_1545 : reservedFreeList2_16; // @[decode.scala 352:28 316:30]
  wire  _GEN_2193 = branchEvalIn_fired ? _GEN_1546 : reservedFreeList2_17; // @[decode.scala 352:28 316:30]
  wire  _GEN_2194 = branchEvalIn_fired ? _GEN_1547 : reservedFreeList2_18; // @[decode.scala 352:28 316:30]
  wire  _GEN_2195 = branchEvalIn_fired ? _GEN_1548 : reservedFreeList2_19; // @[decode.scala 352:28 316:30]
  wire  _GEN_2196 = branchEvalIn_fired ? _GEN_1549 : reservedFreeList2_20; // @[decode.scala 352:28 316:30]
  wire  _GEN_2197 = branchEvalIn_fired ? _GEN_1550 : reservedFreeList2_21; // @[decode.scala 352:28 316:30]
  wire  _GEN_2198 = branchEvalIn_fired ? _GEN_1551 : reservedFreeList2_22; // @[decode.scala 352:28 316:30]
  wire  _GEN_2199 = branchEvalIn_fired ? _GEN_1552 : reservedFreeList2_23; // @[decode.scala 352:28 316:30]
  wire  _GEN_2200 = branchEvalIn_fired ? _GEN_1553 : reservedFreeList2_24; // @[decode.scala 352:28 316:30]
  wire  _GEN_2201 = branchEvalIn_fired ? _GEN_1554 : reservedFreeList2_25; // @[decode.scala 352:28 316:30]
  wire  _GEN_2202 = branchEvalIn_fired ? _GEN_1555 : reservedFreeList2_26; // @[decode.scala 352:28 316:30]
  wire  _GEN_2203 = branchEvalIn_fired ? _GEN_1556 : reservedFreeList2_27; // @[decode.scala 352:28 316:30]
  wire  _GEN_2204 = branchEvalIn_fired ? _GEN_1557 : reservedFreeList2_28; // @[decode.scala 352:28 316:30]
  wire  _GEN_2205 = branchEvalIn_fired ? _GEN_1558 : reservedFreeList2_29; // @[decode.scala 352:28 316:30]
  wire  _GEN_2206 = branchEvalIn_fired ? _GEN_1559 : reservedFreeList2_30; // @[decode.scala 352:28 316:30]
  wire  _GEN_2207 = branchEvalIn_fired ? _GEN_1560 : reservedFreeList2_31; // @[decode.scala 352:28 316:30]
  wire  _GEN_2208 = branchEvalIn_fired ? _GEN_1561 : reservedFreeList2_32; // @[decode.scala 352:28 316:30]
  wire  _GEN_2209 = branchEvalIn_fired ? _GEN_1562 : reservedFreeList2_33; // @[decode.scala 352:28 316:30]
  wire  _GEN_2210 = branchEvalIn_fired ? _GEN_1563 : reservedFreeList2_34; // @[decode.scala 352:28 316:30]
  wire  _GEN_2211 = branchEvalIn_fired ? _GEN_1564 : reservedFreeList2_35; // @[decode.scala 352:28 316:30]
  wire  _GEN_2212 = branchEvalIn_fired ? _GEN_1565 : reservedFreeList2_36; // @[decode.scala 352:28 316:30]
  wire  _GEN_2213 = branchEvalIn_fired ? _GEN_1566 : reservedFreeList2_37; // @[decode.scala 352:28 316:30]
  wire  _GEN_2214 = branchEvalIn_fired ? _GEN_1567 : reservedFreeList2_38; // @[decode.scala 352:28 316:30]
  wire  _GEN_2215 = branchEvalIn_fired ? _GEN_1568 : reservedFreeList2_39; // @[decode.scala 352:28 316:30]
  wire  _GEN_2216 = branchEvalIn_fired ? _GEN_1569 : reservedFreeList2_40; // @[decode.scala 352:28 316:30]
  wire  _GEN_2217 = branchEvalIn_fired ? _GEN_1570 : reservedFreeList2_41; // @[decode.scala 352:28 316:30]
  wire  _GEN_2218 = branchEvalIn_fired ? _GEN_1571 : reservedFreeList2_42; // @[decode.scala 352:28 316:30]
  wire  _GEN_2219 = branchEvalIn_fired ? _GEN_1572 : reservedFreeList2_43; // @[decode.scala 352:28 316:30]
  wire  _GEN_2220 = branchEvalIn_fired ? _GEN_1573 : reservedFreeList2_44; // @[decode.scala 352:28 316:30]
  wire  _GEN_2221 = branchEvalIn_fired ? _GEN_1574 : reservedFreeList2_45; // @[decode.scala 352:28 316:30]
  wire  _GEN_2222 = branchEvalIn_fired ? _GEN_1575 : reservedFreeList2_46; // @[decode.scala 352:28 316:30]
  wire  _GEN_2223 = branchEvalIn_fired ? _GEN_1576 : reservedFreeList2_47; // @[decode.scala 352:28 316:30]
  wire  _GEN_2224 = branchEvalIn_fired ? _GEN_1577 : reservedFreeList2_48; // @[decode.scala 352:28 316:30]
  wire  _GEN_2225 = branchEvalIn_fired ? _GEN_1578 : reservedFreeList2_49; // @[decode.scala 352:28 316:30]
  wire  _GEN_2226 = branchEvalIn_fired ? _GEN_1579 : reservedFreeList2_50; // @[decode.scala 352:28 316:30]
  wire  _GEN_2227 = branchEvalIn_fired ? _GEN_1580 : reservedFreeList2_51; // @[decode.scala 352:28 316:30]
  wire  _GEN_2228 = branchEvalIn_fired ? _GEN_1581 : reservedFreeList2_52; // @[decode.scala 352:28 316:30]
  wire  _GEN_2229 = branchEvalIn_fired ? _GEN_1582 : reservedFreeList2_53; // @[decode.scala 352:28 316:30]
  wire  _GEN_2230 = branchEvalIn_fired ? _GEN_1583 : reservedFreeList2_54; // @[decode.scala 352:28 316:30]
  wire  _GEN_2231 = branchEvalIn_fired ? _GEN_1584 : reservedFreeList2_55; // @[decode.scala 352:28 316:30]
  wire  _GEN_2232 = branchEvalIn_fired ? _GEN_1585 : reservedFreeList2_56; // @[decode.scala 352:28 316:30]
  wire  _GEN_2233 = branchEvalIn_fired ? _GEN_1586 : reservedFreeList2_57; // @[decode.scala 352:28 316:30]
  wire  _GEN_2234 = branchEvalIn_fired ? _GEN_1587 : reservedFreeList2_58; // @[decode.scala 352:28 316:30]
  wire  _GEN_2235 = branchEvalIn_fired ? _GEN_1588 : reservedFreeList2_59; // @[decode.scala 352:28 316:30]
  wire  _GEN_2236 = branchEvalIn_fired ? _GEN_1589 : reservedFreeList2_60; // @[decode.scala 352:28 316:30]
  wire  _GEN_2237 = branchEvalIn_fired ? _GEN_1590 : reservedFreeList2_61; // @[decode.scala 352:28 316:30]
  wire  _GEN_2238 = branchEvalIn_fired ? _GEN_1591 : reservedFreeList2_62; // @[decode.scala 352:28 316:30]
  wire  _GEN_2240 = branchEvalIn_fired ? _GEN_1593 : reservedFreeList3_0; // @[decode.scala 352:28 317:30]
  wire  _GEN_2241 = branchEvalIn_fired ? _GEN_1594 : reservedFreeList3_1; // @[decode.scala 352:28 317:30]
  wire  _GEN_2242 = branchEvalIn_fired ? _GEN_1595 : reservedFreeList3_2; // @[decode.scala 352:28 317:30]
  wire  _GEN_2243 = branchEvalIn_fired ? _GEN_1596 : reservedFreeList3_3; // @[decode.scala 352:28 317:30]
  wire  _GEN_2244 = branchEvalIn_fired ? _GEN_1597 : reservedFreeList3_4; // @[decode.scala 352:28 317:30]
  wire  _GEN_2245 = branchEvalIn_fired ? _GEN_1598 : reservedFreeList3_5; // @[decode.scala 352:28 317:30]
  wire  _GEN_2246 = branchEvalIn_fired ? _GEN_1599 : reservedFreeList3_6; // @[decode.scala 352:28 317:30]
  wire  _GEN_2247 = branchEvalIn_fired ? _GEN_1600 : reservedFreeList3_7; // @[decode.scala 352:28 317:30]
  wire  _GEN_2248 = branchEvalIn_fired ? _GEN_1601 : reservedFreeList3_8; // @[decode.scala 352:28 317:30]
  wire  _GEN_2249 = branchEvalIn_fired ? _GEN_1602 : reservedFreeList3_9; // @[decode.scala 352:28 317:30]
  wire  _GEN_2250 = branchEvalIn_fired ? _GEN_1603 : reservedFreeList3_10; // @[decode.scala 352:28 317:30]
  wire  _GEN_2251 = branchEvalIn_fired ? _GEN_1604 : reservedFreeList3_11; // @[decode.scala 352:28 317:30]
  wire  _GEN_2252 = branchEvalIn_fired ? _GEN_1605 : reservedFreeList3_12; // @[decode.scala 352:28 317:30]
  wire  _GEN_2253 = branchEvalIn_fired ? _GEN_1606 : reservedFreeList3_13; // @[decode.scala 352:28 317:30]
  wire  _GEN_2254 = branchEvalIn_fired ? _GEN_1607 : reservedFreeList3_14; // @[decode.scala 352:28 317:30]
  wire  _GEN_2255 = branchEvalIn_fired ? _GEN_1608 : reservedFreeList3_15; // @[decode.scala 352:28 317:30]
  wire  _GEN_2256 = branchEvalIn_fired ? _GEN_1609 : reservedFreeList3_16; // @[decode.scala 352:28 317:30]
  wire  _GEN_2257 = branchEvalIn_fired ? _GEN_1610 : reservedFreeList3_17; // @[decode.scala 352:28 317:30]
  wire  _GEN_2258 = branchEvalIn_fired ? _GEN_1611 : reservedFreeList3_18; // @[decode.scala 352:28 317:30]
  wire  _GEN_2259 = branchEvalIn_fired ? _GEN_1612 : reservedFreeList3_19; // @[decode.scala 352:28 317:30]
  wire  _GEN_2260 = branchEvalIn_fired ? _GEN_1613 : reservedFreeList3_20; // @[decode.scala 352:28 317:30]
  wire  _GEN_2261 = branchEvalIn_fired ? _GEN_1614 : reservedFreeList3_21; // @[decode.scala 352:28 317:30]
  wire  _GEN_2262 = branchEvalIn_fired ? _GEN_1615 : reservedFreeList3_22; // @[decode.scala 352:28 317:30]
  wire  _GEN_2263 = branchEvalIn_fired ? _GEN_1616 : reservedFreeList3_23; // @[decode.scala 352:28 317:30]
  wire  _GEN_2264 = branchEvalIn_fired ? _GEN_1617 : reservedFreeList3_24; // @[decode.scala 352:28 317:30]
  wire  _GEN_2265 = branchEvalIn_fired ? _GEN_1618 : reservedFreeList3_25; // @[decode.scala 352:28 317:30]
  wire  _GEN_2266 = branchEvalIn_fired ? _GEN_1619 : reservedFreeList3_26; // @[decode.scala 352:28 317:30]
  wire  _GEN_2267 = branchEvalIn_fired ? _GEN_1620 : reservedFreeList3_27; // @[decode.scala 352:28 317:30]
  wire  _GEN_2268 = branchEvalIn_fired ? _GEN_1621 : reservedFreeList3_28; // @[decode.scala 352:28 317:30]
  wire  _GEN_2269 = branchEvalIn_fired ? _GEN_1622 : reservedFreeList3_29; // @[decode.scala 352:28 317:30]
  wire  _GEN_2270 = branchEvalIn_fired ? _GEN_1623 : reservedFreeList3_30; // @[decode.scala 352:28 317:30]
  wire  _GEN_2271 = branchEvalIn_fired ? _GEN_1624 : reservedFreeList3_31; // @[decode.scala 352:28 317:30]
  wire  _GEN_2272 = branchEvalIn_fired ? _GEN_1625 : reservedFreeList3_32; // @[decode.scala 352:28 317:30]
  wire  _GEN_2273 = branchEvalIn_fired ? _GEN_1626 : reservedFreeList3_33; // @[decode.scala 352:28 317:30]
  wire  _GEN_2274 = branchEvalIn_fired ? _GEN_1627 : reservedFreeList3_34; // @[decode.scala 352:28 317:30]
  wire  _GEN_2275 = branchEvalIn_fired ? _GEN_1628 : reservedFreeList3_35; // @[decode.scala 352:28 317:30]
  wire  _GEN_2276 = branchEvalIn_fired ? _GEN_1629 : reservedFreeList3_36; // @[decode.scala 352:28 317:30]
  wire  _GEN_2277 = branchEvalIn_fired ? _GEN_1630 : reservedFreeList3_37; // @[decode.scala 352:28 317:30]
  wire  _GEN_2278 = branchEvalIn_fired ? _GEN_1631 : reservedFreeList3_38; // @[decode.scala 352:28 317:30]
  wire  _GEN_2279 = branchEvalIn_fired ? _GEN_1632 : reservedFreeList3_39; // @[decode.scala 352:28 317:30]
  wire  _GEN_2280 = branchEvalIn_fired ? _GEN_1633 : reservedFreeList3_40; // @[decode.scala 352:28 317:30]
  wire  _GEN_2281 = branchEvalIn_fired ? _GEN_1634 : reservedFreeList3_41; // @[decode.scala 352:28 317:30]
  wire  _GEN_2282 = branchEvalIn_fired ? _GEN_1635 : reservedFreeList3_42; // @[decode.scala 352:28 317:30]
  wire  _GEN_2283 = branchEvalIn_fired ? _GEN_1636 : reservedFreeList3_43; // @[decode.scala 352:28 317:30]
  wire  _GEN_2284 = branchEvalIn_fired ? _GEN_1637 : reservedFreeList3_44; // @[decode.scala 352:28 317:30]
  wire  _GEN_2285 = branchEvalIn_fired ? _GEN_1638 : reservedFreeList3_45; // @[decode.scala 352:28 317:30]
  wire  _GEN_2286 = branchEvalIn_fired ? _GEN_1639 : reservedFreeList3_46; // @[decode.scala 352:28 317:30]
  wire  _GEN_2287 = branchEvalIn_fired ? _GEN_1640 : reservedFreeList3_47; // @[decode.scala 352:28 317:30]
  wire  _GEN_2288 = branchEvalIn_fired ? _GEN_1641 : reservedFreeList3_48; // @[decode.scala 352:28 317:30]
  wire  _GEN_2289 = branchEvalIn_fired ? _GEN_1642 : reservedFreeList3_49; // @[decode.scala 352:28 317:30]
  wire  _GEN_2290 = branchEvalIn_fired ? _GEN_1643 : reservedFreeList3_50; // @[decode.scala 352:28 317:30]
  wire  _GEN_2291 = branchEvalIn_fired ? _GEN_1644 : reservedFreeList3_51; // @[decode.scala 352:28 317:30]
  wire  _GEN_2292 = branchEvalIn_fired ? _GEN_1645 : reservedFreeList3_52; // @[decode.scala 352:28 317:30]
  wire  _GEN_2293 = branchEvalIn_fired ? _GEN_1646 : reservedFreeList3_53; // @[decode.scala 352:28 317:30]
  wire  _GEN_2294 = branchEvalIn_fired ? _GEN_1647 : reservedFreeList3_54; // @[decode.scala 352:28 317:30]
  wire  _GEN_2295 = branchEvalIn_fired ? _GEN_1648 : reservedFreeList3_55; // @[decode.scala 352:28 317:30]
  wire  _GEN_2296 = branchEvalIn_fired ? _GEN_1649 : reservedFreeList3_56; // @[decode.scala 352:28 317:30]
  wire  _GEN_2297 = branchEvalIn_fired ? _GEN_1650 : reservedFreeList3_57; // @[decode.scala 352:28 317:30]
  wire  _GEN_2298 = branchEvalIn_fired ? _GEN_1651 : reservedFreeList3_58; // @[decode.scala 352:28 317:30]
  wire  _GEN_2299 = branchEvalIn_fired ? _GEN_1652 : reservedFreeList3_59; // @[decode.scala 352:28 317:30]
  wire  _GEN_2300 = branchEvalIn_fired ? _GEN_1653 : reservedFreeList3_60; // @[decode.scala 352:28 317:30]
  wire  _GEN_2301 = branchEvalIn_fired ? _GEN_1654 : reservedFreeList3_61; // @[decode.scala 352:28 317:30]
  wire  _GEN_2302 = branchEvalIn_fired ? _GEN_1655 : reservedFreeList3_62; // @[decode.scala 352:28 317:30]
  wire  _GEN_2304 = branchEvalIn_fired ? _GEN_1657 : reservedValidList1_0; // @[decode.scala 352:28 320:31]
  wire  _GEN_2305 = branchEvalIn_fired ? _GEN_1658 : reservedValidList1_1; // @[decode.scala 352:28 320:31]
  wire  _GEN_2306 = branchEvalIn_fired ? _GEN_1659 : reservedValidList1_2; // @[decode.scala 352:28 320:31]
  wire  _GEN_2307 = branchEvalIn_fired ? _GEN_1660 : reservedValidList1_3; // @[decode.scala 352:28 320:31]
  wire  _GEN_2308 = branchEvalIn_fired ? _GEN_1661 : reservedValidList1_4; // @[decode.scala 352:28 320:31]
  wire  _GEN_2309 = branchEvalIn_fired ? _GEN_1662 : reservedValidList1_5; // @[decode.scala 352:28 320:31]
  wire  _GEN_2310 = branchEvalIn_fired ? _GEN_1663 : reservedValidList1_6; // @[decode.scala 352:28 320:31]
  wire  _GEN_2311 = branchEvalIn_fired ? _GEN_1664 : reservedValidList1_7; // @[decode.scala 352:28 320:31]
  wire  _GEN_2312 = branchEvalIn_fired ? _GEN_1665 : reservedValidList1_8; // @[decode.scala 352:28 320:31]
  wire  _GEN_2313 = branchEvalIn_fired ? _GEN_1666 : reservedValidList1_9; // @[decode.scala 352:28 320:31]
  wire  _GEN_2314 = branchEvalIn_fired ? _GEN_1667 : reservedValidList1_10; // @[decode.scala 352:28 320:31]
  wire  _GEN_2315 = branchEvalIn_fired ? _GEN_1668 : reservedValidList1_11; // @[decode.scala 352:28 320:31]
  wire  _GEN_2316 = branchEvalIn_fired ? _GEN_1669 : reservedValidList1_12; // @[decode.scala 352:28 320:31]
  wire  _GEN_2317 = branchEvalIn_fired ? _GEN_1670 : reservedValidList1_13; // @[decode.scala 352:28 320:31]
  wire  _GEN_2318 = branchEvalIn_fired ? _GEN_1671 : reservedValidList1_14; // @[decode.scala 352:28 320:31]
  wire  _GEN_2319 = branchEvalIn_fired ? _GEN_1672 : reservedValidList1_15; // @[decode.scala 352:28 320:31]
  wire  _GEN_2320 = branchEvalIn_fired ? _GEN_1673 : reservedValidList1_16; // @[decode.scala 352:28 320:31]
  wire  _GEN_2321 = branchEvalIn_fired ? _GEN_1674 : reservedValidList1_17; // @[decode.scala 352:28 320:31]
  wire  _GEN_2322 = branchEvalIn_fired ? _GEN_1675 : reservedValidList1_18; // @[decode.scala 352:28 320:31]
  wire  _GEN_2323 = branchEvalIn_fired ? _GEN_1676 : reservedValidList1_19; // @[decode.scala 352:28 320:31]
  wire  _GEN_2324 = branchEvalIn_fired ? _GEN_1677 : reservedValidList1_20; // @[decode.scala 352:28 320:31]
  wire  _GEN_2325 = branchEvalIn_fired ? _GEN_1678 : reservedValidList1_21; // @[decode.scala 352:28 320:31]
  wire  _GEN_2326 = branchEvalIn_fired ? _GEN_1679 : reservedValidList1_22; // @[decode.scala 352:28 320:31]
  wire  _GEN_2327 = branchEvalIn_fired ? _GEN_1680 : reservedValidList1_23; // @[decode.scala 352:28 320:31]
  wire  _GEN_2328 = branchEvalIn_fired ? _GEN_1681 : reservedValidList1_24; // @[decode.scala 352:28 320:31]
  wire  _GEN_2329 = branchEvalIn_fired ? _GEN_1682 : reservedValidList1_25; // @[decode.scala 352:28 320:31]
  wire  _GEN_2330 = branchEvalIn_fired ? _GEN_1683 : reservedValidList1_26; // @[decode.scala 352:28 320:31]
  wire  _GEN_2331 = branchEvalIn_fired ? _GEN_1684 : reservedValidList1_27; // @[decode.scala 352:28 320:31]
  wire  _GEN_2332 = branchEvalIn_fired ? _GEN_1685 : reservedValidList1_28; // @[decode.scala 352:28 320:31]
  wire  _GEN_2333 = branchEvalIn_fired ? _GEN_1686 : reservedValidList1_29; // @[decode.scala 352:28 320:31]
  wire  _GEN_2334 = branchEvalIn_fired ? _GEN_1687 : reservedValidList1_30; // @[decode.scala 352:28 320:31]
  wire  _GEN_2335 = branchEvalIn_fired ? _GEN_1688 : reservedValidList1_31; // @[decode.scala 352:28 320:31]
  wire  _GEN_2336 = branchEvalIn_fired ? _GEN_1689 : reservedValidList1_32; // @[decode.scala 352:28 320:31]
  wire  _GEN_2337 = branchEvalIn_fired ? _GEN_1690 : reservedValidList1_33; // @[decode.scala 352:28 320:31]
  wire  _GEN_2338 = branchEvalIn_fired ? _GEN_1691 : reservedValidList1_34; // @[decode.scala 352:28 320:31]
  wire  _GEN_2339 = branchEvalIn_fired ? _GEN_1692 : reservedValidList1_35; // @[decode.scala 352:28 320:31]
  wire  _GEN_2340 = branchEvalIn_fired ? _GEN_1693 : reservedValidList1_36; // @[decode.scala 352:28 320:31]
  wire  _GEN_2341 = branchEvalIn_fired ? _GEN_1694 : reservedValidList1_37; // @[decode.scala 352:28 320:31]
  wire  _GEN_2342 = branchEvalIn_fired ? _GEN_1695 : reservedValidList1_38; // @[decode.scala 352:28 320:31]
  wire  _GEN_2343 = branchEvalIn_fired ? _GEN_1696 : reservedValidList1_39; // @[decode.scala 352:28 320:31]
  wire  _GEN_2344 = branchEvalIn_fired ? _GEN_1697 : reservedValidList1_40; // @[decode.scala 352:28 320:31]
  wire  _GEN_2345 = branchEvalIn_fired ? _GEN_1698 : reservedValidList1_41; // @[decode.scala 352:28 320:31]
  wire  _GEN_2346 = branchEvalIn_fired ? _GEN_1699 : reservedValidList1_42; // @[decode.scala 352:28 320:31]
  wire  _GEN_2347 = branchEvalIn_fired ? _GEN_1700 : reservedValidList1_43; // @[decode.scala 352:28 320:31]
  wire  _GEN_2348 = branchEvalIn_fired ? _GEN_1701 : reservedValidList1_44; // @[decode.scala 352:28 320:31]
  wire  _GEN_2349 = branchEvalIn_fired ? _GEN_1702 : reservedValidList1_45; // @[decode.scala 352:28 320:31]
  wire  _GEN_2350 = branchEvalIn_fired ? _GEN_1703 : reservedValidList1_46; // @[decode.scala 352:28 320:31]
  wire  _GEN_2351 = branchEvalIn_fired ? _GEN_1704 : reservedValidList1_47; // @[decode.scala 352:28 320:31]
  wire  _GEN_2352 = branchEvalIn_fired ? _GEN_1705 : reservedValidList1_48; // @[decode.scala 352:28 320:31]
  wire  _GEN_2353 = branchEvalIn_fired ? _GEN_1706 : reservedValidList1_49; // @[decode.scala 352:28 320:31]
  wire  _GEN_2354 = branchEvalIn_fired ? _GEN_1707 : reservedValidList1_50; // @[decode.scala 352:28 320:31]
  wire  _GEN_2355 = branchEvalIn_fired ? _GEN_1708 : reservedValidList1_51; // @[decode.scala 352:28 320:31]
  wire  _GEN_2356 = branchEvalIn_fired ? _GEN_1709 : reservedValidList1_52; // @[decode.scala 352:28 320:31]
  wire  _GEN_2357 = branchEvalIn_fired ? _GEN_1710 : reservedValidList1_53; // @[decode.scala 352:28 320:31]
  wire  _GEN_2358 = branchEvalIn_fired ? _GEN_1711 : reservedValidList1_54; // @[decode.scala 352:28 320:31]
  wire  _GEN_2359 = branchEvalIn_fired ? _GEN_1712 : reservedValidList1_55; // @[decode.scala 352:28 320:31]
  wire  _GEN_2360 = branchEvalIn_fired ? _GEN_1713 : reservedValidList1_56; // @[decode.scala 352:28 320:31]
  wire  _GEN_2361 = branchEvalIn_fired ? _GEN_1714 : reservedValidList1_57; // @[decode.scala 352:28 320:31]
  wire  _GEN_2362 = branchEvalIn_fired ? _GEN_1715 : reservedValidList1_58; // @[decode.scala 352:28 320:31]
  wire  _GEN_2363 = branchEvalIn_fired ? _GEN_1716 : reservedValidList1_59; // @[decode.scala 352:28 320:31]
  wire  _GEN_2364 = branchEvalIn_fired ? _GEN_1717 : reservedValidList1_60; // @[decode.scala 352:28 320:31]
  wire  _GEN_2365 = branchEvalIn_fired ? _GEN_1718 : reservedValidList1_61; // @[decode.scala 352:28 320:31]
  wire  _GEN_2366 = branchEvalIn_fired ? _GEN_1719 : reservedValidList1_62; // @[decode.scala 352:28 320:31]
  wire  _GEN_2367 = branchEvalIn_fired ? _GEN_1720 : reservedValidList1_63; // @[decode.scala 352:28 320:31]
  wire  _GEN_2368 = branchEvalIn_fired ? _GEN_1721 : reservedValidList2_0; // @[decode.scala 352:28 321:31]
  wire  _GEN_2369 = branchEvalIn_fired ? _GEN_1722 : reservedValidList2_1; // @[decode.scala 352:28 321:31]
  wire  _GEN_2370 = branchEvalIn_fired ? _GEN_1723 : reservedValidList2_2; // @[decode.scala 352:28 321:31]
  wire  _GEN_2371 = branchEvalIn_fired ? _GEN_1724 : reservedValidList2_3; // @[decode.scala 352:28 321:31]
  wire  _GEN_2372 = branchEvalIn_fired ? _GEN_1725 : reservedValidList2_4; // @[decode.scala 352:28 321:31]
  wire  _GEN_2373 = branchEvalIn_fired ? _GEN_1726 : reservedValidList2_5; // @[decode.scala 352:28 321:31]
  wire  _GEN_2374 = branchEvalIn_fired ? _GEN_1727 : reservedValidList2_6; // @[decode.scala 352:28 321:31]
  wire  _GEN_2375 = branchEvalIn_fired ? _GEN_1728 : reservedValidList2_7; // @[decode.scala 352:28 321:31]
  wire  _GEN_2376 = branchEvalIn_fired ? _GEN_1729 : reservedValidList2_8; // @[decode.scala 352:28 321:31]
  wire  _GEN_2377 = branchEvalIn_fired ? _GEN_1730 : reservedValidList2_9; // @[decode.scala 352:28 321:31]
  wire  _GEN_2378 = branchEvalIn_fired ? _GEN_1731 : reservedValidList2_10; // @[decode.scala 352:28 321:31]
  wire  _GEN_2379 = branchEvalIn_fired ? _GEN_1732 : reservedValidList2_11; // @[decode.scala 352:28 321:31]
  wire  _GEN_2380 = branchEvalIn_fired ? _GEN_1733 : reservedValidList2_12; // @[decode.scala 352:28 321:31]
  wire  _GEN_2381 = branchEvalIn_fired ? _GEN_1734 : reservedValidList2_13; // @[decode.scala 352:28 321:31]
  wire  _GEN_2382 = branchEvalIn_fired ? _GEN_1735 : reservedValidList2_14; // @[decode.scala 352:28 321:31]
  wire  _GEN_2383 = branchEvalIn_fired ? _GEN_1736 : reservedValidList2_15; // @[decode.scala 352:28 321:31]
  wire  _GEN_2384 = branchEvalIn_fired ? _GEN_1737 : reservedValidList2_16; // @[decode.scala 352:28 321:31]
  wire  _GEN_2385 = branchEvalIn_fired ? _GEN_1738 : reservedValidList2_17; // @[decode.scala 352:28 321:31]
  wire  _GEN_2386 = branchEvalIn_fired ? _GEN_1739 : reservedValidList2_18; // @[decode.scala 352:28 321:31]
  wire  _GEN_2387 = branchEvalIn_fired ? _GEN_1740 : reservedValidList2_19; // @[decode.scala 352:28 321:31]
  wire  _GEN_2388 = branchEvalIn_fired ? _GEN_1741 : reservedValidList2_20; // @[decode.scala 352:28 321:31]
  wire  _GEN_2389 = branchEvalIn_fired ? _GEN_1742 : reservedValidList2_21; // @[decode.scala 352:28 321:31]
  wire  _GEN_2390 = branchEvalIn_fired ? _GEN_1743 : reservedValidList2_22; // @[decode.scala 352:28 321:31]
  wire  _GEN_2391 = branchEvalIn_fired ? _GEN_1744 : reservedValidList2_23; // @[decode.scala 352:28 321:31]
  wire  _GEN_2392 = branchEvalIn_fired ? _GEN_1745 : reservedValidList2_24; // @[decode.scala 352:28 321:31]
  wire  _GEN_2393 = branchEvalIn_fired ? _GEN_1746 : reservedValidList2_25; // @[decode.scala 352:28 321:31]
  wire  _GEN_2394 = branchEvalIn_fired ? _GEN_1747 : reservedValidList2_26; // @[decode.scala 352:28 321:31]
  wire  _GEN_2395 = branchEvalIn_fired ? _GEN_1748 : reservedValidList2_27; // @[decode.scala 352:28 321:31]
  wire  _GEN_2396 = branchEvalIn_fired ? _GEN_1749 : reservedValidList2_28; // @[decode.scala 352:28 321:31]
  wire  _GEN_2397 = branchEvalIn_fired ? _GEN_1750 : reservedValidList2_29; // @[decode.scala 352:28 321:31]
  wire  _GEN_2398 = branchEvalIn_fired ? _GEN_1751 : reservedValidList2_30; // @[decode.scala 352:28 321:31]
  wire  _GEN_2399 = branchEvalIn_fired ? _GEN_1752 : reservedValidList2_31; // @[decode.scala 352:28 321:31]
  wire  _GEN_2400 = branchEvalIn_fired ? _GEN_1753 : reservedValidList2_32; // @[decode.scala 352:28 321:31]
  wire  _GEN_2401 = branchEvalIn_fired ? _GEN_1754 : reservedValidList2_33; // @[decode.scala 352:28 321:31]
  wire  _GEN_2402 = branchEvalIn_fired ? _GEN_1755 : reservedValidList2_34; // @[decode.scala 352:28 321:31]
  wire  _GEN_2403 = branchEvalIn_fired ? _GEN_1756 : reservedValidList2_35; // @[decode.scala 352:28 321:31]
  wire  _GEN_2404 = branchEvalIn_fired ? _GEN_1757 : reservedValidList2_36; // @[decode.scala 352:28 321:31]
  wire  _GEN_2405 = branchEvalIn_fired ? _GEN_1758 : reservedValidList2_37; // @[decode.scala 352:28 321:31]
  wire  _GEN_2406 = branchEvalIn_fired ? _GEN_1759 : reservedValidList2_38; // @[decode.scala 352:28 321:31]
  wire  _GEN_2407 = branchEvalIn_fired ? _GEN_1760 : reservedValidList2_39; // @[decode.scala 352:28 321:31]
  wire  _GEN_2408 = branchEvalIn_fired ? _GEN_1761 : reservedValidList2_40; // @[decode.scala 352:28 321:31]
  wire  _GEN_2409 = branchEvalIn_fired ? _GEN_1762 : reservedValidList2_41; // @[decode.scala 352:28 321:31]
  wire  _GEN_2410 = branchEvalIn_fired ? _GEN_1763 : reservedValidList2_42; // @[decode.scala 352:28 321:31]
  wire  _GEN_2411 = branchEvalIn_fired ? _GEN_1764 : reservedValidList2_43; // @[decode.scala 352:28 321:31]
  wire  _GEN_2412 = branchEvalIn_fired ? _GEN_1765 : reservedValidList2_44; // @[decode.scala 352:28 321:31]
  wire  _GEN_2413 = branchEvalIn_fired ? _GEN_1766 : reservedValidList2_45; // @[decode.scala 352:28 321:31]
  wire  _GEN_2414 = branchEvalIn_fired ? _GEN_1767 : reservedValidList2_46; // @[decode.scala 352:28 321:31]
  wire  _GEN_2415 = branchEvalIn_fired ? _GEN_1768 : reservedValidList2_47; // @[decode.scala 352:28 321:31]
  wire  _GEN_2416 = branchEvalIn_fired ? _GEN_1769 : reservedValidList2_48; // @[decode.scala 352:28 321:31]
  wire  _GEN_2417 = branchEvalIn_fired ? _GEN_1770 : reservedValidList2_49; // @[decode.scala 352:28 321:31]
  wire  _GEN_2418 = branchEvalIn_fired ? _GEN_1771 : reservedValidList2_50; // @[decode.scala 352:28 321:31]
  wire  _GEN_2419 = branchEvalIn_fired ? _GEN_1772 : reservedValidList2_51; // @[decode.scala 352:28 321:31]
  wire  _GEN_2420 = branchEvalIn_fired ? _GEN_1773 : reservedValidList2_52; // @[decode.scala 352:28 321:31]
  wire  _GEN_2421 = branchEvalIn_fired ? _GEN_1774 : reservedValidList2_53; // @[decode.scala 352:28 321:31]
  wire  _GEN_2422 = branchEvalIn_fired ? _GEN_1775 : reservedValidList2_54; // @[decode.scala 352:28 321:31]
  wire  _GEN_2423 = branchEvalIn_fired ? _GEN_1776 : reservedValidList2_55; // @[decode.scala 352:28 321:31]
  wire  _GEN_2424 = branchEvalIn_fired ? _GEN_1777 : reservedValidList2_56; // @[decode.scala 352:28 321:31]
  wire  _GEN_2425 = branchEvalIn_fired ? _GEN_1778 : reservedValidList2_57; // @[decode.scala 352:28 321:31]
  wire  _GEN_2426 = branchEvalIn_fired ? _GEN_1779 : reservedValidList2_58; // @[decode.scala 352:28 321:31]
  wire  _GEN_2427 = branchEvalIn_fired ? _GEN_1780 : reservedValidList2_59; // @[decode.scala 352:28 321:31]
  wire  _GEN_2428 = branchEvalIn_fired ? _GEN_1781 : reservedValidList2_60; // @[decode.scala 352:28 321:31]
  wire  _GEN_2429 = branchEvalIn_fired ? _GEN_1782 : reservedValidList2_61; // @[decode.scala 352:28 321:31]
  wire  _GEN_2430 = branchEvalIn_fired ? _GEN_1783 : reservedValidList2_62; // @[decode.scala 352:28 321:31]
  wire  _GEN_2431 = branchEvalIn_fired ? _GEN_1784 : reservedValidList2_63; // @[decode.scala 352:28 321:31]
  wire  _GEN_2432 = branchEvalIn_fired ? _GEN_1785 : reservedValidList3_0; // @[decode.scala 352:28 322:31]
  wire  _GEN_2433 = branchEvalIn_fired ? _GEN_1786 : reservedValidList3_1; // @[decode.scala 352:28 322:31]
  wire  _GEN_2434 = branchEvalIn_fired ? _GEN_1787 : reservedValidList3_2; // @[decode.scala 352:28 322:31]
  wire  _GEN_2435 = branchEvalIn_fired ? _GEN_1788 : reservedValidList3_3; // @[decode.scala 352:28 322:31]
  wire  _GEN_2436 = branchEvalIn_fired ? _GEN_1789 : reservedValidList3_4; // @[decode.scala 352:28 322:31]
  wire  _GEN_2437 = branchEvalIn_fired ? _GEN_1790 : reservedValidList3_5; // @[decode.scala 352:28 322:31]
  wire  _GEN_2438 = branchEvalIn_fired ? _GEN_1791 : reservedValidList3_6; // @[decode.scala 352:28 322:31]
  wire  _GEN_2439 = branchEvalIn_fired ? _GEN_1792 : reservedValidList3_7; // @[decode.scala 352:28 322:31]
  wire  _GEN_2440 = branchEvalIn_fired ? _GEN_1793 : reservedValidList3_8; // @[decode.scala 352:28 322:31]
  wire  _GEN_2441 = branchEvalIn_fired ? _GEN_1794 : reservedValidList3_9; // @[decode.scala 352:28 322:31]
  wire  _GEN_2442 = branchEvalIn_fired ? _GEN_1795 : reservedValidList3_10; // @[decode.scala 352:28 322:31]
  wire  _GEN_2443 = branchEvalIn_fired ? _GEN_1796 : reservedValidList3_11; // @[decode.scala 352:28 322:31]
  wire  _GEN_2444 = branchEvalIn_fired ? _GEN_1797 : reservedValidList3_12; // @[decode.scala 352:28 322:31]
  wire  _GEN_2445 = branchEvalIn_fired ? _GEN_1798 : reservedValidList3_13; // @[decode.scala 352:28 322:31]
  wire  _GEN_2446 = branchEvalIn_fired ? _GEN_1799 : reservedValidList3_14; // @[decode.scala 352:28 322:31]
  wire  _GEN_2447 = branchEvalIn_fired ? _GEN_1800 : reservedValidList3_15; // @[decode.scala 352:28 322:31]
  wire  _GEN_2448 = branchEvalIn_fired ? _GEN_1801 : reservedValidList3_16; // @[decode.scala 352:28 322:31]
  wire  _GEN_2449 = branchEvalIn_fired ? _GEN_1802 : reservedValidList3_17; // @[decode.scala 352:28 322:31]
  wire  _GEN_2450 = branchEvalIn_fired ? _GEN_1803 : reservedValidList3_18; // @[decode.scala 352:28 322:31]
  wire  _GEN_2451 = branchEvalIn_fired ? _GEN_1804 : reservedValidList3_19; // @[decode.scala 352:28 322:31]
  wire  _GEN_2452 = branchEvalIn_fired ? _GEN_1805 : reservedValidList3_20; // @[decode.scala 352:28 322:31]
  wire  _GEN_2453 = branchEvalIn_fired ? _GEN_1806 : reservedValidList3_21; // @[decode.scala 352:28 322:31]
  wire  _GEN_2454 = branchEvalIn_fired ? _GEN_1807 : reservedValidList3_22; // @[decode.scala 352:28 322:31]
  wire  _GEN_2455 = branchEvalIn_fired ? _GEN_1808 : reservedValidList3_23; // @[decode.scala 352:28 322:31]
  wire  _GEN_2456 = branchEvalIn_fired ? _GEN_1809 : reservedValidList3_24; // @[decode.scala 352:28 322:31]
  wire  _GEN_2457 = branchEvalIn_fired ? _GEN_1810 : reservedValidList3_25; // @[decode.scala 352:28 322:31]
  wire  _GEN_2458 = branchEvalIn_fired ? _GEN_1811 : reservedValidList3_26; // @[decode.scala 352:28 322:31]
  wire  _GEN_2459 = branchEvalIn_fired ? _GEN_1812 : reservedValidList3_27; // @[decode.scala 352:28 322:31]
  wire  _GEN_2460 = branchEvalIn_fired ? _GEN_1813 : reservedValidList3_28; // @[decode.scala 352:28 322:31]
  wire  _GEN_2461 = branchEvalIn_fired ? _GEN_1814 : reservedValidList3_29; // @[decode.scala 352:28 322:31]
  wire  _GEN_2462 = branchEvalIn_fired ? _GEN_1815 : reservedValidList3_30; // @[decode.scala 352:28 322:31]
  wire  _GEN_2463 = branchEvalIn_fired ? _GEN_1816 : reservedValidList3_31; // @[decode.scala 352:28 322:31]
  wire  _GEN_2464 = branchEvalIn_fired ? _GEN_1817 : reservedValidList3_32; // @[decode.scala 352:28 322:31]
  wire  _GEN_2465 = branchEvalIn_fired ? _GEN_1818 : reservedValidList3_33; // @[decode.scala 352:28 322:31]
  wire  _GEN_2466 = branchEvalIn_fired ? _GEN_1819 : reservedValidList3_34; // @[decode.scala 352:28 322:31]
  wire  _GEN_2467 = branchEvalIn_fired ? _GEN_1820 : reservedValidList3_35; // @[decode.scala 352:28 322:31]
  wire  _GEN_2468 = branchEvalIn_fired ? _GEN_1821 : reservedValidList3_36; // @[decode.scala 352:28 322:31]
  wire  _GEN_2469 = branchEvalIn_fired ? _GEN_1822 : reservedValidList3_37; // @[decode.scala 352:28 322:31]
  wire  _GEN_2470 = branchEvalIn_fired ? _GEN_1823 : reservedValidList3_38; // @[decode.scala 352:28 322:31]
  wire  _GEN_2471 = branchEvalIn_fired ? _GEN_1824 : reservedValidList3_39; // @[decode.scala 352:28 322:31]
  wire  _GEN_2472 = branchEvalIn_fired ? _GEN_1825 : reservedValidList3_40; // @[decode.scala 352:28 322:31]
  wire  _GEN_2473 = branchEvalIn_fired ? _GEN_1826 : reservedValidList3_41; // @[decode.scala 352:28 322:31]
  wire  _GEN_2474 = branchEvalIn_fired ? _GEN_1827 : reservedValidList3_42; // @[decode.scala 352:28 322:31]
  wire  _GEN_2475 = branchEvalIn_fired ? _GEN_1828 : reservedValidList3_43; // @[decode.scala 352:28 322:31]
  wire  _GEN_2476 = branchEvalIn_fired ? _GEN_1829 : reservedValidList3_44; // @[decode.scala 352:28 322:31]
  wire  _GEN_2477 = branchEvalIn_fired ? _GEN_1830 : reservedValidList3_45; // @[decode.scala 352:28 322:31]
  wire  _GEN_2478 = branchEvalIn_fired ? _GEN_1831 : reservedValidList3_46; // @[decode.scala 352:28 322:31]
  wire  _GEN_2479 = branchEvalIn_fired ? _GEN_1832 : reservedValidList3_47; // @[decode.scala 352:28 322:31]
  wire  _GEN_2480 = branchEvalIn_fired ? _GEN_1833 : reservedValidList3_48; // @[decode.scala 352:28 322:31]
  wire  _GEN_2481 = branchEvalIn_fired ? _GEN_1834 : reservedValidList3_49; // @[decode.scala 352:28 322:31]
  wire  _GEN_2482 = branchEvalIn_fired ? _GEN_1835 : reservedValidList3_50; // @[decode.scala 352:28 322:31]
  wire  _GEN_2483 = branchEvalIn_fired ? _GEN_1836 : reservedValidList3_51; // @[decode.scala 352:28 322:31]
  wire  _GEN_2484 = branchEvalIn_fired ? _GEN_1837 : reservedValidList3_52; // @[decode.scala 352:28 322:31]
  wire  _GEN_2485 = branchEvalIn_fired ? _GEN_1838 : reservedValidList3_53; // @[decode.scala 352:28 322:31]
  wire  _GEN_2486 = branchEvalIn_fired ? _GEN_1839 : reservedValidList3_54; // @[decode.scala 352:28 322:31]
  wire  _GEN_2487 = branchEvalIn_fired ? _GEN_1840 : reservedValidList3_55; // @[decode.scala 352:28 322:31]
  wire  _GEN_2488 = branchEvalIn_fired ? _GEN_1841 : reservedValidList3_56; // @[decode.scala 352:28 322:31]
  wire  _GEN_2489 = branchEvalIn_fired ? _GEN_1842 : reservedValidList3_57; // @[decode.scala 352:28 322:31]
  wire  _GEN_2490 = branchEvalIn_fired ? _GEN_1843 : reservedValidList3_58; // @[decode.scala 352:28 322:31]
  wire  _GEN_2491 = branchEvalIn_fired ? _GEN_1844 : reservedValidList3_59; // @[decode.scala 352:28 322:31]
  wire  _GEN_2492 = branchEvalIn_fired ? _GEN_1845 : reservedValidList3_60; // @[decode.scala 352:28 322:31]
  wire  _GEN_2493 = branchEvalIn_fired ? _GEN_1846 : reservedValidList3_61; // @[decode.scala 352:28 322:31]
  wire  _GEN_2494 = branchEvalIn_fired ? _GEN_1847 : reservedValidList3_62; // @[decode.scala 352:28 322:31]
  wire  _GEN_2495 = branchEvalIn_fired ? _GEN_1848 : reservedValidList3_63; // @[decode.scala 352:28 322:31]
  wire [3:0] _bitPosition_T_1 = ~_toExec_branchMask_T; // @[decode.scala 386:34]
  wire [1:0] _bitPosition_T_6 = _bitPosition_T_1[2] ? 2'h2 : 2'h3; // @[Mux.scala 47:70]
  wire [1:0] _bitPosition_T_7 = _bitPosition_T_1[1] ? 2'h1 : _bitPosition_T_6; // @[Mux.scala 47:70]
  wire [1:0] bitPosition = _bitPosition_T_1[0] ? 2'h0 : _bitPosition_T_7; // @[Mux.scala 47:70]
  wire  _T_181 = _T_432 | _T_434 | _T_431; // @[decode.scala 389:50]
  wire  _GEN_9879 = 2'h0 == bitPosition; // @[decode.scala 392:{44,44}]
  wire  _GEN_2496 = 2'h0 == bitPosition | _GEN_1850; // @[decode.scala 392:{44,44}]
  wire  _GEN_9880 = 2'h1 == bitPosition; // @[decode.scala 392:{44,44}]
  wire  _GEN_2497 = 2'h1 == bitPosition | _GEN_1851; // @[decode.scala 392:{44,44}]
  wire  _GEN_9881 = 2'h2 == bitPosition; // @[decode.scala 392:{44,44}]
  wire  _GEN_2498 = 2'h2 == bitPosition | _GEN_1852; // @[decode.scala 392:{44,44}]
  wire  _GEN_9882 = 2'h3 == bitPosition; // @[decode.scala 392:{44,44}]
  wire  _GEN_2499 = 2'h3 == bitPosition | _GEN_1853; // @[decode.scala 392:{44,44}]
  wire [3:0] _GEN_2500 = _GEN_9882 ? 4'h8 : branchPCMask; // @[decode.scala 393:27 219:29 397:32]
  wire [3:0] _GEN_2501 = _GEN_9881 ? 4'h4 : _GEN_2500; // @[decode.scala 393:27 396:32]
  wire [3:0] _GEN_2502 = _GEN_9880 ? 4'h2 : _GEN_2501; // @[decode.scala 393:27 395:32]
  wire  _GEN_2536 = 6'h0 == freeRegAddr ? 1'h0 : PRFFreeList_0; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2537 = 6'h1 == freeRegAddr ? 1'h0 : PRFFreeList_1; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2538 = 6'h2 == freeRegAddr ? 1'h0 : PRFFreeList_2; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2539 = 6'h3 == freeRegAddr ? 1'h0 : PRFFreeList_3; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2540 = 6'h4 == freeRegAddr ? 1'h0 : PRFFreeList_4; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2541 = 6'h5 == freeRegAddr ? 1'h0 : PRFFreeList_5; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2542 = 6'h6 == freeRegAddr ? 1'h0 : PRFFreeList_6; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2543 = 6'h7 == freeRegAddr ? 1'h0 : PRFFreeList_7; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2544 = 6'h8 == freeRegAddr ? 1'h0 : PRFFreeList_8; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2545 = 6'h9 == freeRegAddr ? 1'h0 : PRFFreeList_9; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2546 = 6'ha == freeRegAddr ? 1'h0 : PRFFreeList_10; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2547 = 6'hb == freeRegAddr ? 1'h0 : PRFFreeList_11; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2548 = 6'hc == freeRegAddr ? 1'h0 : PRFFreeList_12; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2549 = 6'hd == freeRegAddr ? 1'h0 : PRFFreeList_13; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2550 = 6'he == freeRegAddr ? 1'h0 : PRFFreeList_14; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2551 = 6'hf == freeRegAddr ? 1'h0 : PRFFreeList_15; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2552 = 6'h10 == freeRegAddr ? 1'h0 : PRFFreeList_16; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2553 = 6'h11 == freeRegAddr ? 1'h0 : PRFFreeList_17; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2554 = 6'h12 == freeRegAddr ? 1'h0 : PRFFreeList_18; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2555 = 6'h13 == freeRegAddr ? 1'h0 : PRFFreeList_19; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2556 = 6'h14 == freeRegAddr ? 1'h0 : PRFFreeList_20; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2557 = 6'h15 == freeRegAddr ? 1'h0 : PRFFreeList_21; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2558 = 6'h16 == freeRegAddr ? 1'h0 : PRFFreeList_22; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2559 = 6'h17 == freeRegAddr ? 1'h0 : PRFFreeList_23; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2560 = 6'h18 == freeRegAddr ? 1'h0 : PRFFreeList_24; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2561 = 6'h19 == freeRegAddr ? 1'h0 : PRFFreeList_25; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2562 = 6'h1a == freeRegAddr ? 1'h0 : PRFFreeList_26; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2563 = 6'h1b == freeRegAddr ? 1'h0 : PRFFreeList_27; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2564 = 6'h1c == freeRegAddr ? 1'h0 : PRFFreeList_28; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2565 = 6'h1d == freeRegAddr ? 1'h0 : PRFFreeList_29; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2566 = 6'h1e == freeRegAddr ? 1'h0 : PRFFreeList_30; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2567 = 6'h1f == freeRegAddr ? 1'h0 : PRFFreeList_31; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2568 = 6'h20 == freeRegAddr ? 1'h0 : PRFFreeList_32; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2569 = 6'h21 == freeRegAddr ? 1'h0 : PRFFreeList_33; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2570 = 6'h22 == freeRegAddr ? 1'h0 : PRFFreeList_34; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2571 = 6'h23 == freeRegAddr ? 1'h0 : PRFFreeList_35; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2572 = 6'h24 == freeRegAddr ? 1'h0 : PRFFreeList_36; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2573 = 6'h25 == freeRegAddr ? 1'h0 : PRFFreeList_37; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2574 = 6'h26 == freeRegAddr ? 1'h0 : PRFFreeList_38; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2575 = 6'h27 == freeRegAddr ? 1'h0 : PRFFreeList_39; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2576 = 6'h28 == freeRegAddr ? 1'h0 : PRFFreeList_40; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2577 = 6'h29 == freeRegAddr ? 1'h0 : PRFFreeList_41; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2578 = 6'h2a == freeRegAddr ? 1'h0 : PRFFreeList_42; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2579 = 6'h2b == freeRegAddr ? 1'h0 : PRFFreeList_43; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2580 = 6'h2c == freeRegAddr ? 1'h0 : PRFFreeList_44; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2581 = 6'h2d == freeRegAddr ? 1'h0 : PRFFreeList_45; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2582 = 6'h2e == freeRegAddr ? 1'h0 : PRFFreeList_46; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2583 = 6'h2f == freeRegAddr ? 1'h0 : PRFFreeList_47; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2584 = 6'h30 == freeRegAddr ? 1'h0 : PRFFreeList_48; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2585 = 6'h31 == freeRegAddr ? 1'h0 : PRFFreeList_49; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2586 = 6'h32 == freeRegAddr ? 1'h0 : PRFFreeList_50; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2587 = 6'h33 == freeRegAddr ? 1'h0 : PRFFreeList_51; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2588 = 6'h34 == freeRegAddr ? 1'h0 : PRFFreeList_52; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2589 = 6'h35 == freeRegAddr ? 1'h0 : PRFFreeList_53; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2590 = 6'h36 == freeRegAddr ? 1'h0 : PRFFreeList_54; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2591 = 6'h37 == freeRegAddr ? 1'h0 : PRFFreeList_55; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2592 = 6'h38 == freeRegAddr ? 1'h0 : PRFFreeList_56; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2593 = 6'h39 == freeRegAddr ? 1'h0 : PRFFreeList_57; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2594 = 6'h3a == freeRegAddr ? 1'h0 : PRFFreeList_58; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2595 = 6'h3b == freeRegAddr ? 1'h0 : PRFFreeList_59; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2596 = 6'h3c == freeRegAddr ? 1'h0 : PRFFreeList_60; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2597 = 6'h3d == freeRegAddr ? 1'h0 : PRFFreeList_61; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2598 = 6'h3e == freeRegAddr ? 1'h0 : PRFFreeList_62; // @[decode.scala 403:30 407:{45,45}]
  wire  _GEN_2600 = 6'h0 == freeRegAddr ? 1'h0 : PRFValidList_0; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2601 = 6'h1 == freeRegAddr ? 1'h0 : PRFValidList_1; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2602 = 6'h2 == freeRegAddr ? 1'h0 : PRFValidList_2; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2603 = 6'h3 == freeRegAddr ? 1'h0 : PRFValidList_3; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2604 = 6'h4 == freeRegAddr ? 1'h0 : PRFValidList_4; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2605 = 6'h5 == freeRegAddr ? 1'h0 : PRFValidList_5; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2606 = 6'h6 == freeRegAddr ? 1'h0 : PRFValidList_6; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2607 = 6'h7 == freeRegAddr ? 1'h0 : PRFValidList_7; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2608 = 6'h8 == freeRegAddr ? 1'h0 : PRFValidList_8; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2609 = 6'h9 == freeRegAddr ? 1'h0 : PRFValidList_9; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2610 = 6'ha == freeRegAddr ? 1'h0 : PRFValidList_10; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2611 = 6'hb == freeRegAddr ? 1'h0 : PRFValidList_11; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2612 = 6'hc == freeRegAddr ? 1'h0 : PRFValidList_12; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2613 = 6'hd == freeRegAddr ? 1'h0 : PRFValidList_13; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2614 = 6'he == freeRegAddr ? 1'h0 : PRFValidList_14; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2615 = 6'hf == freeRegAddr ? 1'h0 : PRFValidList_15; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2616 = 6'h10 == freeRegAddr ? 1'h0 : PRFValidList_16; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2617 = 6'h11 == freeRegAddr ? 1'h0 : PRFValidList_17; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2618 = 6'h12 == freeRegAddr ? 1'h0 : PRFValidList_18; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2619 = 6'h13 == freeRegAddr ? 1'h0 : PRFValidList_19; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2620 = 6'h14 == freeRegAddr ? 1'h0 : PRFValidList_20; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2621 = 6'h15 == freeRegAddr ? 1'h0 : PRFValidList_21; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2622 = 6'h16 == freeRegAddr ? 1'h0 : PRFValidList_22; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2623 = 6'h17 == freeRegAddr ? 1'h0 : PRFValidList_23; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2624 = 6'h18 == freeRegAddr ? 1'h0 : PRFValidList_24; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2625 = 6'h19 == freeRegAddr ? 1'h0 : PRFValidList_25; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2626 = 6'h1a == freeRegAddr ? 1'h0 : PRFValidList_26; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2627 = 6'h1b == freeRegAddr ? 1'h0 : PRFValidList_27; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2628 = 6'h1c == freeRegAddr ? 1'h0 : PRFValidList_28; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2629 = 6'h1d == freeRegAddr ? 1'h0 : PRFValidList_29; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2630 = 6'h1e == freeRegAddr ? 1'h0 : PRFValidList_30; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2631 = 6'h1f == freeRegAddr ? 1'h0 : PRFValidList_31; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2632 = 6'h20 == freeRegAddr ? 1'h0 : PRFValidList_32; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2633 = 6'h21 == freeRegAddr ? 1'h0 : PRFValidList_33; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2634 = 6'h22 == freeRegAddr ? 1'h0 : PRFValidList_34; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2635 = 6'h23 == freeRegAddr ? 1'h0 : PRFValidList_35; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2636 = 6'h24 == freeRegAddr ? 1'h0 : PRFValidList_36; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2637 = 6'h25 == freeRegAddr ? 1'h0 : PRFValidList_37; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2638 = 6'h26 == freeRegAddr ? 1'h0 : PRFValidList_38; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2639 = 6'h27 == freeRegAddr ? 1'h0 : PRFValidList_39; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2640 = 6'h28 == freeRegAddr ? 1'h0 : PRFValidList_40; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2641 = 6'h29 == freeRegAddr ? 1'h0 : PRFValidList_41; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2642 = 6'h2a == freeRegAddr ? 1'h0 : PRFValidList_42; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2643 = 6'h2b == freeRegAddr ? 1'h0 : PRFValidList_43; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2644 = 6'h2c == freeRegAddr ? 1'h0 : PRFValidList_44; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2645 = 6'h2d == freeRegAddr ? 1'h0 : PRFValidList_45; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2646 = 6'h2e == freeRegAddr ? 1'h0 : PRFValidList_46; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2647 = 6'h2f == freeRegAddr ? 1'h0 : PRFValidList_47; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2648 = 6'h30 == freeRegAddr ? 1'h0 : PRFValidList_48; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2649 = 6'h31 == freeRegAddr ? 1'h0 : PRFValidList_49; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2650 = 6'h32 == freeRegAddr ? 1'h0 : PRFValidList_50; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2651 = 6'h33 == freeRegAddr ? 1'h0 : PRFValidList_51; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2652 = 6'h34 == freeRegAddr ? 1'h0 : PRFValidList_52; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2653 = 6'h35 == freeRegAddr ? 1'h0 : PRFValidList_53; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2654 = 6'h36 == freeRegAddr ? 1'h0 : PRFValidList_54; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2655 = 6'h37 == freeRegAddr ? 1'h0 : PRFValidList_55; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2656 = 6'h38 == freeRegAddr ? 1'h0 : PRFValidList_56; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2657 = 6'h39 == freeRegAddr ? 1'h0 : PRFValidList_57; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2658 = 6'h3a == freeRegAddr ? 1'h0 : PRFValidList_58; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2659 = 6'h3b == freeRegAddr ? 1'h0 : PRFValidList_59; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2660 = 6'h3c == freeRegAddr ? 1'h0 : PRFValidList_60; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2661 = 6'h3d == freeRegAddr ? 1'h0 : PRFValidList_61; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2662 = 6'h3e == freeRegAddr ? 1'h0 : PRFValidList_62; // @[decode.scala 404:30 408:{45,45}]
  wire  _GEN_2663 = 6'h3f == freeRegAddr ? 1'h0 : PRFValidList_63; // @[decode.scala 404:30 408:{45,45}]
  wire [5:0] _GEN_2664 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_850 : frontEndRegMap_0; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2665 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_851 : frontEndRegMap_1; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2666 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_852 : frontEndRegMap_2; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2667 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_853 : frontEndRegMap_3; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2668 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_854 : frontEndRegMap_4; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2669 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_855 : frontEndRegMap_5; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2670 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_856 : frontEndRegMap_6; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2671 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_857 : frontEndRegMap_7; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2672 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_858 : frontEndRegMap_8; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2673 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_859 : frontEndRegMap_9; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2674 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_860 : frontEndRegMap_10; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2675 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_861 : frontEndRegMap_11; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2676 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_862 : frontEndRegMap_12; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2677 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_863 : frontEndRegMap_13; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2678 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_864 : frontEndRegMap_14; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2679 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_865 : frontEndRegMap_15; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2680 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_866 : frontEndRegMap_16; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2681 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_867 : frontEndRegMap_17; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2682 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_868 : frontEndRegMap_18; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2683 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_869 : frontEndRegMap_19; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2684 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_870 : frontEndRegMap_20; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2685 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_871 : frontEndRegMap_21; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2686 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_872 : frontEndRegMap_22; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2687 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_873 : frontEndRegMap_23; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2688 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_874 : frontEndRegMap_24; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2689 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_875 : frontEndRegMap_25; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2690 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_876 : frontEndRegMap_26; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2691 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_877 : frontEndRegMap_27; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2692 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_878 : frontEndRegMap_28; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2693 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_879 : frontEndRegMap_29; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2694 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_880 : frontEndRegMap_30; // @[decode.scala 402:30 405:44]
  wire [5:0] _GEN_2695 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_881 : frontEndRegMap_31; // @[decode.scala 402:30 405:44]
  wire  _GEN_2696 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2536 : PRFFreeList_0; // @[decode.scala 403:30 405:44]
  wire  _GEN_2697 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2537 : PRFFreeList_1; // @[decode.scala 403:30 405:44]
  wire  _GEN_2698 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2538 : PRFFreeList_2; // @[decode.scala 403:30 405:44]
  wire  _GEN_2699 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2539 : PRFFreeList_3; // @[decode.scala 403:30 405:44]
  wire  _GEN_2700 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2540 : PRFFreeList_4; // @[decode.scala 403:30 405:44]
  wire  _GEN_2701 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2541 : PRFFreeList_5; // @[decode.scala 403:30 405:44]
  wire  _GEN_2702 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2542 : PRFFreeList_6; // @[decode.scala 403:30 405:44]
  wire  _GEN_2703 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2543 : PRFFreeList_7; // @[decode.scala 403:30 405:44]
  wire  _GEN_2704 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2544 : PRFFreeList_8; // @[decode.scala 403:30 405:44]
  wire  _GEN_2705 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2545 : PRFFreeList_9; // @[decode.scala 403:30 405:44]
  wire  _GEN_2706 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2546 : PRFFreeList_10; // @[decode.scala 403:30 405:44]
  wire  _GEN_2707 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2547 : PRFFreeList_11; // @[decode.scala 403:30 405:44]
  wire  _GEN_2708 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2548 : PRFFreeList_12; // @[decode.scala 403:30 405:44]
  wire  _GEN_2709 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2549 : PRFFreeList_13; // @[decode.scala 403:30 405:44]
  wire  _GEN_2710 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2550 : PRFFreeList_14; // @[decode.scala 403:30 405:44]
  wire  _GEN_2711 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2551 : PRFFreeList_15; // @[decode.scala 403:30 405:44]
  wire  _GEN_2712 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2552 : PRFFreeList_16; // @[decode.scala 403:30 405:44]
  wire  _GEN_2713 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2553 : PRFFreeList_17; // @[decode.scala 403:30 405:44]
  wire  _GEN_2714 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2554 : PRFFreeList_18; // @[decode.scala 403:30 405:44]
  wire  _GEN_2715 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2555 : PRFFreeList_19; // @[decode.scala 403:30 405:44]
  wire  _GEN_2716 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2556 : PRFFreeList_20; // @[decode.scala 403:30 405:44]
  wire  _GEN_2717 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2557 : PRFFreeList_21; // @[decode.scala 403:30 405:44]
  wire  _GEN_2718 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2558 : PRFFreeList_22; // @[decode.scala 403:30 405:44]
  wire  _GEN_2719 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2559 : PRFFreeList_23; // @[decode.scala 403:30 405:44]
  wire  _GEN_2720 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2560 : PRFFreeList_24; // @[decode.scala 403:30 405:44]
  wire  _GEN_2721 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2561 : PRFFreeList_25; // @[decode.scala 403:30 405:44]
  wire  _GEN_2722 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2562 : PRFFreeList_26; // @[decode.scala 403:30 405:44]
  wire  _GEN_2723 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2563 : PRFFreeList_27; // @[decode.scala 403:30 405:44]
  wire  _GEN_2724 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2564 : PRFFreeList_28; // @[decode.scala 403:30 405:44]
  wire  _GEN_2725 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2565 : PRFFreeList_29; // @[decode.scala 403:30 405:44]
  wire  _GEN_2726 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2566 : PRFFreeList_30; // @[decode.scala 403:30 405:44]
  wire  _GEN_2727 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2567 : PRFFreeList_31; // @[decode.scala 403:30 405:44]
  wire  _GEN_2728 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2568 : PRFFreeList_32; // @[decode.scala 403:30 405:44]
  wire  _GEN_2729 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2569 : PRFFreeList_33; // @[decode.scala 403:30 405:44]
  wire  _GEN_2730 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2570 : PRFFreeList_34; // @[decode.scala 403:30 405:44]
  wire  _GEN_2731 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2571 : PRFFreeList_35; // @[decode.scala 403:30 405:44]
  wire  _GEN_2732 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2572 : PRFFreeList_36; // @[decode.scala 403:30 405:44]
  wire  _GEN_2733 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2573 : PRFFreeList_37; // @[decode.scala 403:30 405:44]
  wire  _GEN_2734 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2574 : PRFFreeList_38; // @[decode.scala 403:30 405:44]
  wire  _GEN_2735 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2575 : PRFFreeList_39; // @[decode.scala 403:30 405:44]
  wire  _GEN_2736 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2576 : PRFFreeList_40; // @[decode.scala 403:30 405:44]
  wire  _GEN_2737 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2577 : PRFFreeList_41; // @[decode.scala 403:30 405:44]
  wire  _GEN_2738 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2578 : PRFFreeList_42; // @[decode.scala 403:30 405:44]
  wire  _GEN_2739 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2579 : PRFFreeList_43; // @[decode.scala 403:30 405:44]
  wire  _GEN_2740 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2580 : PRFFreeList_44; // @[decode.scala 403:30 405:44]
  wire  _GEN_2741 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2581 : PRFFreeList_45; // @[decode.scala 403:30 405:44]
  wire  _GEN_2742 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2582 : PRFFreeList_46; // @[decode.scala 403:30 405:44]
  wire  _GEN_2743 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2583 : PRFFreeList_47; // @[decode.scala 403:30 405:44]
  wire  _GEN_2744 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2584 : PRFFreeList_48; // @[decode.scala 403:30 405:44]
  wire  _GEN_2745 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2585 : PRFFreeList_49; // @[decode.scala 403:30 405:44]
  wire  _GEN_2746 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2586 : PRFFreeList_50; // @[decode.scala 403:30 405:44]
  wire  _GEN_2747 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2587 : PRFFreeList_51; // @[decode.scala 403:30 405:44]
  wire  _GEN_2748 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2588 : PRFFreeList_52; // @[decode.scala 403:30 405:44]
  wire  _GEN_2749 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2589 : PRFFreeList_53; // @[decode.scala 403:30 405:44]
  wire  _GEN_2750 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2590 : PRFFreeList_54; // @[decode.scala 403:30 405:44]
  wire  _GEN_2751 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2591 : PRFFreeList_55; // @[decode.scala 403:30 405:44]
  wire  _GEN_2752 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2592 : PRFFreeList_56; // @[decode.scala 403:30 405:44]
  wire  _GEN_2753 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2593 : PRFFreeList_57; // @[decode.scala 403:30 405:44]
  wire  _GEN_2754 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2594 : PRFFreeList_58; // @[decode.scala 403:30 405:44]
  wire  _GEN_2755 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2595 : PRFFreeList_59; // @[decode.scala 403:30 405:44]
  wire  _GEN_2756 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2596 : PRFFreeList_60; // @[decode.scala 403:30 405:44]
  wire  _GEN_2757 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2597 : PRFFreeList_61; // @[decode.scala 403:30 405:44]
  wire  _GEN_2758 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2598 : PRFFreeList_62; // @[decode.scala 403:30 405:44]
  wire  _GEN_2760 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2600 : PRFValidList_0; // @[decode.scala 404:30 405:44]
  wire  _GEN_2761 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2601 : PRFValidList_1; // @[decode.scala 404:30 405:44]
  wire  _GEN_2762 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2602 : PRFValidList_2; // @[decode.scala 404:30 405:44]
  wire  _GEN_2763 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2603 : PRFValidList_3; // @[decode.scala 404:30 405:44]
  wire  _GEN_2764 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2604 : PRFValidList_4; // @[decode.scala 404:30 405:44]
  wire  _GEN_2765 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2605 : PRFValidList_5; // @[decode.scala 404:30 405:44]
  wire  _GEN_2766 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2606 : PRFValidList_6; // @[decode.scala 404:30 405:44]
  wire  _GEN_2767 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2607 : PRFValidList_7; // @[decode.scala 404:30 405:44]
  wire  _GEN_2768 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2608 : PRFValidList_8; // @[decode.scala 404:30 405:44]
  wire  _GEN_2769 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2609 : PRFValidList_9; // @[decode.scala 404:30 405:44]
  wire  _GEN_2770 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2610 : PRFValidList_10; // @[decode.scala 404:30 405:44]
  wire  _GEN_2771 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2611 : PRFValidList_11; // @[decode.scala 404:30 405:44]
  wire  _GEN_2772 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2612 : PRFValidList_12; // @[decode.scala 404:30 405:44]
  wire  _GEN_2773 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2613 : PRFValidList_13; // @[decode.scala 404:30 405:44]
  wire  _GEN_2774 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2614 : PRFValidList_14; // @[decode.scala 404:30 405:44]
  wire  _GEN_2775 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2615 : PRFValidList_15; // @[decode.scala 404:30 405:44]
  wire  _GEN_2776 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2616 : PRFValidList_16; // @[decode.scala 404:30 405:44]
  wire  _GEN_2777 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2617 : PRFValidList_17; // @[decode.scala 404:30 405:44]
  wire  _GEN_2778 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2618 : PRFValidList_18; // @[decode.scala 404:30 405:44]
  wire  _GEN_2779 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2619 : PRFValidList_19; // @[decode.scala 404:30 405:44]
  wire  _GEN_2780 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2620 : PRFValidList_20; // @[decode.scala 404:30 405:44]
  wire  _GEN_2781 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2621 : PRFValidList_21; // @[decode.scala 404:30 405:44]
  wire  _GEN_2782 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2622 : PRFValidList_22; // @[decode.scala 404:30 405:44]
  wire  _GEN_2783 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2623 : PRFValidList_23; // @[decode.scala 404:30 405:44]
  wire  _GEN_2784 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2624 : PRFValidList_24; // @[decode.scala 404:30 405:44]
  wire  _GEN_2785 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2625 : PRFValidList_25; // @[decode.scala 404:30 405:44]
  wire  _GEN_2786 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2626 : PRFValidList_26; // @[decode.scala 404:30 405:44]
  wire  _GEN_2787 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2627 : PRFValidList_27; // @[decode.scala 404:30 405:44]
  wire  _GEN_2788 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2628 : PRFValidList_28; // @[decode.scala 404:30 405:44]
  wire  _GEN_2789 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2629 : PRFValidList_29; // @[decode.scala 404:30 405:44]
  wire  _GEN_2790 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2630 : PRFValidList_30; // @[decode.scala 404:30 405:44]
  wire  _GEN_2791 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2631 : PRFValidList_31; // @[decode.scala 404:30 405:44]
  wire  _GEN_2792 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2632 : PRFValidList_32; // @[decode.scala 404:30 405:44]
  wire  _GEN_2793 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2633 : PRFValidList_33; // @[decode.scala 404:30 405:44]
  wire  _GEN_2794 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2634 : PRFValidList_34; // @[decode.scala 404:30 405:44]
  wire  _GEN_2795 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2635 : PRFValidList_35; // @[decode.scala 404:30 405:44]
  wire  _GEN_2796 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2636 : PRFValidList_36; // @[decode.scala 404:30 405:44]
  wire  _GEN_2797 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2637 : PRFValidList_37; // @[decode.scala 404:30 405:44]
  wire  _GEN_2798 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2638 : PRFValidList_38; // @[decode.scala 404:30 405:44]
  wire  _GEN_2799 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2639 : PRFValidList_39; // @[decode.scala 404:30 405:44]
  wire  _GEN_2800 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2640 : PRFValidList_40; // @[decode.scala 404:30 405:44]
  wire  _GEN_2801 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2641 : PRFValidList_41; // @[decode.scala 404:30 405:44]
  wire  _GEN_2802 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2642 : PRFValidList_42; // @[decode.scala 404:30 405:44]
  wire  _GEN_2803 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2643 : PRFValidList_43; // @[decode.scala 404:30 405:44]
  wire  _GEN_2804 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2644 : PRFValidList_44; // @[decode.scala 404:30 405:44]
  wire  _GEN_2805 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2645 : PRFValidList_45; // @[decode.scala 404:30 405:44]
  wire  _GEN_2806 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2646 : PRFValidList_46; // @[decode.scala 404:30 405:44]
  wire  _GEN_2807 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2647 : PRFValidList_47; // @[decode.scala 404:30 405:44]
  wire  _GEN_2808 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2648 : PRFValidList_48; // @[decode.scala 404:30 405:44]
  wire  _GEN_2809 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2649 : PRFValidList_49; // @[decode.scala 404:30 405:44]
  wire  _GEN_2810 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2650 : PRFValidList_50; // @[decode.scala 404:30 405:44]
  wire  _GEN_2811 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2651 : PRFValidList_51; // @[decode.scala 404:30 405:44]
  wire  _GEN_2812 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2652 : PRFValidList_52; // @[decode.scala 404:30 405:44]
  wire  _GEN_2813 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2653 : PRFValidList_53; // @[decode.scala 404:30 405:44]
  wire  _GEN_2814 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2654 : PRFValidList_54; // @[decode.scala 404:30 405:44]
  wire  _GEN_2815 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2655 : PRFValidList_55; // @[decode.scala 404:30 405:44]
  wire  _GEN_2816 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2656 : PRFValidList_56; // @[decode.scala 404:30 405:44]
  wire  _GEN_2817 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2657 : PRFValidList_57; // @[decode.scala 404:30 405:44]
  wire  _GEN_2818 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2658 : PRFValidList_58; // @[decode.scala 404:30 405:44]
  wire  _GEN_2819 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2659 : PRFValidList_59; // @[decode.scala 404:30 405:44]
  wire  _GEN_2820 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2660 : PRFValidList_60; // @[decode.scala 404:30 405:44]
  wire  _GEN_2821 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2661 : PRFValidList_61; // @[decode.scala 404:30 405:44]
  wire  _GEN_2822 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2662 : PRFValidList_62; // @[decode.scala 404:30 405:44]
  wire  _GEN_2823 = opcode[2] & |inputBuffer_instruction[11:7] ? _GEN_2663 : PRFValidList_63; // @[decode.scala 404:30 405:44]
  wire [5:0] _GEN_3784 = 3'h3 == branchTracker ? _GEN_2664 : reservedRegMap4_0; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3785 = 3'h3 == branchTracker ? _GEN_2665 : reservedRegMap4_1; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3786 = 3'h3 == branchTracker ? _GEN_2666 : reservedRegMap4_2; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3787 = 3'h3 == branchTracker ? _GEN_2667 : reservedRegMap4_3; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3788 = 3'h3 == branchTracker ? _GEN_2668 : reservedRegMap4_4; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3789 = 3'h3 == branchTracker ? _GEN_2669 : reservedRegMap4_5; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3790 = 3'h3 == branchTracker ? _GEN_2670 : reservedRegMap4_6; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3791 = 3'h3 == branchTracker ? _GEN_2671 : reservedRegMap4_7; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3792 = 3'h3 == branchTracker ? _GEN_2672 : reservedRegMap4_8; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3793 = 3'h3 == branchTracker ? _GEN_2673 : reservedRegMap4_9; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3794 = 3'h3 == branchTracker ? _GEN_2674 : reservedRegMap4_10; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3795 = 3'h3 == branchTracker ? _GEN_2675 : reservedRegMap4_11; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3796 = 3'h3 == branchTracker ? _GEN_2676 : reservedRegMap4_12; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3797 = 3'h3 == branchTracker ? _GEN_2677 : reservedRegMap4_13; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3798 = 3'h3 == branchTracker ? _GEN_2678 : reservedRegMap4_14; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3799 = 3'h3 == branchTracker ? _GEN_2679 : reservedRegMap4_15; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3800 = 3'h3 == branchTracker ? _GEN_2680 : reservedRegMap4_16; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3801 = 3'h3 == branchTracker ? _GEN_2681 : reservedRegMap4_17; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3802 = 3'h3 == branchTracker ? _GEN_2682 : reservedRegMap4_18; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3803 = 3'h3 == branchTracker ? _GEN_2683 : reservedRegMap4_19; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3804 = 3'h3 == branchTracker ? _GEN_2684 : reservedRegMap4_20; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3805 = 3'h3 == branchTracker ? _GEN_2685 : reservedRegMap4_21; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3806 = 3'h3 == branchTracker ? _GEN_2686 : reservedRegMap4_22; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3807 = 3'h3 == branchTracker ? _GEN_2687 : reservedRegMap4_23; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3808 = 3'h3 == branchTracker ? _GEN_2688 : reservedRegMap4_24; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3809 = 3'h3 == branchTracker ? _GEN_2689 : reservedRegMap4_25; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3810 = 3'h3 == branchTracker ? _GEN_2690 : reservedRegMap4_26; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3811 = 3'h3 == branchTracker ? _GEN_2691 : reservedRegMap4_27; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3812 = 3'h3 == branchTracker ? _GEN_2692 : reservedRegMap4_28; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3813 = 3'h3 == branchTracker ? _GEN_2693 : reservedRegMap4_29; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3814 = 3'h3 == branchTracker ? _GEN_2694 : reservedRegMap4_30; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_3815 = 3'h3 == branchTracker ? _GEN_2695 : reservedRegMap4_31; // @[decode.scala 313:28 400:29]
  wire  _GEN_3816 = 3'h3 == branchTracker ? _GEN_2696 : reservedFreeList4_0; // @[decode.scala 400:29 318:30]
  wire  _GEN_3817 = 3'h3 == branchTracker ? _GEN_2697 : reservedFreeList4_1; // @[decode.scala 400:29 318:30]
  wire  _GEN_3818 = 3'h3 == branchTracker ? _GEN_2698 : reservedFreeList4_2; // @[decode.scala 400:29 318:30]
  wire  _GEN_3819 = 3'h3 == branchTracker ? _GEN_2699 : reservedFreeList4_3; // @[decode.scala 400:29 318:30]
  wire  _GEN_3820 = 3'h3 == branchTracker ? _GEN_2700 : reservedFreeList4_4; // @[decode.scala 400:29 318:30]
  wire  _GEN_3821 = 3'h3 == branchTracker ? _GEN_2701 : reservedFreeList4_5; // @[decode.scala 400:29 318:30]
  wire  _GEN_3822 = 3'h3 == branchTracker ? _GEN_2702 : reservedFreeList4_6; // @[decode.scala 400:29 318:30]
  wire  _GEN_3823 = 3'h3 == branchTracker ? _GEN_2703 : reservedFreeList4_7; // @[decode.scala 400:29 318:30]
  wire  _GEN_3824 = 3'h3 == branchTracker ? _GEN_2704 : reservedFreeList4_8; // @[decode.scala 400:29 318:30]
  wire  _GEN_3825 = 3'h3 == branchTracker ? _GEN_2705 : reservedFreeList4_9; // @[decode.scala 400:29 318:30]
  wire  _GEN_3826 = 3'h3 == branchTracker ? _GEN_2706 : reservedFreeList4_10; // @[decode.scala 400:29 318:30]
  wire  _GEN_3827 = 3'h3 == branchTracker ? _GEN_2707 : reservedFreeList4_11; // @[decode.scala 400:29 318:30]
  wire  _GEN_3828 = 3'h3 == branchTracker ? _GEN_2708 : reservedFreeList4_12; // @[decode.scala 400:29 318:30]
  wire  _GEN_3829 = 3'h3 == branchTracker ? _GEN_2709 : reservedFreeList4_13; // @[decode.scala 400:29 318:30]
  wire  _GEN_3830 = 3'h3 == branchTracker ? _GEN_2710 : reservedFreeList4_14; // @[decode.scala 400:29 318:30]
  wire  _GEN_3831 = 3'h3 == branchTracker ? _GEN_2711 : reservedFreeList4_15; // @[decode.scala 400:29 318:30]
  wire  _GEN_3832 = 3'h3 == branchTracker ? _GEN_2712 : reservedFreeList4_16; // @[decode.scala 400:29 318:30]
  wire  _GEN_3833 = 3'h3 == branchTracker ? _GEN_2713 : reservedFreeList4_17; // @[decode.scala 400:29 318:30]
  wire  _GEN_3834 = 3'h3 == branchTracker ? _GEN_2714 : reservedFreeList4_18; // @[decode.scala 400:29 318:30]
  wire  _GEN_3835 = 3'h3 == branchTracker ? _GEN_2715 : reservedFreeList4_19; // @[decode.scala 400:29 318:30]
  wire  _GEN_3836 = 3'h3 == branchTracker ? _GEN_2716 : reservedFreeList4_20; // @[decode.scala 400:29 318:30]
  wire  _GEN_3837 = 3'h3 == branchTracker ? _GEN_2717 : reservedFreeList4_21; // @[decode.scala 400:29 318:30]
  wire  _GEN_3838 = 3'h3 == branchTracker ? _GEN_2718 : reservedFreeList4_22; // @[decode.scala 400:29 318:30]
  wire  _GEN_3839 = 3'h3 == branchTracker ? _GEN_2719 : reservedFreeList4_23; // @[decode.scala 400:29 318:30]
  wire  _GEN_3840 = 3'h3 == branchTracker ? _GEN_2720 : reservedFreeList4_24; // @[decode.scala 400:29 318:30]
  wire  _GEN_3841 = 3'h3 == branchTracker ? _GEN_2721 : reservedFreeList4_25; // @[decode.scala 400:29 318:30]
  wire  _GEN_3842 = 3'h3 == branchTracker ? _GEN_2722 : reservedFreeList4_26; // @[decode.scala 400:29 318:30]
  wire  _GEN_3843 = 3'h3 == branchTracker ? _GEN_2723 : reservedFreeList4_27; // @[decode.scala 400:29 318:30]
  wire  _GEN_3844 = 3'h3 == branchTracker ? _GEN_2724 : reservedFreeList4_28; // @[decode.scala 400:29 318:30]
  wire  _GEN_3845 = 3'h3 == branchTracker ? _GEN_2725 : reservedFreeList4_29; // @[decode.scala 400:29 318:30]
  wire  _GEN_3846 = 3'h3 == branchTracker ? _GEN_2726 : reservedFreeList4_30; // @[decode.scala 400:29 318:30]
  wire  _GEN_3847 = 3'h3 == branchTracker ? _GEN_2727 : reservedFreeList4_31; // @[decode.scala 400:29 318:30]
  wire  _GEN_3848 = 3'h3 == branchTracker ? _GEN_2728 : reservedFreeList4_32; // @[decode.scala 400:29 318:30]
  wire  _GEN_3849 = 3'h3 == branchTracker ? _GEN_2729 : reservedFreeList4_33; // @[decode.scala 400:29 318:30]
  wire  _GEN_3850 = 3'h3 == branchTracker ? _GEN_2730 : reservedFreeList4_34; // @[decode.scala 400:29 318:30]
  wire  _GEN_3851 = 3'h3 == branchTracker ? _GEN_2731 : reservedFreeList4_35; // @[decode.scala 400:29 318:30]
  wire  _GEN_3852 = 3'h3 == branchTracker ? _GEN_2732 : reservedFreeList4_36; // @[decode.scala 400:29 318:30]
  wire  _GEN_3853 = 3'h3 == branchTracker ? _GEN_2733 : reservedFreeList4_37; // @[decode.scala 400:29 318:30]
  wire  _GEN_3854 = 3'h3 == branchTracker ? _GEN_2734 : reservedFreeList4_38; // @[decode.scala 400:29 318:30]
  wire  _GEN_3855 = 3'h3 == branchTracker ? _GEN_2735 : reservedFreeList4_39; // @[decode.scala 400:29 318:30]
  wire  _GEN_3856 = 3'h3 == branchTracker ? _GEN_2736 : reservedFreeList4_40; // @[decode.scala 400:29 318:30]
  wire  _GEN_3857 = 3'h3 == branchTracker ? _GEN_2737 : reservedFreeList4_41; // @[decode.scala 400:29 318:30]
  wire  _GEN_3858 = 3'h3 == branchTracker ? _GEN_2738 : reservedFreeList4_42; // @[decode.scala 400:29 318:30]
  wire  _GEN_3859 = 3'h3 == branchTracker ? _GEN_2739 : reservedFreeList4_43; // @[decode.scala 400:29 318:30]
  wire  _GEN_3860 = 3'h3 == branchTracker ? _GEN_2740 : reservedFreeList4_44; // @[decode.scala 400:29 318:30]
  wire  _GEN_3861 = 3'h3 == branchTracker ? _GEN_2741 : reservedFreeList4_45; // @[decode.scala 400:29 318:30]
  wire  _GEN_3862 = 3'h3 == branchTracker ? _GEN_2742 : reservedFreeList4_46; // @[decode.scala 400:29 318:30]
  wire  _GEN_3863 = 3'h3 == branchTracker ? _GEN_2743 : reservedFreeList4_47; // @[decode.scala 400:29 318:30]
  wire  _GEN_3864 = 3'h3 == branchTracker ? _GEN_2744 : reservedFreeList4_48; // @[decode.scala 400:29 318:30]
  wire  _GEN_3865 = 3'h3 == branchTracker ? _GEN_2745 : reservedFreeList4_49; // @[decode.scala 400:29 318:30]
  wire  _GEN_3866 = 3'h3 == branchTracker ? _GEN_2746 : reservedFreeList4_50; // @[decode.scala 400:29 318:30]
  wire  _GEN_3867 = 3'h3 == branchTracker ? _GEN_2747 : reservedFreeList4_51; // @[decode.scala 400:29 318:30]
  wire  _GEN_3868 = 3'h3 == branchTracker ? _GEN_2748 : reservedFreeList4_52; // @[decode.scala 400:29 318:30]
  wire  _GEN_3869 = 3'h3 == branchTracker ? _GEN_2749 : reservedFreeList4_53; // @[decode.scala 400:29 318:30]
  wire  _GEN_3870 = 3'h3 == branchTracker ? _GEN_2750 : reservedFreeList4_54; // @[decode.scala 400:29 318:30]
  wire  _GEN_3871 = 3'h3 == branchTracker ? _GEN_2751 : reservedFreeList4_55; // @[decode.scala 400:29 318:30]
  wire  _GEN_3872 = 3'h3 == branchTracker ? _GEN_2752 : reservedFreeList4_56; // @[decode.scala 400:29 318:30]
  wire  _GEN_3873 = 3'h3 == branchTracker ? _GEN_2753 : reservedFreeList4_57; // @[decode.scala 400:29 318:30]
  wire  _GEN_3874 = 3'h3 == branchTracker ? _GEN_2754 : reservedFreeList4_58; // @[decode.scala 400:29 318:30]
  wire  _GEN_3875 = 3'h3 == branchTracker ? _GEN_2755 : reservedFreeList4_59; // @[decode.scala 400:29 318:30]
  wire  _GEN_3876 = 3'h3 == branchTracker ? _GEN_2756 : reservedFreeList4_60; // @[decode.scala 400:29 318:30]
  wire  _GEN_3877 = 3'h3 == branchTracker ? _GEN_2757 : reservedFreeList4_61; // @[decode.scala 400:29 318:30]
  wire  _GEN_3878 = 3'h3 == branchTracker ? _GEN_2758 : reservedFreeList4_62; // @[decode.scala 400:29 318:30]
  wire  _GEN_3880 = 3'h3 == branchTracker ? _GEN_2760 : reservedValidList4_0; // @[decode.scala 400:29 323:31]
  wire  _GEN_3881 = 3'h3 == branchTracker ? _GEN_2761 : reservedValidList4_1; // @[decode.scala 400:29 323:31]
  wire  _GEN_3882 = 3'h3 == branchTracker ? _GEN_2762 : reservedValidList4_2; // @[decode.scala 400:29 323:31]
  wire  _GEN_3883 = 3'h3 == branchTracker ? _GEN_2763 : reservedValidList4_3; // @[decode.scala 400:29 323:31]
  wire  _GEN_3884 = 3'h3 == branchTracker ? _GEN_2764 : reservedValidList4_4; // @[decode.scala 400:29 323:31]
  wire  _GEN_3885 = 3'h3 == branchTracker ? _GEN_2765 : reservedValidList4_5; // @[decode.scala 400:29 323:31]
  wire  _GEN_3886 = 3'h3 == branchTracker ? _GEN_2766 : reservedValidList4_6; // @[decode.scala 400:29 323:31]
  wire  _GEN_3887 = 3'h3 == branchTracker ? _GEN_2767 : reservedValidList4_7; // @[decode.scala 400:29 323:31]
  wire  _GEN_3888 = 3'h3 == branchTracker ? _GEN_2768 : reservedValidList4_8; // @[decode.scala 400:29 323:31]
  wire  _GEN_3889 = 3'h3 == branchTracker ? _GEN_2769 : reservedValidList4_9; // @[decode.scala 400:29 323:31]
  wire  _GEN_3890 = 3'h3 == branchTracker ? _GEN_2770 : reservedValidList4_10; // @[decode.scala 400:29 323:31]
  wire  _GEN_3891 = 3'h3 == branchTracker ? _GEN_2771 : reservedValidList4_11; // @[decode.scala 400:29 323:31]
  wire  _GEN_3892 = 3'h3 == branchTracker ? _GEN_2772 : reservedValidList4_12; // @[decode.scala 400:29 323:31]
  wire  _GEN_3893 = 3'h3 == branchTracker ? _GEN_2773 : reservedValidList4_13; // @[decode.scala 400:29 323:31]
  wire  _GEN_3894 = 3'h3 == branchTracker ? _GEN_2774 : reservedValidList4_14; // @[decode.scala 400:29 323:31]
  wire  _GEN_3895 = 3'h3 == branchTracker ? _GEN_2775 : reservedValidList4_15; // @[decode.scala 400:29 323:31]
  wire  _GEN_3896 = 3'h3 == branchTracker ? _GEN_2776 : reservedValidList4_16; // @[decode.scala 400:29 323:31]
  wire  _GEN_3897 = 3'h3 == branchTracker ? _GEN_2777 : reservedValidList4_17; // @[decode.scala 400:29 323:31]
  wire  _GEN_3898 = 3'h3 == branchTracker ? _GEN_2778 : reservedValidList4_18; // @[decode.scala 400:29 323:31]
  wire  _GEN_3899 = 3'h3 == branchTracker ? _GEN_2779 : reservedValidList4_19; // @[decode.scala 400:29 323:31]
  wire  _GEN_3900 = 3'h3 == branchTracker ? _GEN_2780 : reservedValidList4_20; // @[decode.scala 400:29 323:31]
  wire  _GEN_3901 = 3'h3 == branchTracker ? _GEN_2781 : reservedValidList4_21; // @[decode.scala 400:29 323:31]
  wire  _GEN_3902 = 3'h3 == branchTracker ? _GEN_2782 : reservedValidList4_22; // @[decode.scala 400:29 323:31]
  wire  _GEN_3903 = 3'h3 == branchTracker ? _GEN_2783 : reservedValidList4_23; // @[decode.scala 400:29 323:31]
  wire  _GEN_3904 = 3'h3 == branchTracker ? _GEN_2784 : reservedValidList4_24; // @[decode.scala 400:29 323:31]
  wire  _GEN_3905 = 3'h3 == branchTracker ? _GEN_2785 : reservedValidList4_25; // @[decode.scala 400:29 323:31]
  wire  _GEN_3906 = 3'h3 == branchTracker ? _GEN_2786 : reservedValidList4_26; // @[decode.scala 400:29 323:31]
  wire  _GEN_3907 = 3'h3 == branchTracker ? _GEN_2787 : reservedValidList4_27; // @[decode.scala 400:29 323:31]
  wire  _GEN_3908 = 3'h3 == branchTracker ? _GEN_2788 : reservedValidList4_28; // @[decode.scala 400:29 323:31]
  wire  _GEN_3909 = 3'h3 == branchTracker ? _GEN_2789 : reservedValidList4_29; // @[decode.scala 400:29 323:31]
  wire  _GEN_3910 = 3'h3 == branchTracker ? _GEN_2790 : reservedValidList4_30; // @[decode.scala 400:29 323:31]
  wire  _GEN_3911 = 3'h3 == branchTracker ? _GEN_2791 : reservedValidList4_31; // @[decode.scala 400:29 323:31]
  wire  _GEN_3912 = 3'h3 == branchTracker ? _GEN_2792 : reservedValidList4_32; // @[decode.scala 400:29 323:31]
  wire  _GEN_3913 = 3'h3 == branchTracker ? _GEN_2793 : reservedValidList4_33; // @[decode.scala 400:29 323:31]
  wire  _GEN_3914 = 3'h3 == branchTracker ? _GEN_2794 : reservedValidList4_34; // @[decode.scala 400:29 323:31]
  wire  _GEN_3915 = 3'h3 == branchTracker ? _GEN_2795 : reservedValidList4_35; // @[decode.scala 400:29 323:31]
  wire  _GEN_3916 = 3'h3 == branchTracker ? _GEN_2796 : reservedValidList4_36; // @[decode.scala 400:29 323:31]
  wire  _GEN_3917 = 3'h3 == branchTracker ? _GEN_2797 : reservedValidList4_37; // @[decode.scala 400:29 323:31]
  wire  _GEN_3918 = 3'h3 == branchTracker ? _GEN_2798 : reservedValidList4_38; // @[decode.scala 400:29 323:31]
  wire  _GEN_3919 = 3'h3 == branchTracker ? _GEN_2799 : reservedValidList4_39; // @[decode.scala 400:29 323:31]
  wire  _GEN_3920 = 3'h3 == branchTracker ? _GEN_2800 : reservedValidList4_40; // @[decode.scala 400:29 323:31]
  wire  _GEN_3921 = 3'h3 == branchTracker ? _GEN_2801 : reservedValidList4_41; // @[decode.scala 400:29 323:31]
  wire  _GEN_3922 = 3'h3 == branchTracker ? _GEN_2802 : reservedValidList4_42; // @[decode.scala 400:29 323:31]
  wire  _GEN_3923 = 3'h3 == branchTracker ? _GEN_2803 : reservedValidList4_43; // @[decode.scala 400:29 323:31]
  wire  _GEN_3924 = 3'h3 == branchTracker ? _GEN_2804 : reservedValidList4_44; // @[decode.scala 400:29 323:31]
  wire  _GEN_3925 = 3'h3 == branchTracker ? _GEN_2805 : reservedValidList4_45; // @[decode.scala 400:29 323:31]
  wire  _GEN_3926 = 3'h3 == branchTracker ? _GEN_2806 : reservedValidList4_46; // @[decode.scala 400:29 323:31]
  wire  _GEN_3927 = 3'h3 == branchTracker ? _GEN_2807 : reservedValidList4_47; // @[decode.scala 400:29 323:31]
  wire  _GEN_3928 = 3'h3 == branchTracker ? _GEN_2808 : reservedValidList4_48; // @[decode.scala 400:29 323:31]
  wire  _GEN_3929 = 3'h3 == branchTracker ? _GEN_2809 : reservedValidList4_49; // @[decode.scala 400:29 323:31]
  wire  _GEN_3930 = 3'h3 == branchTracker ? _GEN_2810 : reservedValidList4_50; // @[decode.scala 400:29 323:31]
  wire  _GEN_3931 = 3'h3 == branchTracker ? _GEN_2811 : reservedValidList4_51; // @[decode.scala 400:29 323:31]
  wire  _GEN_3932 = 3'h3 == branchTracker ? _GEN_2812 : reservedValidList4_52; // @[decode.scala 400:29 323:31]
  wire  _GEN_3933 = 3'h3 == branchTracker ? _GEN_2813 : reservedValidList4_53; // @[decode.scala 400:29 323:31]
  wire  _GEN_3934 = 3'h3 == branchTracker ? _GEN_2814 : reservedValidList4_54; // @[decode.scala 400:29 323:31]
  wire  _GEN_3935 = 3'h3 == branchTracker ? _GEN_2815 : reservedValidList4_55; // @[decode.scala 400:29 323:31]
  wire  _GEN_3936 = 3'h3 == branchTracker ? _GEN_2816 : reservedValidList4_56; // @[decode.scala 400:29 323:31]
  wire  _GEN_3937 = 3'h3 == branchTracker ? _GEN_2817 : reservedValidList4_57; // @[decode.scala 400:29 323:31]
  wire  _GEN_3938 = 3'h3 == branchTracker ? _GEN_2818 : reservedValidList4_58; // @[decode.scala 400:29 323:31]
  wire  _GEN_3939 = 3'h3 == branchTracker ? _GEN_2819 : reservedValidList4_59; // @[decode.scala 400:29 323:31]
  wire  _GEN_3940 = 3'h3 == branchTracker ? _GEN_2820 : reservedValidList4_60; // @[decode.scala 400:29 323:31]
  wire  _GEN_3941 = 3'h3 == branchTracker ? _GEN_2821 : reservedValidList4_61; // @[decode.scala 400:29 323:31]
  wire  _GEN_3942 = 3'h3 == branchTracker ? _GEN_2822 : reservedValidList4_62; // @[decode.scala 400:29 323:31]
  wire  _GEN_3943 = 3'h3 == branchTracker ? _GEN_2823 : reservedValidList4_63; // @[decode.scala 400:29 323:31]
  wire [5:0] _GEN_3944 = 3'h2 == branchTracker ? _GEN_2664 : _GEN_2080; // @[decode.scala 400:29]
  wire [5:0] _GEN_3945 = 3'h2 == branchTracker ? _GEN_2665 : _GEN_2081; // @[decode.scala 400:29]
  wire [5:0] _GEN_3946 = 3'h2 == branchTracker ? _GEN_2666 : _GEN_2082; // @[decode.scala 400:29]
  wire [5:0] _GEN_3947 = 3'h2 == branchTracker ? _GEN_2667 : _GEN_2083; // @[decode.scala 400:29]
  wire [5:0] _GEN_3948 = 3'h2 == branchTracker ? _GEN_2668 : _GEN_2084; // @[decode.scala 400:29]
  wire [5:0] _GEN_3949 = 3'h2 == branchTracker ? _GEN_2669 : _GEN_2085; // @[decode.scala 400:29]
  wire [5:0] _GEN_3950 = 3'h2 == branchTracker ? _GEN_2670 : _GEN_2086; // @[decode.scala 400:29]
  wire [5:0] _GEN_3951 = 3'h2 == branchTracker ? _GEN_2671 : _GEN_2087; // @[decode.scala 400:29]
  wire [5:0] _GEN_3952 = 3'h2 == branchTracker ? _GEN_2672 : _GEN_2088; // @[decode.scala 400:29]
  wire [5:0] _GEN_3953 = 3'h2 == branchTracker ? _GEN_2673 : _GEN_2089; // @[decode.scala 400:29]
  wire [5:0] _GEN_3954 = 3'h2 == branchTracker ? _GEN_2674 : _GEN_2090; // @[decode.scala 400:29]
  wire [5:0] _GEN_3955 = 3'h2 == branchTracker ? _GEN_2675 : _GEN_2091; // @[decode.scala 400:29]
  wire [5:0] _GEN_3956 = 3'h2 == branchTracker ? _GEN_2676 : _GEN_2092; // @[decode.scala 400:29]
  wire [5:0] _GEN_3957 = 3'h2 == branchTracker ? _GEN_2677 : _GEN_2093; // @[decode.scala 400:29]
  wire [5:0] _GEN_3958 = 3'h2 == branchTracker ? _GEN_2678 : _GEN_2094; // @[decode.scala 400:29]
  wire [5:0] _GEN_3959 = 3'h2 == branchTracker ? _GEN_2679 : _GEN_2095; // @[decode.scala 400:29]
  wire [5:0] _GEN_3960 = 3'h2 == branchTracker ? _GEN_2680 : _GEN_2096; // @[decode.scala 400:29]
  wire [5:0] _GEN_3961 = 3'h2 == branchTracker ? _GEN_2681 : _GEN_2097; // @[decode.scala 400:29]
  wire [5:0] _GEN_3962 = 3'h2 == branchTracker ? _GEN_2682 : _GEN_2098; // @[decode.scala 400:29]
  wire [5:0] _GEN_3963 = 3'h2 == branchTracker ? _GEN_2683 : _GEN_2099; // @[decode.scala 400:29]
  wire [5:0] _GEN_3964 = 3'h2 == branchTracker ? _GEN_2684 : _GEN_2100; // @[decode.scala 400:29]
  wire [5:0] _GEN_3965 = 3'h2 == branchTracker ? _GEN_2685 : _GEN_2101; // @[decode.scala 400:29]
  wire [5:0] _GEN_3966 = 3'h2 == branchTracker ? _GEN_2686 : _GEN_2102; // @[decode.scala 400:29]
  wire [5:0] _GEN_3967 = 3'h2 == branchTracker ? _GEN_2687 : _GEN_2103; // @[decode.scala 400:29]
  wire [5:0] _GEN_3968 = 3'h2 == branchTracker ? _GEN_2688 : _GEN_2104; // @[decode.scala 400:29]
  wire [5:0] _GEN_3969 = 3'h2 == branchTracker ? _GEN_2689 : _GEN_2105; // @[decode.scala 400:29]
  wire [5:0] _GEN_3970 = 3'h2 == branchTracker ? _GEN_2690 : _GEN_2106; // @[decode.scala 400:29]
  wire [5:0] _GEN_3971 = 3'h2 == branchTracker ? _GEN_2691 : _GEN_2107; // @[decode.scala 400:29]
  wire [5:0] _GEN_3972 = 3'h2 == branchTracker ? _GEN_2692 : _GEN_2108; // @[decode.scala 400:29]
  wire [5:0] _GEN_3973 = 3'h2 == branchTracker ? _GEN_2693 : _GEN_2109; // @[decode.scala 400:29]
  wire [5:0] _GEN_3974 = 3'h2 == branchTracker ? _GEN_2694 : _GEN_2110; // @[decode.scala 400:29]
  wire [5:0] _GEN_3975 = 3'h2 == branchTracker ? _GEN_2695 : _GEN_2111; // @[decode.scala 400:29]
  wire  _GEN_3976 = 3'h2 == branchTracker ? _GEN_2696 : _GEN_2240; // @[decode.scala 400:29]
  wire  _GEN_3977 = 3'h2 == branchTracker ? _GEN_2697 : _GEN_2241; // @[decode.scala 400:29]
  wire  _GEN_3978 = 3'h2 == branchTracker ? _GEN_2698 : _GEN_2242; // @[decode.scala 400:29]
  wire  _GEN_3979 = 3'h2 == branchTracker ? _GEN_2699 : _GEN_2243; // @[decode.scala 400:29]
  wire  _GEN_3980 = 3'h2 == branchTracker ? _GEN_2700 : _GEN_2244; // @[decode.scala 400:29]
  wire  _GEN_3981 = 3'h2 == branchTracker ? _GEN_2701 : _GEN_2245; // @[decode.scala 400:29]
  wire  _GEN_3982 = 3'h2 == branchTracker ? _GEN_2702 : _GEN_2246; // @[decode.scala 400:29]
  wire  _GEN_3983 = 3'h2 == branchTracker ? _GEN_2703 : _GEN_2247; // @[decode.scala 400:29]
  wire  _GEN_3984 = 3'h2 == branchTracker ? _GEN_2704 : _GEN_2248; // @[decode.scala 400:29]
  wire  _GEN_3985 = 3'h2 == branchTracker ? _GEN_2705 : _GEN_2249; // @[decode.scala 400:29]
  wire  _GEN_3986 = 3'h2 == branchTracker ? _GEN_2706 : _GEN_2250; // @[decode.scala 400:29]
  wire  _GEN_3987 = 3'h2 == branchTracker ? _GEN_2707 : _GEN_2251; // @[decode.scala 400:29]
  wire  _GEN_3988 = 3'h2 == branchTracker ? _GEN_2708 : _GEN_2252; // @[decode.scala 400:29]
  wire  _GEN_3989 = 3'h2 == branchTracker ? _GEN_2709 : _GEN_2253; // @[decode.scala 400:29]
  wire  _GEN_3990 = 3'h2 == branchTracker ? _GEN_2710 : _GEN_2254; // @[decode.scala 400:29]
  wire  _GEN_3991 = 3'h2 == branchTracker ? _GEN_2711 : _GEN_2255; // @[decode.scala 400:29]
  wire  _GEN_3992 = 3'h2 == branchTracker ? _GEN_2712 : _GEN_2256; // @[decode.scala 400:29]
  wire  _GEN_3993 = 3'h2 == branchTracker ? _GEN_2713 : _GEN_2257; // @[decode.scala 400:29]
  wire  _GEN_3994 = 3'h2 == branchTracker ? _GEN_2714 : _GEN_2258; // @[decode.scala 400:29]
  wire  _GEN_3995 = 3'h2 == branchTracker ? _GEN_2715 : _GEN_2259; // @[decode.scala 400:29]
  wire  _GEN_3996 = 3'h2 == branchTracker ? _GEN_2716 : _GEN_2260; // @[decode.scala 400:29]
  wire  _GEN_3997 = 3'h2 == branchTracker ? _GEN_2717 : _GEN_2261; // @[decode.scala 400:29]
  wire  _GEN_3998 = 3'h2 == branchTracker ? _GEN_2718 : _GEN_2262; // @[decode.scala 400:29]
  wire  _GEN_3999 = 3'h2 == branchTracker ? _GEN_2719 : _GEN_2263; // @[decode.scala 400:29]
  wire  _GEN_4000 = 3'h2 == branchTracker ? _GEN_2720 : _GEN_2264; // @[decode.scala 400:29]
  wire  _GEN_4001 = 3'h2 == branchTracker ? _GEN_2721 : _GEN_2265; // @[decode.scala 400:29]
  wire  _GEN_4002 = 3'h2 == branchTracker ? _GEN_2722 : _GEN_2266; // @[decode.scala 400:29]
  wire  _GEN_4003 = 3'h2 == branchTracker ? _GEN_2723 : _GEN_2267; // @[decode.scala 400:29]
  wire  _GEN_4004 = 3'h2 == branchTracker ? _GEN_2724 : _GEN_2268; // @[decode.scala 400:29]
  wire  _GEN_4005 = 3'h2 == branchTracker ? _GEN_2725 : _GEN_2269; // @[decode.scala 400:29]
  wire  _GEN_4006 = 3'h2 == branchTracker ? _GEN_2726 : _GEN_2270; // @[decode.scala 400:29]
  wire  _GEN_4007 = 3'h2 == branchTracker ? _GEN_2727 : _GEN_2271; // @[decode.scala 400:29]
  wire  _GEN_4008 = 3'h2 == branchTracker ? _GEN_2728 : _GEN_2272; // @[decode.scala 400:29]
  wire  _GEN_4009 = 3'h2 == branchTracker ? _GEN_2729 : _GEN_2273; // @[decode.scala 400:29]
  wire  _GEN_4010 = 3'h2 == branchTracker ? _GEN_2730 : _GEN_2274; // @[decode.scala 400:29]
  wire  _GEN_4011 = 3'h2 == branchTracker ? _GEN_2731 : _GEN_2275; // @[decode.scala 400:29]
  wire  _GEN_4012 = 3'h2 == branchTracker ? _GEN_2732 : _GEN_2276; // @[decode.scala 400:29]
  wire  _GEN_4013 = 3'h2 == branchTracker ? _GEN_2733 : _GEN_2277; // @[decode.scala 400:29]
  wire  _GEN_4014 = 3'h2 == branchTracker ? _GEN_2734 : _GEN_2278; // @[decode.scala 400:29]
  wire  _GEN_4015 = 3'h2 == branchTracker ? _GEN_2735 : _GEN_2279; // @[decode.scala 400:29]
  wire  _GEN_4016 = 3'h2 == branchTracker ? _GEN_2736 : _GEN_2280; // @[decode.scala 400:29]
  wire  _GEN_4017 = 3'h2 == branchTracker ? _GEN_2737 : _GEN_2281; // @[decode.scala 400:29]
  wire  _GEN_4018 = 3'h2 == branchTracker ? _GEN_2738 : _GEN_2282; // @[decode.scala 400:29]
  wire  _GEN_4019 = 3'h2 == branchTracker ? _GEN_2739 : _GEN_2283; // @[decode.scala 400:29]
  wire  _GEN_4020 = 3'h2 == branchTracker ? _GEN_2740 : _GEN_2284; // @[decode.scala 400:29]
  wire  _GEN_4021 = 3'h2 == branchTracker ? _GEN_2741 : _GEN_2285; // @[decode.scala 400:29]
  wire  _GEN_4022 = 3'h2 == branchTracker ? _GEN_2742 : _GEN_2286; // @[decode.scala 400:29]
  wire  _GEN_4023 = 3'h2 == branchTracker ? _GEN_2743 : _GEN_2287; // @[decode.scala 400:29]
  wire  _GEN_4024 = 3'h2 == branchTracker ? _GEN_2744 : _GEN_2288; // @[decode.scala 400:29]
  wire  _GEN_4025 = 3'h2 == branchTracker ? _GEN_2745 : _GEN_2289; // @[decode.scala 400:29]
  wire  _GEN_4026 = 3'h2 == branchTracker ? _GEN_2746 : _GEN_2290; // @[decode.scala 400:29]
  wire  _GEN_4027 = 3'h2 == branchTracker ? _GEN_2747 : _GEN_2291; // @[decode.scala 400:29]
  wire  _GEN_4028 = 3'h2 == branchTracker ? _GEN_2748 : _GEN_2292; // @[decode.scala 400:29]
  wire  _GEN_4029 = 3'h2 == branchTracker ? _GEN_2749 : _GEN_2293; // @[decode.scala 400:29]
  wire  _GEN_4030 = 3'h2 == branchTracker ? _GEN_2750 : _GEN_2294; // @[decode.scala 400:29]
  wire  _GEN_4031 = 3'h2 == branchTracker ? _GEN_2751 : _GEN_2295; // @[decode.scala 400:29]
  wire  _GEN_4032 = 3'h2 == branchTracker ? _GEN_2752 : _GEN_2296; // @[decode.scala 400:29]
  wire  _GEN_4033 = 3'h2 == branchTracker ? _GEN_2753 : _GEN_2297; // @[decode.scala 400:29]
  wire  _GEN_4034 = 3'h2 == branchTracker ? _GEN_2754 : _GEN_2298; // @[decode.scala 400:29]
  wire  _GEN_4035 = 3'h2 == branchTracker ? _GEN_2755 : _GEN_2299; // @[decode.scala 400:29]
  wire  _GEN_4036 = 3'h2 == branchTracker ? _GEN_2756 : _GEN_2300; // @[decode.scala 400:29]
  wire  _GEN_4037 = 3'h2 == branchTracker ? _GEN_2757 : _GEN_2301; // @[decode.scala 400:29]
  wire  _GEN_4038 = 3'h2 == branchTracker ? _GEN_2758 : _GEN_2302; // @[decode.scala 400:29]
  wire  _GEN_4040 = 3'h2 == branchTracker ? _GEN_2760 : _GEN_2432; // @[decode.scala 400:29]
  wire  _GEN_4041 = 3'h2 == branchTracker ? _GEN_2761 : _GEN_2433; // @[decode.scala 400:29]
  wire  _GEN_4042 = 3'h2 == branchTracker ? _GEN_2762 : _GEN_2434; // @[decode.scala 400:29]
  wire  _GEN_4043 = 3'h2 == branchTracker ? _GEN_2763 : _GEN_2435; // @[decode.scala 400:29]
  wire  _GEN_4044 = 3'h2 == branchTracker ? _GEN_2764 : _GEN_2436; // @[decode.scala 400:29]
  wire  _GEN_4045 = 3'h2 == branchTracker ? _GEN_2765 : _GEN_2437; // @[decode.scala 400:29]
  wire  _GEN_4046 = 3'h2 == branchTracker ? _GEN_2766 : _GEN_2438; // @[decode.scala 400:29]
  wire  _GEN_4047 = 3'h2 == branchTracker ? _GEN_2767 : _GEN_2439; // @[decode.scala 400:29]
  wire  _GEN_4048 = 3'h2 == branchTracker ? _GEN_2768 : _GEN_2440; // @[decode.scala 400:29]
  wire  _GEN_4049 = 3'h2 == branchTracker ? _GEN_2769 : _GEN_2441; // @[decode.scala 400:29]
  wire  _GEN_4050 = 3'h2 == branchTracker ? _GEN_2770 : _GEN_2442; // @[decode.scala 400:29]
  wire  _GEN_4051 = 3'h2 == branchTracker ? _GEN_2771 : _GEN_2443; // @[decode.scala 400:29]
  wire  _GEN_4052 = 3'h2 == branchTracker ? _GEN_2772 : _GEN_2444; // @[decode.scala 400:29]
  wire  _GEN_4053 = 3'h2 == branchTracker ? _GEN_2773 : _GEN_2445; // @[decode.scala 400:29]
  wire  _GEN_4054 = 3'h2 == branchTracker ? _GEN_2774 : _GEN_2446; // @[decode.scala 400:29]
  wire  _GEN_4055 = 3'h2 == branchTracker ? _GEN_2775 : _GEN_2447; // @[decode.scala 400:29]
  wire  _GEN_4056 = 3'h2 == branchTracker ? _GEN_2776 : _GEN_2448; // @[decode.scala 400:29]
  wire  _GEN_4057 = 3'h2 == branchTracker ? _GEN_2777 : _GEN_2449; // @[decode.scala 400:29]
  wire  _GEN_4058 = 3'h2 == branchTracker ? _GEN_2778 : _GEN_2450; // @[decode.scala 400:29]
  wire  _GEN_4059 = 3'h2 == branchTracker ? _GEN_2779 : _GEN_2451; // @[decode.scala 400:29]
  wire  _GEN_4060 = 3'h2 == branchTracker ? _GEN_2780 : _GEN_2452; // @[decode.scala 400:29]
  wire  _GEN_4061 = 3'h2 == branchTracker ? _GEN_2781 : _GEN_2453; // @[decode.scala 400:29]
  wire  _GEN_4062 = 3'h2 == branchTracker ? _GEN_2782 : _GEN_2454; // @[decode.scala 400:29]
  wire  _GEN_4063 = 3'h2 == branchTracker ? _GEN_2783 : _GEN_2455; // @[decode.scala 400:29]
  wire  _GEN_4064 = 3'h2 == branchTracker ? _GEN_2784 : _GEN_2456; // @[decode.scala 400:29]
  wire  _GEN_4065 = 3'h2 == branchTracker ? _GEN_2785 : _GEN_2457; // @[decode.scala 400:29]
  wire  _GEN_4066 = 3'h2 == branchTracker ? _GEN_2786 : _GEN_2458; // @[decode.scala 400:29]
  wire  _GEN_4067 = 3'h2 == branchTracker ? _GEN_2787 : _GEN_2459; // @[decode.scala 400:29]
  wire  _GEN_4068 = 3'h2 == branchTracker ? _GEN_2788 : _GEN_2460; // @[decode.scala 400:29]
  wire  _GEN_4069 = 3'h2 == branchTracker ? _GEN_2789 : _GEN_2461; // @[decode.scala 400:29]
  wire  _GEN_4070 = 3'h2 == branchTracker ? _GEN_2790 : _GEN_2462; // @[decode.scala 400:29]
  wire  _GEN_4071 = 3'h2 == branchTracker ? _GEN_2791 : _GEN_2463; // @[decode.scala 400:29]
  wire  _GEN_4072 = 3'h2 == branchTracker ? _GEN_2792 : _GEN_2464; // @[decode.scala 400:29]
  wire  _GEN_4073 = 3'h2 == branchTracker ? _GEN_2793 : _GEN_2465; // @[decode.scala 400:29]
  wire  _GEN_4074 = 3'h2 == branchTracker ? _GEN_2794 : _GEN_2466; // @[decode.scala 400:29]
  wire  _GEN_4075 = 3'h2 == branchTracker ? _GEN_2795 : _GEN_2467; // @[decode.scala 400:29]
  wire  _GEN_4076 = 3'h2 == branchTracker ? _GEN_2796 : _GEN_2468; // @[decode.scala 400:29]
  wire  _GEN_4077 = 3'h2 == branchTracker ? _GEN_2797 : _GEN_2469; // @[decode.scala 400:29]
  wire  _GEN_4078 = 3'h2 == branchTracker ? _GEN_2798 : _GEN_2470; // @[decode.scala 400:29]
  wire  _GEN_4079 = 3'h2 == branchTracker ? _GEN_2799 : _GEN_2471; // @[decode.scala 400:29]
  wire  _GEN_4080 = 3'h2 == branchTracker ? _GEN_2800 : _GEN_2472; // @[decode.scala 400:29]
  wire  _GEN_4081 = 3'h2 == branchTracker ? _GEN_2801 : _GEN_2473; // @[decode.scala 400:29]
  wire  _GEN_4082 = 3'h2 == branchTracker ? _GEN_2802 : _GEN_2474; // @[decode.scala 400:29]
  wire  _GEN_4083 = 3'h2 == branchTracker ? _GEN_2803 : _GEN_2475; // @[decode.scala 400:29]
  wire  _GEN_4084 = 3'h2 == branchTracker ? _GEN_2804 : _GEN_2476; // @[decode.scala 400:29]
  wire  _GEN_4085 = 3'h2 == branchTracker ? _GEN_2805 : _GEN_2477; // @[decode.scala 400:29]
  wire  _GEN_4086 = 3'h2 == branchTracker ? _GEN_2806 : _GEN_2478; // @[decode.scala 400:29]
  wire  _GEN_4087 = 3'h2 == branchTracker ? _GEN_2807 : _GEN_2479; // @[decode.scala 400:29]
  wire  _GEN_4088 = 3'h2 == branchTracker ? _GEN_2808 : _GEN_2480; // @[decode.scala 400:29]
  wire  _GEN_4089 = 3'h2 == branchTracker ? _GEN_2809 : _GEN_2481; // @[decode.scala 400:29]
  wire  _GEN_4090 = 3'h2 == branchTracker ? _GEN_2810 : _GEN_2482; // @[decode.scala 400:29]
  wire  _GEN_4091 = 3'h2 == branchTracker ? _GEN_2811 : _GEN_2483; // @[decode.scala 400:29]
  wire  _GEN_4092 = 3'h2 == branchTracker ? _GEN_2812 : _GEN_2484; // @[decode.scala 400:29]
  wire  _GEN_4093 = 3'h2 == branchTracker ? _GEN_2813 : _GEN_2485; // @[decode.scala 400:29]
  wire  _GEN_4094 = 3'h2 == branchTracker ? _GEN_2814 : _GEN_2486; // @[decode.scala 400:29]
  wire  _GEN_4095 = 3'h2 == branchTracker ? _GEN_2815 : _GEN_2487; // @[decode.scala 400:29]
  wire  _GEN_4096 = 3'h2 == branchTracker ? _GEN_2816 : _GEN_2488; // @[decode.scala 400:29]
  wire  _GEN_4097 = 3'h2 == branchTracker ? _GEN_2817 : _GEN_2489; // @[decode.scala 400:29]
  wire  _GEN_4098 = 3'h2 == branchTracker ? _GEN_2818 : _GEN_2490; // @[decode.scala 400:29]
  wire  _GEN_4099 = 3'h2 == branchTracker ? _GEN_2819 : _GEN_2491; // @[decode.scala 400:29]
  wire  _GEN_4100 = 3'h2 == branchTracker ? _GEN_2820 : _GEN_2492; // @[decode.scala 400:29]
  wire  _GEN_4101 = 3'h2 == branchTracker ? _GEN_2821 : _GEN_2493; // @[decode.scala 400:29]
  wire  _GEN_4102 = 3'h2 == branchTracker ? _GEN_2822 : _GEN_2494; // @[decode.scala 400:29]
  wire  _GEN_4103 = 3'h2 == branchTracker ? _GEN_2823 : _GEN_2495; // @[decode.scala 400:29]
  wire [5:0] _GEN_4104 = 3'h2 == branchTracker ? reservedRegMap4_0 : _GEN_3784; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4105 = 3'h2 == branchTracker ? reservedRegMap4_1 : _GEN_3785; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4106 = 3'h2 == branchTracker ? reservedRegMap4_2 : _GEN_3786; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4107 = 3'h2 == branchTracker ? reservedRegMap4_3 : _GEN_3787; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4108 = 3'h2 == branchTracker ? reservedRegMap4_4 : _GEN_3788; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4109 = 3'h2 == branchTracker ? reservedRegMap4_5 : _GEN_3789; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4110 = 3'h2 == branchTracker ? reservedRegMap4_6 : _GEN_3790; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4111 = 3'h2 == branchTracker ? reservedRegMap4_7 : _GEN_3791; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4112 = 3'h2 == branchTracker ? reservedRegMap4_8 : _GEN_3792; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4113 = 3'h2 == branchTracker ? reservedRegMap4_9 : _GEN_3793; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4114 = 3'h2 == branchTracker ? reservedRegMap4_10 : _GEN_3794; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4115 = 3'h2 == branchTracker ? reservedRegMap4_11 : _GEN_3795; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4116 = 3'h2 == branchTracker ? reservedRegMap4_12 : _GEN_3796; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4117 = 3'h2 == branchTracker ? reservedRegMap4_13 : _GEN_3797; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4118 = 3'h2 == branchTracker ? reservedRegMap4_14 : _GEN_3798; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4119 = 3'h2 == branchTracker ? reservedRegMap4_15 : _GEN_3799; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4120 = 3'h2 == branchTracker ? reservedRegMap4_16 : _GEN_3800; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4121 = 3'h2 == branchTracker ? reservedRegMap4_17 : _GEN_3801; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4122 = 3'h2 == branchTracker ? reservedRegMap4_18 : _GEN_3802; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4123 = 3'h2 == branchTracker ? reservedRegMap4_19 : _GEN_3803; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4124 = 3'h2 == branchTracker ? reservedRegMap4_20 : _GEN_3804; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4125 = 3'h2 == branchTracker ? reservedRegMap4_21 : _GEN_3805; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4126 = 3'h2 == branchTracker ? reservedRegMap4_22 : _GEN_3806; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4127 = 3'h2 == branchTracker ? reservedRegMap4_23 : _GEN_3807; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4128 = 3'h2 == branchTracker ? reservedRegMap4_24 : _GEN_3808; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4129 = 3'h2 == branchTracker ? reservedRegMap4_25 : _GEN_3809; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4130 = 3'h2 == branchTracker ? reservedRegMap4_26 : _GEN_3810; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4131 = 3'h2 == branchTracker ? reservedRegMap4_27 : _GEN_3811; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4132 = 3'h2 == branchTracker ? reservedRegMap4_28 : _GEN_3812; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4133 = 3'h2 == branchTracker ? reservedRegMap4_29 : _GEN_3813; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4134 = 3'h2 == branchTracker ? reservedRegMap4_30 : _GEN_3814; // @[decode.scala 313:28 400:29]
  wire [5:0] _GEN_4135 = 3'h2 == branchTracker ? reservedRegMap4_31 : _GEN_3815; // @[decode.scala 313:28 400:29]
  wire  _GEN_4136 = 3'h2 == branchTracker ? reservedFreeList4_0 : _GEN_3816; // @[decode.scala 400:29 318:30]
  wire  _GEN_4137 = 3'h2 == branchTracker ? reservedFreeList4_1 : _GEN_3817; // @[decode.scala 400:29 318:30]
  wire  _GEN_4138 = 3'h2 == branchTracker ? reservedFreeList4_2 : _GEN_3818; // @[decode.scala 400:29 318:30]
  wire  _GEN_4139 = 3'h2 == branchTracker ? reservedFreeList4_3 : _GEN_3819; // @[decode.scala 400:29 318:30]
  wire  _GEN_4140 = 3'h2 == branchTracker ? reservedFreeList4_4 : _GEN_3820; // @[decode.scala 400:29 318:30]
  wire  _GEN_4141 = 3'h2 == branchTracker ? reservedFreeList4_5 : _GEN_3821; // @[decode.scala 400:29 318:30]
  wire  _GEN_4142 = 3'h2 == branchTracker ? reservedFreeList4_6 : _GEN_3822; // @[decode.scala 400:29 318:30]
  wire  _GEN_4143 = 3'h2 == branchTracker ? reservedFreeList4_7 : _GEN_3823; // @[decode.scala 400:29 318:30]
  wire  _GEN_4144 = 3'h2 == branchTracker ? reservedFreeList4_8 : _GEN_3824; // @[decode.scala 400:29 318:30]
  wire  _GEN_4145 = 3'h2 == branchTracker ? reservedFreeList4_9 : _GEN_3825; // @[decode.scala 400:29 318:30]
  wire  _GEN_4146 = 3'h2 == branchTracker ? reservedFreeList4_10 : _GEN_3826; // @[decode.scala 400:29 318:30]
  wire  _GEN_4147 = 3'h2 == branchTracker ? reservedFreeList4_11 : _GEN_3827; // @[decode.scala 400:29 318:30]
  wire  _GEN_4148 = 3'h2 == branchTracker ? reservedFreeList4_12 : _GEN_3828; // @[decode.scala 400:29 318:30]
  wire  _GEN_4149 = 3'h2 == branchTracker ? reservedFreeList4_13 : _GEN_3829; // @[decode.scala 400:29 318:30]
  wire  _GEN_4150 = 3'h2 == branchTracker ? reservedFreeList4_14 : _GEN_3830; // @[decode.scala 400:29 318:30]
  wire  _GEN_4151 = 3'h2 == branchTracker ? reservedFreeList4_15 : _GEN_3831; // @[decode.scala 400:29 318:30]
  wire  _GEN_4152 = 3'h2 == branchTracker ? reservedFreeList4_16 : _GEN_3832; // @[decode.scala 400:29 318:30]
  wire  _GEN_4153 = 3'h2 == branchTracker ? reservedFreeList4_17 : _GEN_3833; // @[decode.scala 400:29 318:30]
  wire  _GEN_4154 = 3'h2 == branchTracker ? reservedFreeList4_18 : _GEN_3834; // @[decode.scala 400:29 318:30]
  wire  _GEN_4155 = 3'h2 == branchTracker ? reservedFreeList4_19 : _GEN_3835; // @[decode.scala 400:29 318:30]
  wire  _GEN_4156 = 3'h2 == branchTracker ? reservedFreeList4_20 : _GEN_3836; // @[decode.scala 400:29 318:30]
  wire  _GEN_4157 = 3'h2 == branchTracker ? reservedFreeList4_21 : _GEN_3837; // @[decode.scala 400:29 318:30]
  wire  _GEN_4158 = 3'h2 == branchTracker ? reservedFreeList4_22 : _GEN_3838; // @[decode.scala 400:29 318:30]
  wire  _GEN_4159 = 3'h2 == branchTracker ? reservedFreeList4_23 : _GEN_3839; // @[decode.scala 400:29 318:30]
  wire  _GEN_4160 = 3'h2 == branchTracker ? reservedFreeList4_24 : _GEN_3840; // @[decode.scala 400:29 318:30]
  wire  _GEN_4161 = 3'h2 == branchTracker ? reservedFreeList4_25 : _GEN_3841; // @[decode.scala 400:29 318:30]
  wire  _GEN_4162 = 3'h2 == branchTracker ? reservedFreeList4_26 : _GEN_3842; // @[decode.scala 400:29 318:30]
  wire  _GEN_4163 = 3'h2 == branchTracker ? reservedFreeList4_27 : _GEN_3843; // @[decode.scala 400:29 318:30]
  wire  _GEN_4164 = 3'h2 == branchTracker ? reservedFreeList4_28 : _GEN_3844; // @[decode.scala 400:29 318:30]
  wire  _GEN_4165 = 3'h2 == branchTracker ? reservedFreeList4_29 : _GEN_3845; // @[decode.scala 400:29 318:30]
  wire  _GEN_4166 = 3'h2 == branchTracker ? reservedFreeList4_30 : _GEN_3846; // @[decode.scala 400:29 318:30]
  wire  _GEN_4167 = 3'h2 == branchTracker ? reservedFreeList4_31 : _GEN_3847; // @[decode.scala 400:29 318:30]
  wire  _GEN_4168 = 3'h2 == branchTracker ? reservedFreeList4_32 : _GEN_3848; // @[decode.scala 400:29 318:30]
  wire  _GEN_4169 = 3'h2 == branchTracker ? reservedFreeList4_33 : _GEN_3849; // @[decode.scala 400:29 318:30]
  wire  _GEN_4170 = 3'h2 == branchTracker ? reservedFreeList4_34 : _GEN_3850; // @[decode.scala 400:29 318:30]
  wire  _GEN_4171 = 3'h2 == branchTracker ? reservedFreeList4_35 : _GEN_3851; // @[decode.scala 400:29 318:30]
  wire  _GEN_4172 = 3'h2 == branchTracker ? reservedFreeList4_36 : _GEN_3852; // @[decode.scala 400:29 318:30]
  wire  _GEN_4173 = 3'h2 == branchTracker ? reservedFreeList4_37 : _GEN_3853; // @[decode.scala 400:29 318:30]
  wire  _GEN_4174 = 3'h2 == branchTracker ? reservedFreeList4_38 : _GEN_3854; // @[decode.scala 400:29 318:30]
  wire  _GEN_4175 = 3'h2 == branchTracker ? reservedFreeList4_39 : _GEN_3855; // @[decode.scala 400:29 318:30]
  wire  _GEN_4176 = 3'h2 == branchTracker ? reservedFreeList4_40 : _GEN_3856; // @[decode.scala 400:29 318:30]
  wire  _GEN_4177 = 3'h2 == branchTracker ? reservedFreeList4_41 : _GEN_3857; // @[decode.scala 400:29 318:30]
  wire  _GEN_4178 = 3'h2 == branchTracker ? reservedFreeList4_42 : _GEN_3858; // @[decode.scala 400:29 318:30]
  wire  _GEN_4179 = 3'h2 == branchTracker ? reservedFreeList4_43 : _GEN_3859; // @[decode.scala 400:29 318:30]
  wire  _GEN_4180 = 3'h2 == branchTracker ? reservedFreeList4_44 : _GEN_3860; // @[decode.scala 400:29 318:30]
  wire  _GEN_4181 = 3'h2 == branchTracker ? reservedFreeList4_45 : _GEN_3861; // @[decode.scala 400:29 318:30]
  wire  _GEN_4182 = 3'h2 == branchTracker ? reservedFreeList4_46 : _GEN_3862; // @[decode.scala 400:29 318:30]
  wire  _GEN_4183 = 3'h2 == branchTracker ? reservedFreeList4_47 : _GEN_3863; // @[decode.scala 400:29 318:30]
  wire  _GEN_4184 = 3'h2 == branchTracker ? reservedFreeList4_48 : _GEN_3864; // @[decode.scala 400:29 318:30]
  wire  _GEN_4185 = 3'h2 == branchTracker ? reservedFreeList4_49 : _GEN_3865; // @[decode.scala 400:29 318:30]
  wire  _GEN_4186 = 3'h2 == branchTracker ? reservedFreeList4_50 : _GEN_3866; // @[decode.scala 400:29 318:30]
  wire  _GEN_4187 = 3'h2 == branchTracker ? reservedFreeList4_51 : _GEN_3867; // @[decode.scala 400:29 318:30]
  wire  _GEN_4188 = 3'h2 == branchTracker ? reservedFreeList4_52 : _GEN_3868; // @[decode.scala 400:29 318:30]
  wire  _GEN_4189 = 3'h2 == branchTracker ? reservedFreeList4_53 : _GEN_3869; // @[decode.scala 400:29 318:30]
  wire  _GEN_4190 = 3'h2 == branchTracker ? reservedFreeList4_54 : _GEN_3870; // @[decode.scala 400:29 318:30]
  wire  _GEN_4191 = 3'h2 == branchTracker ? reservedFreeList4_55 : _GEN_3871; // @[decode.scala 400:29 318:30]
  wire  _GEN_4192 = 3'h2 == branchTracker ? reservedFreeList4_56 : _GEN_3872; // @[decode.scala 400:29 318:30]
  wire  _GEN_4193 = 3'h2 == branchTracker ? reservedFreeList4_57 : _GEN_3873; // @[decode.scala 400:29 318:30]
  wire  _GEN_4194 = 3'h2 == branchTracker ? reservedFreeList4_58 : _GEN_3874; // @[decode.scala 400:29 318:30]
  wire  _GEN_4195 = 3'h2 == branchTracker ? reservedFreeList4_59 : _GEN_3875; // @[decode.scala 400:29 318:30]
  wire  _GEN_4196 = 3'h2 == branchTracker ? reservedFreeList4_60 : _GEN_3876; // @[decode.scala 400:29 318:30]
  wire  _GEN_4197 = 3'h2 == branchTracker ? reservedFreeList4_61 : _GEN_3877; // @[decode.scala 400:29 318:30]
  wire  _GEN_4198 = 3'h2 == branchTracker ? reservedFreeList4_62 : _GEN_3878; // @[decode.scala 400:29 318:30]
  wire  _GEN_4200 = 3'h2 == branchTracker ? reservedValidList4_0 : _GEN_3880; // @[decode.scala 400:29 323:31]
  wire  _GEN_4201 = 3'h2 == branchTracker ? reservedValidList4_1 : _GEN_3881; // @[decode.scala 400:29 323:31]
  wire  _GEN_4202 = 3'h2 == branchTracker ? reservedValidList4_2 : _GEN_3882; // @[decode.scala 400:29 323:31]
  wire  _GEN_4203 = 3'h2 == branchTracker ? reservedValidList4_3 : _GEN_3883; // @[decode.scala 400:29 323:31]
  wire  _GEN_4204 = 3'h2 == branchTracker ? reservedValidList4_4 : _GEN_3884; // @[decode.scala 400:29 323:31]
  wire  _GEN_4205 = 3'h2 == branchTracker ? reservedValidList4_5 : _GEN_3885; // @[decode.scala 400:29 323:31]
  wire  _GEN_4206 = 3'h2 == branchTracker ? reservedValidList4_6 : _GEN_3886; // @[decode.scala 400:29 323:31]
  wire  _GEN_4207 = 3'h2 == branchTracker ? reservedValidList4_7 : _GEN_3887; // @[decode.scala 400:29 323:31]
  wire  _GEN_4208 = 3'h2 == branchTracker ? reservedValidList4_8 : _GEN_3888; // @[decode.scala 400:29 323:31]
  wire  _GEN_4209 = 3'h2 == branchTracker ? reservedValidList4_9 : _GEN_3889; // @[decode.scala 400:29 323:31]
  wire  _GEN_4210 = 3'h2 == branchTracker ? reservedValidList4_10 : _GEN_3890; // @[decode.scala 400:29 323:31]
  wire  _GEN_4211 = 3'h2 == branchTracker ? reservedValidList4_11 : _GEN_3891; // @[decode.scala 400:29 323:31]
  wire  _GEN_4212 = 3'h2 == branchTracker ? reservedValidList4_12 : _GEN_3892; // @[decode.scala 400:29 323:31]
  wire  _GEN_4213 = 3'h2 == branchTracker ? reservedValidList4_13 : _GEN_3893; // @[decode.scala 400:29 323:31]
  wire  _GEN_4214 = 3'h2 == branchTracker ? reservedValidList4_14 : _GEN_3894; // @[decode.scala 400:29 323:31]
  wire  _GEN_4215 = 3'h2 == branchTracker ? reservedValidList4_15 : _GEN_3895; // @[decode.scala 400:29 323:31]
  wire  _GEN_4216 = 3'h2 == branchTracker ? reservedValidList4_16 : _GEN_3896; // @[decode.scala 400:29 323:31]
  wire  _GEN_4217 = 3'h2 == branchTracker ? reservedValidList4_17 : _GEN_3897; // @[decode.scala 400:29 323:31]
  wire  _GEN_4218 = 3'h2 == branchTracker ? reservedValidList4_18 : _GEN_3898; // @[decode.scala 400:29 323:31]
  wire  _GEN_4219 = 3'h2 == branchTracker ? reservedValidList4_19 : _GEN_3899; // @[decode.scala 400:29 323:31]
  wire  _GEN_4220 = 3'h2 == branchTracker ? reservedValidList4_20 : _GEN_3900; // @[decode.scala 400:29 323:31]
  wire  _GEN_4221 = 3'h2 == branchTracker ? reservedValidList4_21 : _GEN_3901; // @[decode.scala 400:29 323:31]
  wire  _GEN_4222 = 3'h2 == branchTracker ? reservedValidList4_22 : _GEN_3902; // @[decode.scala 400:29 323:31]
  wire  _GEN_4223 = 3'h2 == branchTracker ? reservedValidList4_23 : _GEN_3903; // @[decode.scala 400:29 323:31]
  wire  _GEN_4224 = 3'h2 == branchTracker ? reservedValidList4_24 : _GEN_3904; // @[decode.scala 400:29 323:31]
  wire  _GEN_4225 = 3'h2 == branchTracker ? reservedValidList4_25 : _GEN_3905; // @[decode.scala 400:29 323:31]
  wire  _GEN_4226 = 3'h2 == branchTracker ? reservedValidList4_26 : _GEN_3906; // @[decode.scala 400:29 323:31]
  wire  _GEN_4227 = 3'h2 == branchTracker ? reservedValidList4_27 : _GEN_3907; // @[decode.scala 400:29 323:31]
  wire  _GEN_4228 = 3'h2 == branchTracker ? reservedValidList4_28 : _GEN_3908; // @[decode.scala 400:29 323:31]
  wire  _GEN_4229 = 3'h2 == branchTracker ? reservedValidList4_29 : _GEN_3909; // @[decode.scala 400:29 323:31]
  wire  _GEN_4230 = 3'h2 == branchTracker ? reservedValidList4_30 : _GEN_3910; // @[decode.scala 400:29 323:31]
  wire  _GEN_4231 = 3'h2 == branchTracker ? reservedValidList4_31 : _GEN_3911; // @[decode.scala 400:29 323:31]
  wire  _GEN_4232 = 3'h2 == branchTracker ? reservedValidList4_32 : _GEN_3912; // @[decode.scala 400:29 323:31]
  wire  _GEN_4233 = 3'h2 == branchTracker ? reservedValidList4_33 : _GEN_3913; // @[decode.scala 400:29 323:31]
  wire  _GEN_4234 = 3'h2 == branchTracker ? reservedValidList4_34 : _GEN_3914; // @[decode.scala 400:29 323:31]
  wire  _GEN_4235 = 3'h2 == branchTracker ? reservedValidList4_35 : _GEN_3915; // @[decode.scala 400:29 323:31]
  wire  _GEN_4236 = 3'h2 == branchTracker ? reservedValidList4_36 : _GEN_3916; // @[decode.scala 400:29 323:31]
  wire  _GEN_4237 = 3'h2 == branchTracker ? reservedValidList4_37 : _GEN_3917; // @[decode.scala 400:29 323:31]
  wire  _GEN_4238 = 3'h2 == branchTracker ? reservedValidList4_38 : _GEN_3918; // @[decode.scala 400:29 323:31]
  wire  _GEN_4239 = 3'h2 == branchTracker ? reservedValidList4_39 : _GEN_3919; // @[decode.scala 400:29 323:31]
  wire  _GEN_4240 = 3'h2 == branchTracker ? reservedValidList4_40 : _GEN_3920; // @[decode.scala 400:29 323:31]
  wire  _GEN_4241 = 3'h2 == branchTracker ? reservedValidList4_41 : _GEN_3921; // @[decode.scala 400:29 323:31]
  wire  _GEN_4242 = 3'h2 == branchTracker ? reservedValidList4_42 : _GEN_3922; // @[decode.scala 400:29 323:31]
  wire  _GEN_4243 = 3'h2 == branchTracker ? reservedValidList4_43 : _GEN_3923; // @[decode.scala 400:29 323:31]
  wire  _GEN_4244 = 3'h2 == branchTracker ? reservedValidList4_44 : _GEN_3924; // @[decode.scala 400:29 323:31]
  wire  _GEN_4245 = 3'h2 == branchTracker ? reservedValidList4_45 : _GEN_3925; // @[decode.scala 400:29 323:31]
  wire  _GEN_4246 = 3'h2 == branchTracker ? reservedValidList4_46 : _GEN_3926; // @[decode.scala 400:29 323:31]
  wire  _GEN_4247 = 3'h2 == branchTracker ? reservedValidList4_47 : _GEN_3927; // @[decode.scala 400:29 323:31]
  wire  _GEN_4248 = 3'h2 == branchTracker ? reservedValidList4_48 : _GEN_3928; // @[decode.scala 400:29 323:31]
  wire  _GEN_4249 = 3'h2 == branchTracker ? reservedValidList4_49 : _GEN_3929; // @[decode.scala 400:29 323:31]
  wire  _GEN_4250 = 3'h2 == branchTracker ? reservedValidList4_50 : _GEN_3930; // @[decode.scala 400:29 323:31]
  wire  _GEN_4251 = 3'h2 == branchTracker ? reservedValidList4_51 : _GEN_3931; // @[decode.scala 400:29 323:31]
  wire  _GEN_4252 = 3'h2 == branchTracker ? reservedValidList4_52 : _GEN_3932; // @[decode.scala 400:29 323:31]
  wire  _GEN_4253 = 3'h2 == branchTracker ? reservedValidList4_53 : _GEN_3933; // @[decode.scala 400:29 323:31]
  wire  _GEN_4254 = 3'h2 == branchTracker ? reservedValidList4_54 : _GEN_3934; // @[decode.scala 400:29 323:31]
  wire  _GEN_4255 = 3'h2 == branchTracker ? reservedValidList4_55 : _GEN_3935; // @[decode.scala 400:29 323:31]
  wire  _GEN_4256 = 3'h2 == branchTracker ? reservedValidList4_56 : _GEN_3936; // @[decode.scala 400:29 323:31]
  wire  _GEN_4257 = 3'h2 == branchTracker ? reservedValidList4_57 : _GEN_3937; // @[decode.scala 400:29 323:31]
  wire  _GEN_4258 = 3'h2 == branchTracker ? reservedValidList4_58 : _GEN_3938; // @[decode.scala 400:29 323:31]
  wire  _GEN_4259 = 3'h2 == branchTracker ? reservedValidList4_59 : _GEN_3939; // @[decode.scala 400:29 323:31]
  wire  _GEN_4260 = 3'h2 == branchTracker ? reservedValidList4_60 : _GEN_3940; // @[decode.scala 400:29 323:31]
  wire  _GEN_4261 = 3'h2 == branchTracker ? reservedValidList4_61 : _GEN_3941; // @[decode.scala 400:29 323:31]
  wire  _GEN_4262 = 3'h2 == branchTracker ? reservedValidList4_62 : _GEN_3942; // @[decode.scala 400:29 323:31]
  wire  _GEN_4263 = 3'h2 == branchTracker ? reservedValidList4_63 : _GEN_3943; // @[decode.scala 400:29 323:31]
  wire  _GEN_4296 = 3'h1 == branchTracker ? _GEN_2696 : _GEN_2176; // @[decode.scala 400:29]
  wire  _GEN_4297 = 3'h1 == branchTracker ? _GEN_2697 : _GEN_2177; // @[decode.scala 400:29]
  wire  _GEN_4298 = 3'h1 == branchTracker ? _GEN_2698 : _GEN_2178; // @[decode.scala 400:29]
  wire  _GEN_4299 = 3'h1 == branchTracker ? _GEN_2699 : _GEN_2179; // @[decode.scala 400:29]
  wire  _GEN_4300 = 3'h1 == branchTracker ? _GEN_2700 : _GEN_2180; // @[decode.scala 400:29]
  wire  _GEN_4301 = 3'h1 == branchTracker ? _GEN_2701 : _GEN_2181; // @[decode.scala 400:29]
  wire  _GEN_4302 = 3'h1 == branchTracker ? _GEN_2702 : _GEN_2182; // @[decode.scala 400:29]
  wire  _GEN_4303 = 3'h1 == branchTracker ? _GEN_2703 : _GEN_2183; // @[decode.scala 400:29]
  wire  _GEN_4304 = 3'h1 == branchTracker ? _GEN_2704 : _GEN_2184; // @[decode.scala 400:29]
  wire  _GEN_4305 = 3'h1 == branchTracker ? _GEN_2705 : _GEN_2185; // @[decode.scala 400:29]
  wire  _GEN_4306 = 3'h1 == branchTracker ? _GEN_2706 : _GEN_2186; // @[decode.scala 400:29]
  wire  _GEN_4307 = 3'h1 == branchTracker ? _GEN_2707 : _GEN_2187; // @[decode.scala 400:29]
  wire  _GEN_4308 = 3'h1 == branchTracker ? _GEN_2708 : _GEN_2188; // @[decode.scala 400:29]
  wire  _GEN_4309 = 3'h1 == branchTracker ? _GEN_2709 : _GEN_2189; // @[decode.scala 400:29]
  wire  _GEN_4310 = 3'h1 == branchTracker ? _GEN_2710 : _GEN_2190; // @[decode.scala 400:29]
  wire  _GEN_4311 = 3'h1 == branchTracker ? _GEN_2711 : _GEN_2191; // @[decode.scala 400:29]
  wire  _GEN_4312 = 3'h1 == branchTracker ? _GEN_2712 : _GEN_2192; // @[decode.scala 400:29]
  wire  _GEN_4313 = 3'h1 == branchTracker ? _GEN_2713 : _GEN_2193; // @[decode.scala 400:29]
  wire  _GEN_4314 = 3'h1 == branchTracker ? _GEN_2714 : _GEN_2194; // @[decode.scala 400:29]
  wire  _GEN_4315 = 3'h1 == branchTracker ? _GEN_2715 : _GEN_2195; // @[decode.scala 400:29]
  wire  _GEN_4316 = 3'h1 == branchTracker ? _GEN_2716 : _GEN_2196; // @[decode.scala 400:29]
  wire  _GEN_4317 = 3'h1 == branchTracker ? _GEN_2717 : _GEN_2197; // @[decode.scala 400:29]
  wire  _GEN_4318 = 3'h1 == branchTracker ? _GEN_2718 : _GEN_2198; // @[decode.scala 400:29]
  wire  _GEN_4319 = 3'h1 == branchTracker ? _GEN_2719 : _GEN_2199; // @[decode.scala 400:29]
  wire  _GEN_4320 = 3'h1 == branchTracker ? _GEN_2720 : _GEN_2200; // @[decode.scala 400:29]
  wire  _GEN_4321 = 3'h1 == branchTracker ? _GEN_2721 : _GEN_2201; // @[decode.scala 400:29]
  wire  _GEN_4322 = 3'h1 == branchTracker ? _GEN_2722 : _GEN_2202; // @[decode.scala 400:29]
  wire  _GEN_4323 = 3'h1 == branchTracker ? _GEN_2723 : _GEN_2203; // @[decode.scala 400:29]
  wire  _GEN_4324 = 3'h1 == branchTracker ? _GEN_2724 : _GEN_2204; // @[decode.scala 400:29]
  wire  _GEN_4325 = 3'h1 == branchTracker ? _GEN_2725 : _GEN_2205; // @[decode.scala 400:29]
  wire  _GEN_4326 = 3'h1 == branchTracker ? _GEN_2726 : _GEN_2206; // @[decode.scala 400:29]
  wire  _GEN_4327 = 3'h1 == branchTracker ? _GEN_2727 : _GEN_2207; // @[decode.scala 400:29]
  wire  _GEN_4328 = 3'h1 == branchTracker ? _GEN_2728 : _GEN_2208; // @[decode.scala 400:29]
  wire  _GEN_4329 = 3'h1 == branchTracker ? _GEN_2729 : _GEN_2209; // @[decode.scala 400:29]
  wire  _GEN_4330 = 3'h1 == branchTracker ? _GEN_2730 : _GEN_2210; // @[decode.scala 400:29]
  wire  _GEN_4331 = 3'h1 == branchTracker ? _GEN_2731 : _GEN_2211; // @[decode.scala 400:29]
  wire  _GEN_4332 = 3'h1 == branchTracker ? _GEN_2732 : _GEN_2212; // @[decode.scala 400:29]
  wire  _GEN_4333 = 3'h1 == branchTracker ? _GEN_2733 : _GEN_2213; // @[decode.scala 400:29]
  wire  _GEN_4334 = 3'h1 == branchTracker ? _GEN_2734 : _GEN_2214; // @[decode.scala 400:29]
  wire  _GEN_4335 = 3'h1 == branchTracker ? _GEN_2735 : _GEN_2215; // @[decode.scala 400:29]
  wire  _GEN_4336 = 3'h1 == branchTracker ? _GEN_2736 : _GEN_2216; // @[decode.scala 400:29]
  wire  _GEN_4337 = 3'h1 == branchTracker ? _GEN_2737 : _GEN_2217; // @[decode.scala 400:29]
  wire  _GEN_4338 = 3'h1 == branchTracker ? _GEN_2738 : _GEN_2218; // @[decode.scala 400:29]
  wire  _GEN_4339 = 3'h1 == branchTracker ? _GEN_2739 : _GEN_2219; // @[decode.scala 400:29]
  wire  _GEN_4340 = 3'h1 == branchTracker ? _GEN_2740 : _GEN_2220; // @[decode.scala 400:29]
  wire  _GEN_4341 = 3'h1 == branchTracker ? _GEN_2741 : _GEN_2221; // @[decode.scala 400:29]
  wire  _GEN_4342 = 3'h1 == branchTracker ? _GEN_2742 : _GEN_2222; // @[decode.scala 400:29]
  wire  _GEN_4343 = 3'h1 == branchTracker ? _GEN_2743 : _GEN_2223; // @[decode.scala 400:29]
  wire  _GEN_4344 = 3'h1 == branchTracker ? _GEN_2744 : _GEN_2224; // @[decode.scala 400:29]
  wire  _GEN_4345 = 3'h1 == branchTracker ? _GEN_2745 : _GEN_2225; // @[decode.scala 400:29]
  wire  _GEN_4346 = 3'h1 == branchTracker ? _GEN_2746 : _GEN_2226; // @[decode.scala 400:29]
  wire  _GEN_4347 = 3'h1 == branchTracker ? _GEN_2747 : _GEN_2227; // @[decode.scala 400:29]
  wire  _GEN_4348 = 3'h1 == branchTracker ? _GEN_2748 : _GEN_2228; // @[decode.scala 400:29]
  wire  _GEN_4349 = 3'h1 == branchTracker ? _GEN_2749 : _GEN_2229; // @[decode.scala 400:29]
  wire  _GEN_4350 = 3'h1 == branchTracker ? _GEN_2750 : _GEN_2230; // @[decode.scala 400:29]
  wire  _GEN_4351 = 3'h1 == branchTracker ? _GEN_2751 : _GEN_2231; // @[decode.scala 400:29]
  wire  _GEN_4352 = 3'h1 == branchTracker ? _GEN_2752 : _GEN_2232; // @[decode.scala 400:29]
  wire  _GEN_4353 = 3'h1 == branchTracker ? _GEN_2753 : _GEN_2233; // @[decode.scala 400:29]
  wire  _GEN_4354 = 3'h1 == branchTracker ? _GEN_2754 : _GEN_2234; // @[decode.scala 400:29]
  wire  _GEN_4355 = 3'h1 == branchTracker ? _GEN_2755 : _GEN_2235; // @[decode.scala 400:29]
  wire  _GEN_4356 = 3'h1 == branchTracker ? _GEN_2756 : _GEN_2236; // @[decode.scala 400:29]
  wire  _GEN_4357 = 3'h1 == branchTracker ? _GEN_2757 : _GEN_2237; // @[decode.scala 400:29]
  wire  _GEN_4358 = 3'h1 == branchTracker ? _GEN_2758 : _GEN_2238; // @[decode.scala 400:29]
  wire  _GEN_4456 = 3'h1 == branchTracker ? _GEN_2240 : _GEN_3976; // @[decode.scala 400:29]
  wire  _GEN_4457 = 3'h1 == branchTracker ? _GEN_2241 : _GEN_3977; // @[decode.scala 400:29]
  wire  _GEN_4458 = 3'h1 == branchTracker ? _GEN_2242 : _GEN_3978; // @[decode.scala 400:29]
  wire  _GEN_4459 = 3'h1 == branchTracker ? _GEN_2243 : _GEN_3979; // @[decode.scala 400:29]
  wire  _GEN_4460 = 3'h1 == branchTracker ? _GEN_2244 : _GEN_3980; // @[decode.scala 400:29]
  wire  _GEN_4461 = 3'h1 == branchTracker ? _GEN_2245 : _GEN_3981; // @[decode.scala 400:29]
  wire  _GEN_4462 = 3'h1 == branchTracker ? _GEN_2246 : _GEN_3982; // @[decode.scala 400:29]
  wire  _GEN_4463 = 3'h1 == branchTracker ? _GEN_2247 : _GEN_3983; // @[decode.scala 400:29]
  wire  _GEN_4464 = 3'h1 == branchTracker ? _GEN_2248 : _GEN_3984; // @[decode.scala 400:29]
  wire  _GEN_4465 = 3'h1 == branchTracker ? _GEN_2249 : _GEN_3985; // @[decode.scala 400:29]
  wire  _GEN_4466 = 3'h1 == branchTracker ? _GEN_2250 : _GEN_3986; // @[decode.scala 400:29]
  wire  _GEN_4467 = 3'h1 == branchTracker ? _GEN_2251 : _GEN_3987; // @[decode.scala 400:29]
  wire  _GEN_4468 = 3'h1 == branchTracker ? _GEN_2252 : _GEN_3988; // @[decode.scala 400:29]
  wire  _GEN_4469 = 3'h1 == branchTracker ? _GEN_2253 : _GEN_3989; // @[decode.scala 400:29]
  wire  _GEN_4470 = 3'h1 == branchTracker ? _GEN_2254 : _GEN_3990; // @[decode.scala 400:29]
  wire  _GEN_4471 = 3'h1 == branchTracker ? _GEN_2255 : _GEN_3991; // @[decode.scala 400:29]
  wire  _GEN_4472 = 3'h1 == branchTracker ? _GEN_2256 : _GEN_3992; // @[decode.scala 400:29]
  wire  _GEN_4473 = 3'h1 == branchTracker ? _GEN_2257 : _GEN_3993; // @[decode.scala 400:29]
  wire  _GEN_4474 = 3'h1 == branchTracker ? _GEN_2258 : _GEN_3994; // @[decode.scala 400:29]
  wire  _GEN_4475 = 3'h1 == branchTracker ? _GEN_2259 : _GEN_3995; // @[decode.scala 400:29]
  wire  _GEN_4476 = 3'h1 == branchTracker ? _GEN_2260 : _GEN_3996; // @[decode.scala 400:29]
  wire  _GEN_4477 = 3'h1 == branchTracker ? _GEN_2261 : _GEN_3997; // @[decode.scala 400:29]
  wire  _GEN_4478 = 3'h1 == branchTracker ? _GEN_2262 : _GEN_3998; // @[decode.scala 400:29]
  wire  _GEN_4479 = 3'h1 == branchTracker ? _GEN_2263 : _GEN_3999; // @[decode.scala 400:29]
  wire  _GEN_4480 = 3'h1 == branchTracker ? _GEN_2264 : _GEN_4000; // @[decode.scala 400:29]
  wire  _GEN_4481 = 3'h1 == branchTracker ? _GEN_2265 : _GEN_4001; // @[decode.scala 400:29]
  wire  _GEN_4482 = 3'h1 == branchTracker ? _GEN_2266 : _GEN_4002; // @[decode.scala 400:29]
  wire  _GEN_4483 = 3'h1 == branchTracker ? _GEN_2267 : _GEN_4003; // @[decode.scala 400:29]
  wire  _GEN_4484 = 3'h1 == branchTracker ? _GEN_2268 : _GEN_4004; // @[decode.scala 400:29]
  wire  _GEN_4485 = 3'h1 == branchTracker ? _GEN_2269 : _GEN_4005; // @[decode.scala 400:29]
  wire  _GEN_4486 = 3'h1 == branchTracker ? _GEN_2270 : _GEN_4006; // @[decode.scala 400:29]
  wire  _GEN_4487 = 3'h1 == branchTracker ? _GEN_2271 : _GEN_4007; // @[decode.scala 400:29]
  wire  _GEN_4488 = 3'h1 == branchTracker ? _GEN_2272 : _GEN_4008; // @[decode.scala 400:29]
  wire  _GEN_4489 = 3'h1 == branchTracker ? _GEN_2273 : _GEN_4009; // @[decode.scala 400:29]
  wire  _GEN_4490 = 3'h1 == branchTracker ? _GEN_2274 : _GEN_4010; // @[decode.scala 400:29]
  wire  _GEN_4491 = 3'h1 == branchTracker ? _GEN_2275 : _GEN_4011; // @[decode.scala 400:29]
  wire  _GEN_4492 = 3'h1 == branchTracker ? _GEN_2276 : _GEN_4012; // @[decode.scala 400:29]
  wire  _GEN_4493 = 3'h1 == branchTracker ? _GEN_2277 : _GEN_4013; // @[decode.scala 400:29]
  wire  _GEN_4494 = 3'h1 == branchTracker ? _GEN_2278 : _GEN_4014; // @[decode.scala 400:29]
  wire  _GEN_4495 = 3'h1 == branchTracker ? _GEN_2279 : _GEN_4015; // @[decode.scala 400:29]
  wire  _GEN_4496 = 3'h1 == branchTracker ? _GEN_2280 : _GEN_4016; // @[decode.scala 400:29]
  wire  _GEN_4497 = 3'h1 == branchTracker ? _GEN_2281 : _GEN_4017; // @[decode.scala 400:29]
  wire  _GEN_4498 = 3'h1 == branchTracker ? _GEN_2282 : _GEN_4018; // @[decode.scala 400:29]
  wire  _GEN_4499 = 3'h1 == branchTracker ? _GEN_2283 : _GEN_4019; // @[decode.scala 400:29]
  wire  _GEN_4500 = 3'h1 == branchTracker ? _GEN_2284 : _GEN_4020; // @[decode.scala 400:29]
  wire  _GEN_4501 = 3'h1 == branchTracker ? _GEN_2285 : _GEN_4021; // @[decode.scala 400:29]
  wire  _GEN_4502 = 3'h1 == branchTracker ? _GEN_2286 : _GEN_4022; // @[decode.scala 400:29]
  wire  _GEN_4503 = 3'h1 == branchTracker ? _GEN_2287 : _GEN_4023; // @[decode.scala 400:29]
  wire  _GEN_4504 = 3'h1 == branchTracker ? _GEN_2288 : _GEN_4024; // @[decode.scala 400:29]
  wire  _GEN_4505 = 3'h1 == branchTracker ? _GEN_2289 : _GEN_4025; // @[decode.scala 400:29]
  wire  _GEN_4506 = 3'h1 == branchTracker ? _GEN_2290 : _GEN_4026; // @[decode.scala 400:29]
  wire  _GEN_4507 = 3'h1 == branchTracker ? _GEN_2291 : _GEN_4027; // @[decode.scala 400:29]
  wire  _GEN_4508 = 3'h1 == branchTracker ? _GEN_2292 : _GEN_4028; // @[decode.scala 400:29]
  wire  _GEN_4509 = 3'h1 == branchTracker ? _GEN_2293 : _GEN_4029; // @[decode.scala 400:29]
  wire  _GEN_4510 = 3'h1 == branchTracker ? _GEN_2294 : _GEN_4030; // @[decode.scala 400:29]
  wire  _GEN_4511 = 3'h1 == branchTracker ? _GEN_2295 : _GEN_4031; // @[decode.scala 400:29]
  wire  _GEN_4512 = 3'h1 == branchTracker ? _GEN_2296 : _GEN_4032; // @[decode.scala 400:29]
  wire  _GEN_4513 = 3'h1 == branchTracker ? _GEN_2297 : _GEN_4033; // @[decode.scala 400:29]
  wire  _GEN_4514 = 3'h1 == branchTracker ? _GEN_2298 : _GEN_4034; // @[decode.scala 400:29]
  wire  _GEN_4515 = 3'h1 == branchTracker ? _GEN_2299 : _GEN_4035; // @[decode.scala 400:29]
  wire  _GEN_4516 = 3'h1 == branchTracker ? _GEN_2300 : _GEN_4036; // @[decode.scala 400:29]
  wire  _GEN_4517 = 3'h1 == branchTracker ? _GEN_2301 : _GEN_4037; // @[decode.scala 400:29]
  wire  _GEN_4518 = 3'h1 == branchTracker ? _GEN_2302 : _GEN_4038; // @[decode.scala 400:29]
  wire  _GEN_4616 = 3'h1 == branchTracker ? reservedFreeList4_0 : _GEN_4136; // @[decode.scala 400:29 318:30]
  wire  _GEN_4617 = 3'h1 == branchTracker ? reservedFreeList4_1 : _GEN_4137; // @[decode.scala 400:29 318:30]
  wire  _GEN_4618 = 3'h1 == branchTracker ? reservedFreeList4_2 : _GEN_4138; // @[decode.scala 400:29 318:30]
  wire  _GEN_4619 = 3'h1 == branchTracker ? reservedFreeList4_3 : _GEN_4139; // @[decode.scala 400:29 318:30]
  wire  _GEN_4620 = 3'h1 == branchTracker ? reservedFreeList4_4 : _GEN_4140; // @[decode.scala 400:29 318:30]
  wire  _GEN_4621 = 3'h1 == branchTracker ? reservedFreeList4_5 : _GEN_4141; // @[decode.scala 400:29 318:30]
  wire  _GEN_4622 = 3'h1 == branchTracker ? reservedFreeList4_6 : _GEN_4142; // @[decode.scala 400:29 318:30]
  wire  _GEN_4623 = 3'h1 == branchTracker ? reservedFreeList4_7 : _GEN_4143; // @[decode.scala 400:29 318:30]
  wire  _GEN_4624 = 3'h1 == branchTracker ? reservedFreeList4_8 : _GEN_4144; // @[decode.scala 400:29 318:30]
  wire  _GEN_4625 = 3'h1 == branchTracker ? reservedFreeList4_9 : _GEN_4145; // @[decode.scala 400:29 318:30]
  wire  _GEN_4626 = 3'h1 == branchTracker ? reservedFreeList4_10 : _GEN_4146; // @[decode.scala 400:29 318:30]
  wire  _GEN_4627 = 3'h1 == branchTracker ? reservedFreeList4_11 : _GEN_4147; // @[decode.scala 400:29 318:30]
  wire  _GEN_4628 = 3'h1 == branchTracker ? reservedFreeList4_12 : _GEN_4148; // @[decode.scala 400:29 318:30]
  wire  _GEN_4629 = 3'h1 == branchTracker ? reservedFreeList4_13 : _GEN_4149; // @[decode.scala 400:29 318:30]
  wire  _GEN_4630 = 3'h1 == branchTracker ? reservedFreeList4_14 : _GEN_4150; // @[decode.scala 400:29 318:30]
  wire  _GEN_4631 = 3'h1 == branchTracker ? reservedFreeList4_15 : _GEN_4151; // @[decode.scala 400:29 318:30]
  wire  _GEN_4632 = 3'h1 == branchTracker ? reservedFreeList4_16 : _GEN_4152; // @[decode.scala 400:29 318:30]
  wire  _GEN_4633 = 3'h1 == branchTracker ? reservedFreeList4_17 : _GEN_4153; // @[decode.scala 400:29 318:30]
  wire  _GEN_4634 = 3'h1 == branchTracker ? reservedFreeList4_18 : _GEN_4154; // @[decode.scala 400:29 318:30]
  wire  _GEN_4635 = 3'h1 == branchTracker ? reservedFreeList4_19 : _GEN_4155; // @[decode.scala 400:29 318:30]
  wire  _GEN_4636 = 3'h1 == branchTracker ? reservedFreeList4_20 : _GEN_4156; // @[decode.scala 400:29 318:30]
  wire  _GEN_4637 = 3'h1 == branchTracker ? reservedFreeList4_21 : _GEN_4157; // @[decode.scala 400:29 318:30]
  wire  _GEN_4638 = 3'h1 == branchTracker ? reservedFreeList4_22 : _GEN_4158; // @[decode.scala 400:29 318:30]
  wire  _GEN_4639 = 3'h1 == branchTracker ? reservedFreeList4_23 : _GEN_4159; // @[decode.scala 400:29 318:30]
  wire  _GEN_4640 = 3'h1 == branchTracker ? reservedFreeList4_24 : _GEN_4160; // @[decode.scala 400:29 318:30]
  wire  _GEN_4641 = 3'h1 == branchTracker ? reservedFreeList4_25 : _GEN_4161; // @[decode.scala 400:29 318:30]
  wire  _GEN_4642 = 3'h1 == branchTracker ? reservedFreeList4_26 : _GEN_4162; // @[decode.scala 400:29 318:30]
  wire  _GEN_4643 = 3'h1 == branchTracker ? reservedFreeList4_27 : _GEN_4163; // @[decode.scala 400:29 318:30]
  wire  _GEN_4644 = 3'h1 == branchTracker ? reservedFreeList4_28 : _GEN_4164; // @[decode.scala 400:29 318:30]
  wire  _GEN_4645 = 3'h1 == branchTracker ? reservedFreeList4_29 : _GEN_4165; // @[decode.scala 400:29 318:30]
  wire  _GEN_4646 = 3'h1 == branchTracker ? reservedFreeList4_30 : _GEN_4166; // @[decode.scala 400:29 318:30]
  wire  _GEN_4647 = 3'h1 == branchTracker ? reservedFreeList4_31 : _GEN_4167; // @[decode.scala 400:29 318:30]
  wire  _GEN_4648 = 3'h1 == branchTracker ? reservedFreeList4_32 : _GEN_4168; // @[decode.scala 400:29 318:30]
  wire  _GEN_4649 = 3'h1 == branchTracker ? reservedFreeList4_33 : _GEN_4169; // @[decode.scala 400:29 318:30]
  wire  _GEN_4650 = 3'h1 == branchTracker ? reservedFreeList4_34 : _GEN_4170; // @[decode.scala 400:29 318:30]
  wire  _GEN_4651 = 3'h1 == branchTracker ? reservedFreeList4_35 : _GEN_4171; // @[decode.scala 400:29 318:30]
  wire  _GEN_4652 = 3'h1 == branchTracker ? reservedFreeList4_36 : _GEN_4172; // @[decode.scala 400:29 318:30]
  wire  _GEN_4653 = 3'h1 == branchTracker ? reservedFreeList4_37 : _GEN_4173; // @[decode.scala 400:29 318:30]
  wire  _GEN_4654 = 3'h1 == branchTracker ? reservedFreeList4_38 : _GEN_4174; // @[decode.scala 400:29 318:30]
  wire  _GEN_4655 = 3'h1 == branchTracker ? reservedFreeList4_39 : _GEN_4175; // @[decode.scala 400:29 318:30]
  wire  _GEN_4656 = 3'h1 == branchTracker ? reservedFreeList4_40 : _GEN_4176; // @[decode.scala 400:29 318:30]
  wire  _GEN_4657 = 3'h1 == branchTracker ? reservedFreeList4_41 : _GEN_4177; // @[decode.scala 400:29 318:30]
  wire  _GEN_4658 = 3'h1 == branchTracker ? reservedFreeList4_42 : _GEN_4178; // @[decode.scala 400:29 318:30]
  wire  _GEN_4659 = 3'h1 == branchTracker ? reservedFreeList4_43 : _GEN_4179; // @[decode.scala 400:29 318:30]
  wire  _GEN_4660 = 3'h1 == branchTracker ? reservedFreeList4_44 : _GEN_4180; // @[decode.scala 400:29 318:30]
  wire  _GEN_4661 = 3'h1 == branchTracker ? reservedFreeList4_45 : _GEN_4181; // @[decode.scala 400:29 318:30]
  wire  _GEN_4662 = 3'h1 == branchTracker ? reservedFreeList4_46 : _GEN_4182; // @[decode.scala 400:29 318:30]
  wire  _GEN_4663 = 3'h1 == branchTracker ? reservedFreeList4_47 : _GEN_4183; // @[decode.scala 400:29 318:30]
  wire  _GEN_4664 = 3'h1 == branchTracker ? reservedFreeList4_48 : _GEN_4184; // @[decode.scala 400:29 318:30]
  wire  _GEN_4665 = 3'h1 == branchTracker ? reservedFreeList4_49 : _GEN_4185; // @[decode.scala 400:29 318:30]
  wire  _GEN_4666 = 3'h1 == branchTracker ? reservedFreeList4_50 : _GEN_4186; // @[decode.scala 400:29 318:30]
  wire  _GEN_4667 = 3'h1 == branchTracker ? reservedFreeList4_51 : _GEN_4187; // @[decode.scala 400:29 318:30]
  wire  _GEN_4668 = 3'h1 == branchTracker ? reservedFreeList4_52 : _GEN_4188; // @[decode.scala 400:29 318:30]
  wire  _GEN_4669 = 3'h1 == branchTracker ? reservedFreeList4_53 : _GEN_4189; // @[decode.scala 400:29 318:30]
  wire  _GEN_4670 = 3'h1 == branchTracker ? reservedFreeList4_54 : _GEN_4190; // @[decode.scala 400:29 318:30]
  wire  _GEN_4671 = 3'h1 == branchTracker ? reservedFreeList4_55 : _GEN_4191; // @[decode.scala 400:29 318:30]
  wire  _GEN_4672 = 3'h1 == branchTracker ? reservedFreeList4_56 : _GEN_4192; // @[decode.scala 400:29 318:30]
  wire  _GEN_4673 = 3'h1 == branchTracker ? reservedFreeList4_57 : _GEN_4193; // @[decode.scala 400:29 318:30]
  wire  _GEN_4674 = 3'h1 == branchTracker ? reservedFreeList4_58 : _GEN_4194; // @[decode.scala 400:29 318:30]
  wire  _GEN_4675 = 3'h1 == branchTracker ? reservedFreeList4_59 : _GEN_4195; // @[decode.scala 400:29 318:30]
  wire  _GEN_4676 = 3'h1 == branchTracker ? reservedFreeList4_60 : _GEN_4196; // @[decode.scala 400:29 318:30]
  wire  _GEN_4677 = 3'h1 == branchTracker ? reservedFreeList4_61 : _GEN_4197; // @[decode.scala 400:29 318:30]
  wire  _GEN_4678 = 3'h1 == branchTracker ? reservedFreeList4_62 : _GEN_4198; // @[decode.scala 400:29 318:30]
  wire  _GEN_4776 = 3'h0 == branchTracker ? _GEN_2696 : _GEN_2112; // @[decode.scala 400:29]
  wire  _GEN_4777 = 3'h0 == branchTracker ? _GEN_2697 : _GEN_2113; // @[decode.scala 400:29]
  wire  _GEN_4778 = 3'h0 == branchTracker ? _GEN_2698 : _GEN_2114; // @[decode.scala 400:29]
  wire  _GEN_4779 = 3'h0 == branchTracker ? _GEN_2699 : _GEN_2115; // @[decode.scala 400:29]
  wire  _GEN_4780 = 3'h0 == branchTracker ? _GEN_2700 : _GEN_2116; // @[decode.scala 400:29]
  wire  _GEN_4781 = 3'h0 == branchTracker ? _GEN_2701 : _GEN_2117; // @[decode.scala 400:29]
  wire  _GEN_4782 = 3'h0 == branchTracker ? _GEN_2702 : _GEN_2118; // @[decode.scala 400:29]
  wire  _GEN_4783 = 3'h0 == branchTracker ? _GEN_2703 : _GEN_2119; // @[decode.scala 400:29]
  wire  _GEN_4784 = 3'h0 == branchTracker ? _GEN_2704 : _GEN_2120; // @[decode.scala 400:29]
  wire  _GEN_4785 = 3'h0 == branchTracker ? _GEN_2705 : _GEN_2121; // @[decode.scala 400:29]
  wire  _GEN_4786 = 3'h0 == branchTracker ? _GEN_2706 : _GEN_2122; // @[decode.scala 400:29]
  wire  _GEN_4787 = 3'h0 == branchTracker ? _GEN_2707 : _GEN_2123; // @[decode.scala 400:29]
  wire  _GEN_4788 = 3'h0 == branchTracker ? _GEN_2708 : _GEN_2124; // @[decode.scala 400:29]
  wire  _GEN_4789 = 3'h0 == branchTracker ? _GEN_2709 : _GEN_2125; // @[decode.scala 400:29]
  wire  _GEN_4790 = 3'h0 == branchTracker ? _GEN_2710 : _GEN_2126; // @[decode.scala 400:29]
  wire  _GEN_4791 = 3'h0 == branchTracker ? _GEN_2711 : _GEN_2127; // @[decode.scala 400:29]
  wire  _GEN_4792 = 3'h0 == branchTracker ? _GEN_2712 : _GEN_2128; // @[decode.scala 400:29]
  wire  _GEN_4793 = 3'h0 == branchTracker ? _GEN_2713 : _GEN_2129; // @[decode.scala 400:29]
  wire  _GEN_4794 = 3'h0 == branchTracker ? _GEN_2714 : _GEN_2130; // @[decode.scala 400:29]
  wire  _GEN_4795 = 3'h0 == branchTracker ? _GEN_2715 : _GEN_2131; // @[decode.scala 400:29]
  wire  _GEN_4796 = 3'h0 == branchTracker ? _GEN_2716 : _GEN_2132; // @[decode.scala 400:29]
  wire  _GEN_4797 = 3'h0 == branchTracker ? _GEN_2717 : _GEN_2133; // @[decode.scala 400:29]
  wire  _GEN_4798 = 3'h0 == branchTracker ? _GEN_2718 : _GEN_2134; // @[decode.scala 400:29]
  wire  _GEN_4799 = 3'h0 == branchTracker ? _GEN_2719 : _GEN_2135; // @[decode.scala 400:29]
  wire  _GEN_4800 = 3'h0 == branchTracker ? _GEN_2720 : _GEN_2136; // @[decode.scala 400:29]
  wire  _GEN_4801 = 3'h0 == branchTracker ? _GEN_2721 : _GEN_2137; // @[decode.scala 400:29]
  wire  _GEN_4802 = 3'h0 == branchTracker ? _GEN_2722 : _GEN_2138; // @[decode.scala 400:29]
  wire  _GEN_4803 = 3'h0 == branchTracker ? _GEN_2723 : _GEN_2139; // @[decode.scala 400:29]
  wire  _GEN_4804 = 3'h0 == branchTracker ? _GEN_2724 : _GEN_2140; // @[decode.scala 400:29]
  wire  _GEN_4805 = 3'h0 == branchTracker ? _GEN_2725 : _GEN_2141; // @[decode.scala 400:29]
  wire  _GEN_4806 = 3'h0 == branchTracker ? _GEN_2726 : _GEN_2142; // @[decode.scala 400:29]
  wire  _GEN_4807 = 3'h0 == branchTracker ? _GEN_2727 : _GEN_2143; // @[decode.scala 400:29]
  wire  _GEN_4808 = 3'h0 == branchTracker ? _GEN_2728 : _GEN_2144; // @[decode.scala 400:29]
  wire  _GEN_4809 = 3'h0 == branchTracker ? _GEN_2729 : _GEN_2145; // @[decode.scala 400:29]
  wire  _GEN_4810 = 3'h0 == branchTracker ? _GEN_2730 : _GEN_2146; // @[decode.scala 400:29]
  wire  _GEN_4811 = 3'h0 == branchTracker ? _GEN_2731 : _GEN_2147; // @[decode.scala 400:29]
  wire  _GEN_4812 = 3'h0 == branchTracker ? _GEN_2732 : _GEN_2148; // @[decode.scala 400:29]
  wire  _GEN_4813 = 3'h0 == branchTracker ? _GEN_2733 : _GEN_2149; // @[decode.scala 400:29]
  wire  _GEN_4814 = 3'h0 == branchTracker ? _GEN_2734 : _GEN_2150; // @[decode.scala 400:29]
  wire  _GEN_4815 = 3'h0 == branchTracker ? _GEN_2735 : _GEN_2151; // @[decode.scala 400:29]
  wire  _GEN_4816 = 3'h0 == branchTracker ? _GEN_2736 : _GEN_2152; // @[decode.scala 400:29]
  wire  _GEN_4817 = 3'h0 == branchTracker ? _GEN_2737 : _GEN_2153; // @[decode.scala 400:29]
  wire  _GEN_4818 = 3'h0 == branchTracker ? _GEN_2738 : _GEN_2154; // @[decode.scala 400:29]
  wire  _GEN_4819 = 3'h0 == branchTracker ? _GEN_2739 : _GEN_2155; // @[decode.scala 400:29]
  wire  _GEN_4820 = 3'h0 == branchTracker ? _GEN_2740 : _GEN_2156; // @[decode.scala 400:29]
  wire  _GEN_4821 = 3'h0 == branchTracker ? _GEN_2741 : _GEN_2157; // @[decode.scala 400:29]
  wire  _GEN_4822 = 3'h0 == branchTracker ? _GEN_2742 : _GEN_2158; // @[decode.scala 400:29]
  wire  _GEN_4823 = 3'h0 == branchTracker ? _GEN_2743 : _GEN_2159; // @[decode.scala 400:29]
  wire  _GEN_4824 = 3'h0 == branchTracker ? _GEN_2744 : _GEN_2160; // @[decode.scala 400:29]
  wire  _GEN_4825 = 3'h0 == branchTracker ? _GEN_2745 : _GEN_2161; // @[decode.scala 400:29]
  wire  _GEN_4826 = 3'h0 == branchTracker ? _GEN_2746 : _GEN_2162; // @[decode.scala 400:29]
  wire  _GEN_4827 = 3'h0 == branchTracker ? _GEN_2747 : _GEN_2163; // @[decode.scala 400:29]
  wire  _GEN_4828 = 3'h0 == branchTracker ? _GEN_2748 : _GEN_2164; // @[decode.scala 400:29]
  wire  _GEN_4829 = 3'h0 == branchTracker ? _GEN_2749 : _GEN_2165; // @[decode.scala 400:29]
  wire  _GEN_4830 = 3'h0 == branchTracker ? _GEN_2750 : _GEN_2166; // @[decode.scala 400:29]
  wire  _GEN_4831 = 3'h0 == branchTracker ? _GEN_2751 : _GEN_2167; // @[decode.scala 400:29]
  wire  _GEN_4832 = 3'h0 == branchTracker ? _GEN_2752 : _GEN_2168; // @[decode.scala 400:29]
  wire  _GEN_4833 = 3'h0 == branchTracker ? _GEN_2753 : _GEN_2169; // @[decode.scala 400:29]
  wire  _GEN_4834 = 3'h0 == branchTracker ? _GEN_2754 : _GEN_2170; // @[decode.scala 400:29]
  wire  _GEN_4835 = 3'h0 == branchTracker ? _GEN_2755 : _GEN_2171; // @[decode.scala 400:29]
  wire  _GEN_4836 = 3'h0 == branchTracker ? _GEN_2756 : _GEN_2172; // @[decode.scala 400:29]
  wire  _GEN_4837 = 3'h0 == branchTracker ? _GEN_2757 : _GEN_2173; // @[decode.scala 400:29]
  wire  _GEN_4838 = 3'h0 == branchTracker ? _GEN_2758 : _GEN_2174; // @[decode.scala 400:29]
  wire  _GEN_4936 = 3'h0 == branchTracker ? _GEN_2176 : _GEN_4296; // @[decode.scala 400:29]
  wire  _GEN_4937 = 3'h0 == branchTracker ? _GEN_2177 : _GEN_4297; // @[decode.scala 400:29]
  wire  _GEN_4938 = 3'h0 == branchTracker ? _GEN_2178 : _GEN_4298; // @[decode.scala 400:29]
  wire  _GEN_4939 = 3'h0 == branchTracker ? _GEN_2179 : _GEN_4299; // @[decode.scala 400:29]
  wire  _GEN_4940 = 3'h0 == branchTracker ? _GEN_2180 : _GEN_4300; // @[decode.scala 400:29]
  wire  _GEN_4941 = 3'h0 == branchTracker ? _GEN_2181 : _GEN_4301; // @[decode.scala 400:29]
  wire  _GEN_4942 = 3'h0 == branchTracker ? _GEN_2182 : _GEN_4302; // @[decode.scala 400:29]
  wire  _GEN_4943 = 3'h0 == branchTracker ? _GEN_2183 : _GEN_4303; // @[decode.scala 400:29]
  wire  _GEN_4944 = 3'h0 == branchTracker ? _GEN_2184 : _GEN_4304; // @[decode.scala 400:29]
  wire  _GEN_4945 = 3'h0 == branchTracker ? _GEN_2185 : _GEN_4305; // @[decode.scala 400:29]
  wire  _GEN_4946 = 3'h0 == branchTracker ? _GEN_2186 : _GEN_4306; // @[decode.scala 400:29]
  wire  _GEN_4947 = 3'h0 == branchTracker ? _GEN_2187 : _GEN_4307; // @[decode.scala 400:29]
  wire  _GEN_4948 = 3'h0 == branchTracker ? _GEN_2188 : _GEN_4308; // @[decode.scala 400:29]
  wire  _GEN_4949 = 3'h0 == branchTracker ? _GEN_2189 : _GEN_4309; // @[decode.scala 400:29]
  wire  _GEN_4950 = 3'h0 == branchTracker ? _GEN_2190 : _GEN_4310; // @[decode.scala 400:29]
  wire  _GEN_4951 = 3'h0 == branchTracker ? _GEN_2191 : _GEN_4311; // @[decode.scala 400:29]
  wire  _GEN_4952 = 3'h0 == branchTracker ? _GEN_2192 : _GEN_4312; // @[decode.scala 400:29]
  wire  _GEN_4953 = 3'h0 == branchTracker ? _GEN_2193 : _GEN_4313; // @[decode.scala 400:29]
  wire  _GEN_4954 = 3'h0 == branchTracker ? _GEN_2194 : _GEN_4314; // @[decode.scala 400:29]
  wire  _GEN_4955 = 3'h0 == branchTracker ? _GEN_2195 : _GEN_4315; // @[decode.scala 400:29]
  wire  _GEN_4956 = 3'h0 == branchTracker ? _GEN_2196 : _GEN_4316; // @[decode.scala 400:29]
  wire  _GEN_4957 = 3'h0 == branchTracker ? _GEN_2197 : _GEN_4317; // @[decode.scala 400:29]
  wire  _GEN_4958 = 3'h0 == branchTracker ? _GEN_2198 : _GEN_4318; // @[decode.scala 400:29]
  wire  _GEN_4959 = 3'h0 == branchTracker ? _GEN_2199 : _GEN_4319; // @[decode.scala 400:29]
  wire  _GEN_4960 = 3'h0 == branchTracker ? _GEN_2200 : _GEN_4320; // @[decode.scala 400:29]
  wire  _GEN_4961 = 3'h0 == branchTracker ? _GEN_2201 : _GEN_4321; // @[decode.scala 400:29]
  wire  _GEN_4962 = 3'h0 == branchTracker ? _GEN_2202 : _GEN_4322; // @[decode.scala 400:29]
  wire  _GEN_4963 = 3'h0 == branchTracker ? _GEN_2203 : _GEN_4323; // @[decode.scala 400:29]
  wire  _GEN_4964 = 3'h0 == branchTracker ? _GEN_2204 : _GEN_4324; // @[decode.scala 400:29]
  wire  _GEN_4965 = 3'h0 == branchTracker ? _GEN_2205 : _GEN_4325; // @[decode.scala 400:29]
  wire  _GEN_4966 = 3'h0 == branchTracker ? _GEN_2206 : _GEN_4326; // @[decode.scala 400:29]
  wire  _GEN_4967 = 3'h0 == branchTracker ? _GEN_2207 : _GEN_4327; // @[decode.scala 400:29]
  wire  _GEN_4968 = 3'h0 == branchTracker ? _GEN_2208 : _GEN_4328; // @[decode.scala 400:29]
  wire  _GEN_4969 = 3'h0 == branchTracker ? _GEN_2209 : _GEN_4329; // @[decode.scala 400:29]
  wire  _GEN_4970 = 3'h0 == branchTracker ? _GEN_2210 : _GEN_4330; // @[decode.scala 400:29]
  wire  _GEN_4971 = 3'h0 == branchTracker ? _GEN_2211 : _GEN_4331; // @[decode.scala 400:29]
  wire  _GEN_4972 = 3'h0 == branchTracker ? _GEN_2212 : _GEN_4332; // @[decode.scala 400:29]
  wire  _GEN_4973 = 3'h0 == branchTracker ? _GEN_2213 : _GEN_4333; // @[decode.scala 400:29]
  wire  _GEN_4974 = 3'h0 == branchTracker ? _GEN_2214 : _GEN_4334; // @[decode.scala 400:29]
  wire  _GEN_4975 = 3'h0 == branchTracker ? _GEN_2215 : _GEN_4335; // @[decode.scala 400:29]
  wire  _GEN_4976 = 3'h0 == branchTracker ? _GEN_2216 : _GEN_4336; // @[decode.scala 400:29]
  wire  _GEN_4977 = 3'h0 == branchTracker ? _GEN_2217 : _GEN_4337; // @[decode.scala 400:29]
  wire  _GEN_4978 = 3'h0 == branchTracker ? _GEN_2218 : _GEN_4338; // @[decode.scala 400:29]
  wire  _GEN_4979 = 3'h0 == branchTracker ? _GEN_2219 : _GEN_4339; // @[decode.scala 400:29]
  wire  _GEN_4980 = 3'h0 == branchTracker ? _GEN_2220 : _GEN_4340; // @[decode.scala 400:29]
  wire  _GEN_4981 = 3'h0 == branchTracker ? _GEN_2221 : _GEN_4341; // @[decode.scala 400:29]
  wire  _GEN_4982 = 3'h0 == branchTracker ? _GEN_2222 : _GEN_4342; // @[decode.scala 400:29]
  wire  _GEN_4983 = 3'h0 == branchTracker ? _GEN_2223 : _GEN_4343; // @[decode.scala 400:29]
  wire  _GEN_4984 = 3'h0 == branchTracker ? _GEN_2224 : _GEN_4344; // @[decode.scala 400:29]
  wire  _GEN_4985 = 3'h0 == branchTracker ? _GEN_2225 : _GEN_4345; // @[decode.scala 400:29]
  wire  _GEN_4986 = 3'h0 == branchTracker ? _GEN_2226 : _GEN_4346; // @[decode.scala 400:29]
  wire  _GEN_4987 = 3'h0 == branchTracker ? _GEN_2227 : _GEN_4347; // @[decode.scala 400:29]
  wire  _GEN_4988 = 3'h0 == branchTracker ? _GEN_2228 : _GEN_4348; // @[decode.scala 400:29]
  wire  _GEN_4989 = 3'h0 == branchTracker ? _GEN_2229 : _GEN_4349; // @[decode.scala 400:29]
  wire  _GEN_4990 = 3'h0 == branchTracker ? _GEN_2230 : _GEN_4350; // @[decode.scala 400:29]
  wire  _GEN_4991 = 3'h0 == branchTracker ? _GEN_2231 : _GEN_4351; // @[decode.scala 400:29]
  wire  _GEN_4992 = 3'h0 == branchTracker ? _GEN_2232 : _GEN_4352; // @[decode.scala 400:29]
  wire  _GEN_4993 = 3'h0 == branchTracker ? _GEN_2233 : _GEN_4353; // @[decode.scala 400:29]
  wire  _GEN_4994 = 3'h0 == branchTracker ? _GEN_2234 : _GEN_4354; // @[decode.scala 400:29]
  wire  _GEN_4995 = 3'h0 == branchTracker ? _GEN_2235 : _GEN_4355; // @[decode.scala 400:29]
  wire  _GEN_4996 = 3'h0 == branchTracker ? _GEN_2236 : _GEN_4356; // @[decode.scala 400:29]
  wire  _GEN_4997 = 3'h0 == branchTracker ? _GEN_2237 : _GEN_4357; // @[decode.scala 400:29]
  wire  _GEN_4998 = 3'h0 == branchTracker ? _GEN_2238 : _GEN_4358; // @[decode.scala 400:29]
  wire  _GEN_5096 = 3'h0 == branchTracker ? _GEN_2240 : _GEN_4456; // @[decode.scala 400:29]
  wire  _GEN_5097 = 3'h0 == branchTracker ? _GEN_2241 : _GEN_4457; // @[decode.scala 400:29]
  wire  _GEN_5098 = 3'h0 == branchTracker ? _GEN_2242 : _GEN_4458; // @[decode.scala 400:29]
  wire  _GEN_5099 = 3'h0 == branchTracker ? _GEN_2243 : _GEN_4459; // @[decode.scala 400:29]
  wire  _GEN_5100 = 3'h0 == branchTracker ? _GEN_2244 : _GEN_4460; // @[decode.scala 400:29]
  wire  _GEN_5101 = 3'h0 == branchTracker ? _GEN_2245 : _GEN_4461; // @[decode.scala 400:29]
  wire  _GEN_5102 = 3'h0 == branchTracker ? _GEN_2246 : _GEN_4462; // @[decode.scala 400:29]
  wire  _GEN_5103 = 3'h0 == branchTracker ? _GEN_2247 : _GEN_4463; // @[decode.scala 400:29]
  wire  _GEN_5104 = 3'h0 == branchTracker ? _GEN_2248 : _GEN_4464; // @[decode.scala 400:29]
  wire  _GEN_5105 = 3'h0 == branchTracker ? _GEN_2249 : _GEN_4465; // @[decode.scala 400:29]
  wire  _GEN_5106 = 3'h0 == branchTracker ? _GEN_2250 : _GEN_4466; // @[decode.scala 400:29]
  wire  _GEN_5107 = 3'h0 == branchTracker ? _GEN_2251 : _GEN_4467; // @[decode.scala 400:29]
  wire  _GEN_5108 = 3'h0 == branchTracker ? _GEN_2252 : _GEN_4468; // @[decode.scala 400:29]
  wire  _GEN_5109 = 3'h0 == branchTracker ? _GEN_2253 : _GEN_4469; // @[decode.scala 400:29]
  wire  _GEN_5110 = 3'h0 == branchTracker ? _GEN_2254 : _GEN_4470; // @[decode.scala 400:29]
  wire  _GEN_5111 = 3'h0 == branchTracker ? _GEN_2255 : _GEN_4471; // @[decode.scala 400:29]
  wire  _GEN_5112 = 3'h0 == branchTracker ? _GEN_2256 : _GEN_4472; // @[decode.scala 400:29]
  wire  _GEN_5113 = 3'h0 == branchTracker ? _GEN_2257 : _GEN_4473; // @[decode.scala 400:29]
  wire  _GEN_5114 = 3'h0 == branchTracker ? _GEN_2258 : _GEN_4474; // @[decode.scala 400:29]
  wire  _GEN_5115 = 3'h0 == branchTracker ? _GEN_2259 : _GEN_4475; // @[decode.scala 400:29]
  wire  _GEN_5116 = 3'h0 == branchTracker ? _GEN_2260 : _GEN_4476; // @[decode.scala 400:29]
  wire  _GEN_5117 = 3'h0 == branchTracker ? _GEN_2261 : _GEN_4477; // @[decode.scala 400:29]
  wire  _GEN_5118 = 3'h0 == branchTracker ? _GEN_2262 : _GEN_4478; // @[decode.scala 400:29]
  wire  _GEN_5119 = 3'h0 == branchTracker ? _GEN_2263 : _GEN_4479; // @[decode.scala 400:29]
  wire  _GEN_5120 = 3'h0 == branchTracker ? _GEN_2264 : _GEN_4480; // @[decode.scala 400:29]
  wire  _GEN_5121 = 3'h0 == branchTracker ? _GEN_2265 : _GEN_4481; // @[decode.scala 400:29]
  wire  _GEN_5122 = 3'h0 == branchTracker ? _GEN_2266 : _GEN_4482; // @[decode.scala 400:29]
  wire  _GEN_5123 = 3'h0 == branchTracker ? _GEN_2267 : _GEN_4483; // @[decode.scala 400:29]
  wire  _GEN_5124 = 3'h0 == branchTracker ? _GEN_2268 : _GEN_4484; // @[decode.scala 400:29]
  wire  _GEN_5125 = 3'h0 == branchTracker ? _GEN_2269 : _GEN_4485; // @[decode.scala 400:29]
  wire  _GEN_5126 = 3'h0 == branchTracker ? _GEN_2270 : _GEN_4486; // @[decode.scala 400:29]
  wire  _GEN_5127 = 3'h0 == branchTracker ? _GEN_2271 : _GEN_4487; // @[decode.scala 400:29]
  wire  _GEN_5128 = 3'h0 == branchTracker ? _GEN_2272 : _GEN_4488; // @[decode.scala 400:29]
  wire  _GEN_5129 = 3'h0 == branchTracker ? _GEN_2273 : _GEN_4489; // @[decode.scala 400:29]
  wire  _GEN_5130 = 3'h0 == branchTracker ? _GEN_2274 : _GEN_4490; // @[decode.scala 400:29]
  wire  _GEN_5131 = 3'h0 == branchTracker ? _GEN_2275 : _GEN_4491; // @[decode.scala 400:29]
  wire  _GEN_5132 = 3'h0 == branchTracker ? _GEN_2276 : _GEN_4492; // @[decode.scala 400:29]
  wire  _GEN_5133 = 3'h0 == branchTracker ? _GEN_2277 : _GEN_4493; // @[decode.scala 400:29]
  wire  _GEN_5134 = 3'h0 == branchTracker ? _GEN_2278 : _GEN_4494; // @[decode.scala 400:29]
  wire  _GEN_5135 = 3'h0 == branchTracker ? _GEN_2279 : _GEN_4495; // @[decode.scala 400:29]
  wire  _GEN_5136 = 3'h0 == branchTracker ? _GEN_2280 : _GEN_4496; // @[decode.scala 400:29]
  wire  _GEN_5137 = 3'h0 == branchTracker ? _GEN_2281 : _GEN_4497; // @[decode.scala 400:29]
  wire  _GEN_5138 = 3'h0 == branchTracker ? _GEN_2282 : _GEN_4498; // @[decode.scala 400:29]
  wire  _GEN_5139 = 3'h0 == branchTracker ? _GEN_2283 : _GEN_4499; // @[decode.scala 400:29]
  wire  _GEN_5140 = 3'h0 == branchTracker ? _GEN_2284 : _GEN_4500; // @[decode.scala 400:29]
  wire  _GEN_5141 = 3'h0 == branchTracker ? _GEN_2285 : _GEN_4501; // @[decode.scala 400:29]
  wire  _GEN_5142 = 3'h0 == branchTracker ? _GEN_2286 : _GEN_4502; // @[decode.scala 400:29]
  wire  _GEN_5143 = 3'h0 == branchTracker ? _GEN_2287 : _GEN_4503; // @[decode.scala 400:29]
  wire  _GEN_5144 = 3'h0 == branchTracker ? _GEN_2288 : _GEN_4504; // @[decode.scala 400:29]
  wire  _GEN_5145 = 3'h0 == branchTracker ? _GEN_2289 : _GEN_4505; // @[decode.scala 400:29]
  wire  _GEN_5146 = 3'h0 == branchTracker ? _GEN_2290 : _GEN_4506; // @[decode.scala 400:29]
  wire  _GEN_5147 = 3'h0 == branchTracker ? _GEN_2291 : _GEN_4507; // @[decode.scala 400:29]
  wire  _GEN_5148 = 3'h0 == branchTracker ? _GEN_2292 : _GEN_4508; // @[decode.scala 400:29]
  wire  _GEN_5149 = 3'h0 == branchTracker ? _GEN_2293 : _GEN_4509; // @[decode.scala 400:29]
  wire  _GEN_5150 = 3'h0 == branchTracker ? _GEN_2294 : _GEN_4510; // @[decode.scala 400:29]
  wire  _GEN_5151 = 3'h0 == branchTracker ? _GEN_2295 : _GEN_4511; // @[decode.scala 400:29]
  wire  _GEN_5152 = 3'h0 == branchTracker ? _GEN_2296 : _GEN_4512; // @[decode.scala 400:29]
  wire  _GEN_5153 = 3'h0 == branchTracker ? _GEN_2297 : _GEN_4513; // @[decode.scala 400:29]
  wire  _GEN_5154 = 3'h0 == branchTracker ? _GEN_2298 : _GEN_4514; // @[decode.scala 400:29]
  wire  _GEN_5155 = 3'h0 == branchTracker ? _GEN_2299 : _GEN_4515; // @[decode.scala 400:29]
  wire  _GEN_5156 = 3'h0 == branchTracker ? _GEN_2300 : _GEN_4516; // @[decode.scala 400:29]
  wire  _GEN_5157 = 3'h0 == branchTracker ? _GEN_2301 : _GEN_4517; // @[decode.scala 400:29]
  wire  _GEN_5158 = 3'h0 == branchTracker ? _GEN_2302 : _GEN_4518; // @[decode.scala 400:29]
  wire  _GEN_5256 = 3'h0 == branchTracker ? reservedFreeList4_0 : _GEN_4616; // @[decode.scala 400:29 318:30]
  wire  _GEN_5257 = 3'h0 == branchTracker ? reservedFreeList4_1 : _GEN_4617; // @[decode.scala 400:29 318:30]
  wire  _GEN_5258 = 3'h0 == branchTracker ? reservedFreeList4_2 : _GEN_4618; // @[decode.scala 400:29 318:30]
  wire  _GEN_5259 = 3'h0 == branchTracker ? reservedFreeList4_3 : _GEN_4619; // @[decode.scala 400:29 318:30]
  wire  _GEN_5260 = 3'h0 == branchTracker ? reservedFreeList4_4 : _GEN_4620; // @[decode.scala 400:29 318:30]
  wire  _GEN_5261 = 3'h0 == branchTracker ? reservedFreeList4_5 : _GEN_4621; // @[decode.scala 400:29 318:30]
  wire  _GEN_5262 = 3'h0 == branchTracker ? reservedFreeList4_6 : _GEN_4622; // @[decode.scala 400:29 318:30]
  wire  _GEN_5263 = 3'h0 == branchTracker ? reservedFreeList4_7 : _GEN_4623; // @[decode.scala 400:29 318:30]
  wire  _GEN_5264 = 3'h0 == branchTracker ? reservedFreeList4_8 : _GEN_4624; // @[decode.scala 400:29 318:30]
  wire  _GEN_5265 = 3'h0 == branchTracker ? reservedFreeList4_9 : _GEN_4625; // @[decode.scala 400:29 318:30]
  wire  _GEN_5266 = 3'h0 == branchTracker ? reservedFreeList4_10 : _GEN_4626; // @[decode.scala 400:29 318:30]
  wire  _GEN_5267 = 3'h0 == branchTracker ? reservedFreeList4_11 : _GEN_4627; // @[decode.scala 400:29 318:30]
  wire  _GEN_5268 = 3'h0 == branchTracker ? reservedFreeList4_12 : _GEN_4628; // @[decode.scala 400:29 318:30]
  wire  _GEN_5269 = 3'h0 == branchTracker ? reservedFreeList4_13 : _GEN_4629; // @[decode.scala 400:29 318:30]
  wire  _GEN_5270 = 3'h0 == branchTracker ? reservedFreeList4_14 : _GEN_4630; // @[decode.scala 400:29 318:30]
  wire  _GEN_5271 = 3'h0 == branchTracker ? reservedFreeList4_15 : _GEN_4631; // @[decode.scala 400:29 318:30]
  wire  _GEN_5272 = 3'h0 == branchTracker ? reservedFreeList4_16 : _GEN_4632; // @[decode.scala 400:29 318:30]
  wire  _GEN_5273 = 3'h0 == branchTracker ? reservedFreeList4_17 : _GEN_4633; // @[decode.scala 400:29 318:30]
  wire  _GEN_5274 = 3'h0 == branchTracker ? reservedFreeList4_18 : _GEN_4634; // @[decode.scala 400:29 318:30]
  wire  _GEN_5275 = 3'h0 == branchTracker ? reservedFreeList4_19 : _GEN_4635; // @[decode.scala 400:29 318:30]
  wire  _GEN_5276 = 3'h0 == branchTracker ? reservedFreeList4_20 : _GEN_4636; // @[decode.scala 400:29 318:30]
  wire  _GEN_5277 = 3'h0 == branchTracker ? reservedFreeList4_21 : _GEN_4637; // @[decode.scala 400:29 318:30]
  wire  _GEN_5278 = 3'h0 == branchTracker ? reservedFreeList4_22 : _GEN_4638; // @[decode.scala 400:29 318:30]
  wire  _GEN_5279 = 3'h0 == branchTracker ? reservedFreeList4_23 : _GEN_4639; // @[decode.scala 400:29 318:30]
  wire  _GEN_5280 = 3'h0 == branchTracker ? reservedFreeList4_24 : _GEN_4640; // @[decode.scala 400:29 318:30]
  wire  _GEN_5281 = 3'h0 == branchTracker ? reservedFreeList4_25 : _GEN_4641; // @[decode.scala 400:29 318:30]
  wire  _GEN_5282 = 3'h0 == branchTracker ? reservedFreeList4_26 : _GEN_4642; // @[decode.scala 400:29 318:30]
  wire  _GEN_5283 = 3'h0 == branchTracker ? reservedFreeList4_27 : _GEN_4643; // @[decode.scala 400:29 318:30]
  wire  _GEN_5284 = 3'h0 == branchTracker ? reservedFreeList4_28 : _GEN_4644; // @[decode.scala 400:29 318:30]
  wire  _GEN_5285 = 3'h0 == branchTracker ? reservedFreeList4_29 : _GEN_4645; // @[decode.scala 400:29 318:30]
  wire  _GEN_5286 = 3'h0 == branchTracker ? reservedFreeList4_30 : _GEN_4646; // @[decode.scala 400:29 318:30]
  wire  _GEN_5287 = 3'h0 == branchTracker ? reservedFreeList4_31 : _GEN_4647; // @[decode.scala 400:29 318:30]
  wire  _GEN_5288 = 3'h0 == branchTracker ? reservedFreeList4_32 : _GEN_4648; // @[decode.scala 400:29 318:30]
  wire  _GEN_5289 = 3'h0 == branchTracker ? reservedFreeList4_33 : _GEN_4649; // @[decode.scala 400:29 318:30]
  wire  _GEN_5290 = 3'h0 == branchTracker ? reservedFreeList4_34 : _GEN_4650; // @[decode.scala 400:29 318:30]
  wire  _GEN_5291 = 3'h0 == branchTracker ? reservedFreeList4_35 : _GEN_4651; // @[decode.scala 400:29 318:30]
  wire  _GEN_5292 = 3'h0 == branchTracker ? reservedFreeList4_36 : _GEN_4652; // @[decode.scala 400:29 318:30]
  wire  _GEN_5293 = 3'h0 == branchTracker ? reservedFreeList4_37 : _GEN_4653; // @[decode.scala 400:29 318:30]
  wire  _GEN_5294 = 3'h0 == branchTracker ? reservedFreeList4_38 : _GEN_4654; // @[decode.scala 400:29 318:30]
  wire  _GEN_5295 = 3'h0 == branchTracker ? reservedFreeList4_39 : _GEN_4655; // @[decode.scala 400:29 318:30]
  wire  _GEN_5296 = 3'h0 == branchTracker ? reservedFreeList4_40 : _GEN_4656; // @[decode.scala 400:29 318:30]
  wire  _GEN_5297 = 3'h0 == branchTracker ? reservedFreeList4_41 : _GEN_4657; // @[decode.scala 400:29 318:30]
  wire  _GEN_5298 = 3'h0 == branchTracker ? reservedFreeList4_42 : _GEN_4658; // @[decode.scala 400:29 318:30]
  wire  _GEN_5299 = 3'h0 == branchTracker ? reservedFreeList4_43 : _GEN_4659; // @[decode.scala 400:29 318:30]
  wire  _GEN_5300 = 3'h0 == branchTracker ? reservedFreeList4_44 : _GEN_4660; // @[decode.scala 400:29 318:30]
  wire  _GEN_5301 = 3'h0 == branchTracker ? reservedFreeList4_45 : _GEN_4661; // @[decode.scala 400:29 318:30]
  wire  _GEN_5302 = 3'h0 == branchTracker ? reservedFreeList4_46 : _GEN_4662; // @[decode.scala 400:29 318:30]
  wire  _GEN_5303 = 3'h0 == branchTracker ? reservedFreeList4_47 : _GEN_4663; // @[decode.scala 400:29 318:30]
  wire  _GEN_5304 = 3'h0 == branchTracker ? reservedFreeList4_48 : _GEN_4664; // @[decode.scala 400:29 318:30]
  wire  _GEN_5305 = 3'h0 == branchTracker ? reservedFreeList4_49 : _GEN_4665; // @[decode.scala 400:29 318:30]
  wire  _GEN_5306 = 3'h0 == branchTracker ? reservedFreeList4_50 : _GEN_4666; // @[decode.scala 400:29 318:30]
  wire  _GEN_5307 = 3'h0 == branchTracker ? reservedFreeList4_51 : _GEN_4667; // @[decode.scala 400:29 318:30]
  wire  _GEN_5308 = 3'h0 == branchTracker ? reservedFreeList4_52 : _GEN_4668; // @[decode.scala 400:29 318:30]
  wire  _GEN_5309 = 3'h0 == branchTracker ? reservedFreeList4_53 : _GEN_4669; // @[decode.scala 400:29 318:30]
  wire  _GEN_5310 = 3'h0 == branchTracker ? reservedFreeList4_54 : _GEN_4670; // @[decode.scala 400:29 318:30]
  wire  _GEN_5311 = 3'h0 == branchTracker ? reservedFreeList4_55 : _GEN_4671; // @[decode.scala 400:29 318:30]
  wire  _GEN_5312 = 3'h0 == branchTracker ? reservedFreeList4_56 : _GEN_4672; // @[decode.scala 400:29 318:30]
  wire  _GEN_5313 = 3'h0 == branchTracker ? reservedFreeList4_57 : _GEN_4673; // @[decode.scala 400:29 318:30]
  wire  _GEN_5314 = 3'h0 == branchTracker ? reservedFreeList4_58 : _GEN_4674; // @[decode.scala 400:29 318:30]
  wire  _GEN_5315 = 3'h0 == branchTracker ? reservedFreeList4_59 : _GEN_4675; // @[decode.scala 400:29 318:30]
  wire  _GEN_5316 = 3'h0 == branchTracker ? reservedFreeList4_60 : _GEN_4676; // @[decode.scala 400:29 318:30]
  wire  _GEN_5317 = 3'h0 == branchTracker ? reservedFreeList4_61 : _GEN_4677; // @[decode.scala 400:29 318:30]
  wire  _GEN_5318 = 3'h0 == branchTracker ? reservedFreeList4_62 : _GEN_4678; // @[decode.scala 400:29 318:30]
  wire [2:0] _branchTracker_T_3 = branchTracker + 3'h1; // @[decode.scala 442:38]
  wire  _GEN_5423 = _T_432 | _T_434 | _T_431 ? _GEN_4776 : _GEN_2112; // @[decode.scala 389:73]
  wire  _GEN_5424 = _T_432 | _T_434 | _T_431 ? _GEN_4777 : _GEN_2113; // @[decode.scala 389:73]
  wire  _GEN_5425 = _T_432 | _T_434 | _T_431 ? _GEN_4778 : _GEN_2114; // @[decode.scala 389:73]
  wire  _GEN_5426 = _T_432 | _T_434 | _T_431 ? _GEN_4779 : _GEN_2115; // @[decode.scala 389:73]
  wire  _GEN_5427 = _T_432 | _T_434 | _T_431 ? _GEN_4780 : _GEN_2116; // @[decode.scala 389:73]
  wire  _GEN_5428 = _T_432 | _T_434 | _T_431 ? _GEN_4781 : _GEN_2117; // @[decode.scala 389:73]
  wire  _GEN_5429 = _T_432 | _T_434 | _T_431 ? _GEN_4782 : _GEN_2118; // @[decode.scala 389:73]
  wire  _GEN_5430 = _T_432 | _T_434 | _T_431 ? _GEN_4783 : _GEN_2119; // @[decode.scala 389:73]
  wire  _GEN_5431 = _T_432 | _T_434 | _T_431 ? _GEN_4784 : _GEN_2120; // @[decode.scala 389:73]
  wire  _GEN_5432 = _T_432 | _T_434 | _T_431 ? _GEN_4785 : _GEN_2121; // @[decode.scala 389:73]
  wire  _GEN_5433 = _T_432 | _T_434 | _T_431 ? _GEN_4786 : _GEN_2122; // @[decode.scala 389:73]
  wire  _GEN_5434 = _T_432 | _T_434 | _T_431 ? _GEN_4787 : _GEN_2123; // @[decode.scala 389:73]
  wire  _GEN_5435 = _T_432 | _T_434 | _T_431 ? _GEN_4788 : _GEN_2124; // @[decode.scala 389:73]
  wire  _GEN_5436 = _T_432 | _T_434 | _T_431 ? _GEN_4789 : _GEN_2125; // @[decode.scala 389:73]
  wire  _GEN_5437 = _T_432 | _T_434 | _T_431 ? _GEN_4790 : _GEN_2126; // @[decode.scala 389:73]
  wire  _GEN_5438 = _T_432 | _T_434 | _T_431 ? _GEN_4791 : _GEN_2127; // @[decode.scala 389:73]
  wire  _GEN_5439 = _T_432 | _T_434 | _T_431 ? _GEN_4792 : _GEN_2128; // @[decode.scala 389:73]
  wire  _GEN_5440 = _T_432 | _T_434 | _T_431 ? _GEN_4793 : _GEN_2129; // @[decode.scala 389:73]
  wire  _GEN_5441 = _T_432 | _T_434 | _T_431 ? _GEN_4794 : _GEN_2130; // @[decode.scala 389:73]
  wire  _GEN_5442 = _T_432 | _T_434 | _T_431 ? _GEN_4795 : _GEN_2131; // @[decode.scala 389:73]
  wire  _GEN_5443 = _T_432 | _T_434 | _T_431 ? _GEN_4796 : _GEN_2132; // @[decode.scala 389:73]
  wire  _GEN_5444 = _T_432 | _T_434 | _T_431 ? _GEN_4797 : _GEN_2133; // @[decode.scala 389:73]
  wire  _GEN_5445 = _T_432 | _T_434 | _T_431 ? _GEN_4798 : _GEN_2134; // @[decode.scala 389:73]
  wire  _GEN_5446 = _T_432 | _T_434 | _T_431 ? _GEN_4799 : _GEN_2135; // @[decode.scala 389:73]
  wire  _GEN_5447 = _T_432 | _T_434 | _T_431 ? _GEN_4800 : _GEN_2136; // @[decode.scala 389:73]
  wire  _GEN_5448 = _T_432 | _T_434 | _T_431 ? _GEN_4801 : _GEN_2137; // @[decode.scala 389:73]
  wire  _GEN_5449 = _T_432 | _T_434 | _T_431 ? _GEN_4802 : _GEN_2138; // @[decode.scala 389:73]
  wire  _GEN_5450 = _T_432 | _T_434 | _T_431 ? _GEN_4803 : _GEN_2139; // @[decode.scala 389:73]
  wire  _GEN_5451 = _T_432 | _T_434 | _T_431 ? _GEN_4804 : _GEN_2140; // @[decode.scala 389:73]
  wire  _GEN_5452 = _T_432 | _T_434 | _T_431 ? _GEN_4805 : _GEN_2141; // @[decode.scala 389:73]
  wire  _GEN_5453 = _T_432 | _T_434 | _T_431 ? _GEN_4806 : _GEN_2142; // @[decode.scala 389:73]
  wire  _GEN_5454 = _T_432 | _T_434 | _T_431 ? _GEN_4807 : _GEN_2143; // @[decode.scala 389:73]
  wire  _GEN_5455 = _T_432 | _T_434 | _T_431 ? _GEN_4808 : _GEN_2144; // @[decode.scala 389:73]
  wire  _GEN_5456 = _T_432 | _T_434 | _T_431 ? _GEN_4809 : _GEN_2145; // @[decode.scala 389:73]
  wire  _GEN_5457 = _T_432 | _T_434 | _T_431 ? _GEN_4810 : _GEN_2146; // @[decode.scala 389:73]
  wire  _GEN_5458 = _T_432 | _T_434 | _T_431 ? _GEN_4811 : _GEN_2147; // @[decode.scala 389:73]
  wire  _GEN_5459 = _T_432 | _T_434 | _T_431 ? _GEN_4812 : _GEN_2148; // @[decode.scala 389:73]
  wire  _GEN_5460 = _T_432 | _T_434 | _T_431 ? _GEN_4813 : _GEN_2149; // @[decode.scala 389:73]
  wire  _GEN_5461 = _T_432 | _T_434 | _T_431 ? _GEN_4814 : _GEN_2150; // @[decode.scala 389:73]
  wire  _GEN_5462 = _T_432 | _T_434 | _T_431 ? _GEN_4815 : _GEN_2151; // @[decode.scala 389:73]
  wire  _GEN_5463 = _T_432 | _T_434 | _T_431 ? _GEN_4816 : _GEN_2152; // @[decode.scala 389:73]
  wire  _GEN_5464 = _T_432 | _T_434 | _T_431 ? _GEN_4817 : _GEN_2153; // @[decode.scala 389:73]
  wire  _GEN_5465 = _T_432 | _T_434 | _T_431 ? _GEN_4818 : _GEN_2154; // @[decode.scala 389:73]
  wire  _GEN_5466 = _T_432 | _T_434 | _T_431 ? _GEN_4819 : _GEN_2155; // @[decode.scala 389:73]
  wire  _GEN_5467 = _T_432 | _T_434 | _T_431 ? _GEN_4820 : _GEN_2156; // @[decode.scala 389:73]
  wire  _GEN_5468 = _T_432 | _T_434 | _T_431 ? _GEN_4821 : _GEN_2157; // @[decode.scala 389:73]
  wire  _GEN_5469 = _T_432 | _T_434 | _T_431 ? _GEN_4822 : _GEN_2158; // @[decode.scala 389:73]
  wire  _GEN_5470 = _T_432 | _T_434 | _T_431 ? _GEN_4823 : _GEN_2159; // @[decode.scala 389:73]
  wire  _GEN_5471 = _T_432 | _T_434 | _T_431 ? _GEN_4824 : _GEN_2160; // @[decode.scala 389:73]
  wire  _GEN_5472 = _T_432 | _T_434 | _T_431 ? _GEN_4825 : _GEN_2161; // @[decode.scala 389:73]
  wire  _GEN_5473 = _T_432 | _T_434 | _T_431 ? _GEN_4826 : _GEN_2162; // @[decode.scala 389:73]
  wire  _GEN_5474 = _T_432 | _T_434 | _T_431 ? _GEN_4827 : _GEN_2163; // @[decode.scala 389:73]
  wire  _GEN_5475 = _T_432 | _T_434 | _T_431 ? _GEN_4828 : _GEN_2164; // @[decode.scala 389:73]
  wire  _GEN_5476 = _T_432 | _T_434 | _T_431 ? _GEN_4829 : _GEN_2165; // @[decode.scala 389:73]
  wire  _GEN_5477 = _T_432 | _T_434 | _T_431 ? _GEN_4830 : _GEN_2166; // @[decode.scala 389:73]
  wire  _GEN_5478 = _T_432 | _T_434 | _T_431 ? _GEN_4831 : _GEN_2167; // @[decode.scala 389:73]
  wire  _GEN_5479 = _T_432 | _T_434 | _T_431 ? _GEN_4832 : _GEN_2168; // @[decode.scala 389:73]
  wire  _GEN_5480 = _T_432 | _T_434 | _T_431 ? _GEN_4833 : _GEN_2169; // @[decode.scala 389:73]
  wire  _GEN_5481 = _T_432 | _T_434 | _T_431 ? _GEN_4834 : _GEN_2170; // @[decode.scala 389:73]
  wire  _GEN_5482 = _T_432 | _T_434 | _T_431 ? _GEN_4835 : _GEN_2171; // @[decode.scala 389:73]
  wire  _GEN_5483 = _T_432 | _T_434 | _T_431 ? _GEN_4836 : _GEN_2172; // @[decode.scala 389:73]
  wire  _GEN_5484 = _T_432 | _T_434 | _T_431 ? _GEN_4837 : _GEN_2173; // @[decode.scala 389:73]
  wire  _GEN_5485 = _T_432 | _T_434 | _T_431 ? _GEN_4838 : _GEN_2174; // @[decode.scala 389:73]
  wire  _GEN_5583 = _T_432 | _T_434 | _T_431 ? _GEN_4936 : _GEN_2176; // @[decode.scala 389:73]
  wire  _GEN_5584 = _T_432 | _T_434 | _T_431 ? _GEN_4937 : _GEN_2177; // @[decode.scala 389:73]
  wire  _GEN_5585 = _T_432 | _T_434 | _T_431 ? _GEN_4938 : _GEN_2178; // @[decode.scala 389:73]
  wire  _GEN_5586 = _T_432 | _T_434 | _T_431 ? _GEN_4939 : _GEN_2179; // @[decode.scala 389:73]
  wire  _GEN_5587 = _T_432 | _T_434 | _T_431 ? _GEN_4940 : _GEN_2180; // @[decode.scala 389:73]
  wire  _GEN_5588 = _T_432 | _T_434 | _T_431 ? _GEN_4941 : _GEN_2181; // @[decode.scala 389:73]
  wire  _GEN_5589 = _T_432 | _T_434 | _T_431 ? _GEN_4942 : _GEN_2182; // @[decode.scala 389:73]
  wire  _GEN_5590 = _T_432 | _T_434 | _T_431 ? _GEN_4943 : _GEN_2183; // @[decode.scala 389:73]
  wire  _GEN_5591 = _T_432 | _T_434 | _T_431 ? _GEN_4944 : _GEN_2184; // @[decode.scala 389:73]
  wire  _GEN_5592 = _T_432 | _T_434 | _T_431 ? _GEN_4945 : _GEN_2185; // @[decode.scala 389:73]
  wire  _GEN_5593 = _T_432 | _T_434 | _T_431 ? _GEN_4946 : _GEN_2186; // @[decode.scala 389:73]
  wire  _GEN_5594 = _T_432 | _T_434 | _T_431 ? _GEN_4947 : _GEN_2187; // @[decode.scala 389:73]
  wire  _GEN_5595 = _T_432 | _T_434 | _T_431 ? _GEN_4948 : _GEN_2188; // @[decode.scala 389:73]
  wire  _GEN_5596 = _T_432 | _T_434 | _T_431 ? _GEN_4949 : _GEN_2189; // @[decode.scala 389:73]
  wire  _GEN_5597 = _T_432 | _T_434 | _T_431 ? _GEN_4950 : _GEN_2190; // @[decode.scala 389:73]
  wire  _GEN_5598 = _T_432 | _T_434 | _T_431 ? _GEN_4951 : _GEN_2191; // @[decode.scala 389:73]
  wire  _GEN_5599 = _T_432 | _T_434 | _T_431 ? _GEN_4952 : _GEN_2192; // @[decode.scala 389:73]
  wire  _GEN_5600 = _T_432 | _T_434 | _T_431 ? _GEN_4953 : _GEN_2193; // @[decode.scala 389:73]
  wire  _GEN_5601 = _T_432 | _T_434 | _T_431 ? _GEN_4954 : _GEN_2194; // @[decode.scala 389:73]
  wire  _GEN_5602 = _T_432 | _T_434 | _T_431 ? _GEN_4955 : _GEN_2195; // @[decode.scala 389:73]
  wire  _GEN_5603 = _T_432 | _T_434 | _T_431 ? _GEN_4956 : _GEN_2196; // @[decode.scala 389:73]
  wire  _GEN_5604 = _T_432 | _T_434 | _T_431 ? _GEN_4957 : _GEN_2197; // @[decode.scala 389:73]
  wire  _GEN_5605 = _T_432 | _T_434 | _T_431 ? _GEN_4958 : _GEN_2198; // @[decode.scala 389:73]
  wire  _GEN_5606 = _T_432 | _T_434 | _T_431 ? _GEN_4959 : _GEN_2199; // @[decode.scala 389:73]
  wire  _GEN_5607 = _T_432 | _T_434 | _T_431 ? _GEN_4960 : _GEN_2200; // @[decode.scala 389:73]
  wire  _GEN_5608 = _T_432 | _T_434 | _T_431 ? _GEN_4961 : _GEN_2201; // @[decode.scala 389:73]
  wire  _GEN_5609 = _T_432 | _T_434 | _T_431 ? _GEN_4962 : _GEN_2202; // @[decode.scala 389:73]
  wire  _GEN_5610 = _T_432 | _T_434 | _T_431 ? _GEN_4963 : _GEN_2203; // @[decode.scala 389:73]
  wire  _GEN_5611 = _T_432 | _T_434 | _T_431 ? _GEN_4964 : _GEN_2204; // @[decode.scala 389:73]
  wire  _GEN_5612 = _T_432 | _T_434 | _T_431 ? _GEN_4965 : _GEN_2205; // @[decode.scala 389:73]
  wire  _GEN_5613 = _T_432 | _T_434 | _T_431 ? _GEN_4966 : _GEN_2206; // @[decode.scala 389:73]
  wire  _GEN_5614 = _T_432 | _T_434 | _T_431 ? _GEN_4967 : _GEN_2207; // @[decode.scala 389:73]
  wire  _GEN_5615 = _T_432 | _T_434 | _T_431 ? _GEN_4968 : _GEN_2208; // @[decode.scala 389:73]
  wire  _GEN_5616 = _T_432 | _T_434 | _T_431 ? _GEN_4969 : _GEN_2209; // @[decode.scala 389:73]
  wire  _GEN_5617 = _T_432 | _T_434 | _T_431 ? _GEN_4970 : _GEN_2210; // @[decode.scala 389:73]
  wire  _GEN_5618 = _T_432 | _T_434 | _T_431 ? _GEN_4971 : _GEN_2211; // @[decode.scala 389:73]
  wire  _GEN_5619 = _T_432 | _T_434 | _T_431 ? _GEN_4972 : _GEN_2212; // @[decode.scala 389:73]
  wire  _GEN_5620 = _T_432 | _T_434 | _T_431 ? _GEN_4973 : _GEN_2213; // @[decode.scala 389:73]
  wire  _GEN_5621 = _T_432 | _T_434 | _T_431 ? _GEN_4974 : _GEN_2214; // @[decode.scala 389:73]
  wire  _GEN_5622 = _T_432 | _T_434 | _T_431 ? _GEN_4975 : _GEN_2215; // @[decode.scala 389:73]
  wire  _GEN_5623 = _T_432 | _T_434 | _T_431 ? _GEN_4976 : _GEN_2216; // @[decode.scala 389:73]
  wire  _GEN_5624 = _T_432 | _T_434 | _T_431 ? _GEN_4977 : _GEN_2217; // @[decode.scala 389:73]
  wire  _GEN_5625 = _T_432 | _T_434 | _T_431 ? _GEN_4978 : _GEN_2218; // @[decode.scala 389:73]
  wire  _GEN_5626 = _T_432 | _T_434 | _T_431 ? _GEN_4979 : _GEN_2219; // @[decode.scala 389:73]
  wire  _GEN_5627 = _T_432 | _T_434 | _T_431 ? _GEN_4980 : _GEN_2220; // @[decode.scala 389:73]
  wire  _GEN_5628 = _T_432 | _T_434 | _T_431 ? _GEN_4981 : _GEN_2221; // @[decode.scala 389:73]
  wire  _GEN_5629 = _T_432 | _T_434 | _T_431 ? _GEN_4982 : _GEN_2222; // @[decode.scala 389:73]
  wire  _GEN_5630 = _T_432 | _T_434 | _T_431 ? _GEN_4983 : _GEN_2223; // @[decode.scala 389:73]
  wire  _GEN_5631 = _T_432 | _T_434 | _T_431 ? _GEN_4984 : _GEN_2224; // @[decode.scala 389:73]
  wire  _GEN_5632 = _T_432 | _T_434 | _T_431 ? _GEN_4985 : _GEN_2225; // @[decode.scala 389:73]
  wire  _GEN_5633 = _T_432 | _T_434 | _T_431 ? _GEN_4986 : _GEN_2226; // @[decode.scala 389:73]
  wire  _GEN_5634 = _T_432 | _T_434 | _T_431 ? _GEN_4987 : _GEN_2227; // @[decode.scala 389:73]
  wire  _GEN_5635 = _T_432 | _T_434 | _T_431 ? _GEN_4988 : _GEN_2228; // @[decode.scala 389:73]
  wire  _GEN_5636 = _T_432 | _T_434 | _T_431 ? _GEN_4989 : _GEN_2229; // @[decode.scala 389:73]
  wire  _GEN_5637 = _T_432 | _T_434 | _T_431 ? _GEN_4990 : _GEN_2230; // @[decode.scala 389:73]
  wire  _GEN_5638 = _T_432 | _T_434 | _T_431 ? _GEN_4991 : _GEN_2231; // @[decode.scala 389:73]
  wire  _GEN_5639 = _T_432 | _T_434 | _T_431 ? _GEN_4992 : _GEN_2232; // @[decode.scala 389:73]
  wire  _GEN_5640 = _T_432 | _T_434 | _T_431 ? _GEN_4993 : _GEN_2233; // @[decode.scala 389:73]
  wire  _GEN_5641 = _T_432 | _T_434 | _T_431 ? _GEN_4994 : _GEN_2234; // @[decode.scala 389:73]
  wire  _GEN_5642 = _T_432 | _T_434 | _T_431 ? _GEN_4995 : _GEN_2235; // @[decode.scala 389:73]
  wire  _GEN_5643 = _T_432 | _T_434 | _T_431 ? _GEN_4996 : _GEN_2236; // @[decode.scala 389:73]
  wire  _GEN_5644 = _T_432 | _T_434 | _T_431 ? _GEN_4997 : _GEN_2237; // @[decode.scala 389:73]
  wire  _GEN_5645 = _T_432 | _T_434 | _T_431 ? _GEN_4998 : _GEN_2238; // @[decode.scala 389:73]
  wire  _GEN_5743 = _T_432 | _T_434 | _T_431 ? _GEN_5096 : _GEN_2240; // @[decode.scala 389:73]
  wire  _GEN_5744 = _T_432 | _T_434 | _T_431 ? _GEN_5097 : _GEN_2241; // @[decode.scala 389:73]
  wire  _GEN_5745 = _T_432 | _T_434 | _T_431 ? _GEN_5098 : _GEN_2242; // @[decode.scala 389:73]
  wire  _GEN_5746 = _T_432 | _T_434 | _T_431 ? _GEN_5099 : _GEN_2243; // @[decode.scala 389:73]
  wire  _GEN_5747 = _T_432 | _T_434 | _T_431 ? _GEN_5100 : _GEN_2244; // @[decode.scala 389:73]
  wire  _GEN_5748 = _T_432 | _T_434 | _T_431 ? _GEN_5101 : _GEN_2245; // @[decode.scala 389:73]
  wire  _GEN_5749 = _T_432 | _T_434 | _T_431 ? _GEN_5102 : _GEN_2246; // @[decode.scala 389:73]
  wire  _GEN_5750 = _T_432 | _T_434 | _T_431 ? _GEN_5103 : _GEN_2247; // @[decode.scala 389:73]
  wire  _GEN_5751 = _T_432 | _T_434 | _T_431 ? _GEN_5104 : _GEN_2248; // @[decode.scala 389:73]
  wire  _GEN_5752 = _T_432 | _T_434 | _T_431 ? _GEN_5105 : _GEN_2249; // @[decode.scala 389:73]
  wire  _GEN_5753 = _T_432 | _T_434 | _T_431 ? _GEN_5106 : _GEN_2250; // @[decode.scala 389:73]
  wire  _GEN_5754 = _T_432 | _T_434 | _T_431 ? _GEN_5107 : _GEN_2251; // @[decode.scala 389:73]
  wire  _GEN_5755 = _T_432 | _T_434 | _T_431 ? _GEN_5108 : _GEN_2252; // @[decode.scala 389:73]
  wire  _GEN_5756 = _T_432 | _T_434 | _T_431 ? _GEN_5109 : _GEN_2253; // @[decode.scala 389:73]
  wire  _GEN_5757 = _T_432 | _T_434 | _T_431 ? _GEN_5110 : _GEN_2254; // @[decode.scala 389:73]
  wire  _GEN_5758 = _T_432 | _T_434 | _T_431 ? _GEN_5111 : _GEN_2255; // @[decode.scala 389:73]
  wire  _GEN_5759 = _T_432 | _T_434 | _T_431 ? _GEN_5112 : _GEN_2256; // @[decode.scala 389:73]
  wire  _GEN_5760 = _T_432 | _T_434 | _T_431 ? _GEN_5113 : _GEN_2257; // @[decode.scala 389:73]
  wire  _GEN_5761 = _T_432 | _T_434 | _T_431 ? _GEN_5114 : _GEN_2258; // @[decode.scala 389:73]
  wire  _GEN_5762 = _T_432 | _T_434 | _T_431 ? _GEN_5115 : _GEN_2259; // @[decode.scala 389:73]
  wire  _GEN_5763 = _T_432 | _T_434 | _T_431 ? _GEN_5116 : _GEN_2260; // @[decode.scala 389:73]
  wire  _GEN_5764 = _T_432 | _T_434 | _T_431 ? _GEN_5117 : _GEN_2261; // @[decode.scala 389:73]
  wire  _GEN_5765 = _T_432 | _T_434 | _T_431 ? _GEN_5118 : _GEN_2262; // @[decode.scala 389:73]
  wire  _GEN_5766 = _T_432 | _T_434 | _T_431 ? _GEN_5119 : _GEN_2263; // @[decode.scala 389:73]
  wire  _GEN_5767 = _T_432 | _T_434 | _T_431 ? _GEN_5120 : _GEN_2264; // @[decode.scala 389:73]
  wire  _GEN_5768 = _T_432 | _T_434 | _T_431 ? _GEN_5121 : _GEN_2265; // @[decode.scala 389:73]
  wire  _GEN_5769 = _T_432 | _T_434 | _T_431 ? _GEN_5122 : _GEN_2266; // @[decode.scala 389:73]
  wire  _GEN_5770 = _T_432 | _T_434 | _T_431 ? _GEN_5123 : _GEN_2267; // @[decode.scala 389:73]
  wire  _GEN_5771 = _T_432 | _T_434 | _T_431 ? _GEN_5124 : _GEN_2268; // @[decode.scala 389:73]
  wire  _GEN_5772 = _T_432 | _T_434 | _T_431 ? _GEN_5125 : _GEN_2269; // @[decode.scala 389:73]
  wire  _GEN_5773 = _T_432 | _T_434 | _T_431 ? _GEN_5126 : _GEN_2270; // @[decode.scala 389:73]
  wire  _GEN_5774 = _T_432 | _T_434 | _T_431 ? _GEN_5127 : _GEN_2271; // @[decode.scala 389:73]
  wire  _GEN_5775 = _T_432 | _T_434 | _T_431 ? _GEN_5128 : _GEN_2272; // @[decode.scala 389:73]
  wire  _GEN_5776 = _T_432 | _T_434 | _T_431 ? _GEN_5129 : _GEN_2273; // @[decode.scala 389:73]
  wire  _GEN_5777 = _T_432 | _T_434 | _T_431 ? _GEN_5130 : _GEN_2274; // @[decode.scala 389:73]
  wire  _GEN_5778 = _T_432 | _T_434 | _T_431 ? _GEN_5131 : _GEN_2275; // @[decode.scala 389:73]
  wire  _GEN_5779 = _T_432 | _T_434 | _T_431 ? _GEN_5132 : _GEN_2276; // @[decode.scala 389:73]
  wire  _GEN_5780 = _T_432 | _T_434 | _T_431 ? _GEN_5133 : _GEN_2277; // @[decode.scala 389:73]
  wire  _GEN_5781 = _T_432 | _T_434 | _T_431 ? _GEN_5134 : _GEN_2278; // @[decode.scala 389:73]
  wire  _GEN_5782 = _T_432 | _T_434 | _T_431 ? _GEN_5135 : _GEN_2279; // @[decode.scala 389:73]
  wire  _GEN_5783 = _T_432 | _T_434 | _T_431 ? _GEN_5136 : _GEN_2280; // @[decode.scala 389:73]
  wire  _GEN_5784 = _T_432 | _T_434 | _T_431 ? _GEN_5137 : _GEN_2281; // @[decode.scala 389:73]
  wire  _GEN_5785 = _T_432 | _T_434 | _T_431 ? _GEN_5138 : _GEN_2282; // @[decode.scala 389:73]
  wire  _GEN_5786 = _T_432 | _T_434 | _T_431 ? _GEN_5139 : _GEN_2283; // @[decode.scala 389:73]
  wire  _GEN_5787 = _T_432 | _T_434 | _T_431 ? _GEN_5140 : _GEN_2284; // @[decode.scala 389:73]
  wire  _GEN_5788 = _T_432 | _T_434 | _T_431 ? _GEN_5141 : _GEN_2285; // @[decode.scala 389:73]
  wire  _GEN_5789 = _T_432 | _T_434 | _T_431 ? _GEN_5142 : _GEN_2286; // @[decode.scala 389:73]
  wire  _GEN_5790 = _T_432 | _T_434 | _T_431 ? _GEN_5143 : _GEN_2287; // @[decode.scala 389:73]
  wire  _GEN_5791 = _T_432 | _T_434 | _T_431 ? _GEN_5144 : _GEN_2288; // @[decode.scala 389:73]
  wire  _GEN_5792 = _T_432 | _T_434 | _T_431 ? _GEN_5145 : _GEN_2289; // @[decode.scala 389:73]
  wire  _GEN_5793 = _T_432 | _T_434 | _T_431 ? _GEN_5146 : _GEN_2290; // @[decode.scala 389:73]
  wire  _GEN_5794 = _T_432 | _T_434 | _T_431 ? _GEN_5147 : _GEN_2291; // @[decode.scala 389:73]
  wire  _GEN_5795 = _T_432 | _T_434 | _T_431 ? _GEN_5148 : _GEN_2292; // @[decode.scala 389:73]
  wire  _GEN_5796 = _T_432 | _T_434 | _T_431 ? _GEN_5149 : _GEN_2293; // @[decode.scala 389:73]
  wire  _GEN_5797 = _T_432 | _T_434 | _T_431 ? _GEN_5150 : _GEN_2294; // @[decode.scala 389:73]
  wire  _GEN_5798 = _T_432 | _T_434 | _T_431 ? _GEN_5151 : _GEN_2295; // @[decode.scala 389:73]
  wire  _GEN_5799 = _T_432 | _T_434 | _T_431 ? _GEN_5152 : _GEN_2296; // @[decode.scala 389:73]
  wire  _GEN_5800 = _T_432 | _T_434 | _T_431 ? _GEN_5153 : _GEN_2297; // @[decode.scala 389:73]
  wire  _GEN_5801 = _T_432 | _T_434 | _T_431 ? _GEN_5154 : _GEN_2298; // @[decode.scala 389:73]
  wire  _GEN_5802 = _T_432 | _T_434 | _T_431 ? _GEN_5155 : _GEN_2299; // @[decode.scala 389:73]
  wire  _GEN_5803 = _T_432 | _T_434 | _T_431 ? _GEN_5156 : _GEN_2300; // @[decode.scala 389:73]
  wire  _GEN_5804 = _T_432 | _T_434 | _T_431 ? _GEN_5157 : _GEN_2301; // @[decode.scala 389:73]
  wire  _GEN_5805 = _T_432 | _T_434 | _T_431 ? _GEN_5158 : _GEN_2302; // @[decode.scala 389:73]
  wire  _GEN_5903 = _T_432 | _T_434 | _T_431 ? _GEN_5256 : reservedFreeList4_0; // @[decode.scala 318:30 389:73]
  wire  _GEN_5904 = _T_432 | _T_434 | _T_431 ? _GEN_5257 : reservedFreeList4_1; // @[decode.scala 318:30 389:73]
  wire  _GEN_5905 = _T_432 | _T_434 | _T_431 ? _GEN_5258 : reservedFreeList4_2; // @[decode.scala 318:30 389:73]
  wire  _GEN_5906 = _T_432 | _T_434 | _T_431 ? _GEN_5259 : reservedFreeList4_3; // @[decode.scala 318:30 389:73]
  wire  _GEN_5907 = _T_432 | _T_434 | _T_431 ? _GEN_5260 : reservedFreeList4_4; // @[decode.scala 318:30 389:73]
  wire  _GEN_5908 = _T_432 | _T_434 | _T_431 ? _GEN_5261 : reservedFreeList4_5; // @[decode.scala 318:30 389:73]
  wire  _GEN_5909 = _T_432 | _T_434 | _T_431 ? _GEN_5262 : reservedFreeList4_6; // @[decode.scala 318:30 389:73]
  wire  _GEN_5910 = _T_432 | _T_434 | _T_431 ? _GEN_5263 : reservedFreeList4_7; // @[decode.scala 318:30 389:73]
  wire  _GEN_5911 = _T_432 | _T_434 | _T_431 ? _GEN_5264 : reservedFreeList4_8; // @[decode.scala 318:30 389:73]
  wire  _GEN_5912 = _T_432 | _T_434 | _T_431 ? _GEN_5265 : reservedFreeList4_9; // @[decode.scala 318:30 389:73]
  wire  _GEN_5913 = _T_432 | _T_434 | _T_431 ? _GEN_5266 : reservedFreeList4_10; // @[decode.scala 318:30 389:73]
  wire  _GEN_5914 = _T_432 | _T_434 | _T_431 ? _GEN_5267 : reservedFreeList4_11; // @[decode.scala 318:30 389:73]
  wire  _GEN_5915 = _T_432 | _T_434 | _T_431 ? _GEN_5268 : reservedFreeList4_12; // @[decode.scala 318:30 389:73]
  wire  _GEN_5916 = _T_432 | _T_434 | _T_431 ? _GEN_5269 : reservedFreeList4_13; // @[decode.scala 318:30 389:73]
  wire  _GEN_5917 = _T_432 | _T_434 | _T_431 ? _GEN_5270 : reservedFreeList4_14; // @[decode.scala 318:30 389:73]
  wire  _GEN_5918 = _T_432 | _T_434 | _T_431 ? _GEN_5271 : reservedFreeList4_15; // @[decode.scala 318:30 389:73]
  wire  _GEN_5919 = _T_432 | _T_434 | _T_431 ? _GEN_5272 : reservedFreeList4_16; // @[decode.scala 318:30 389:73]
  wire  _GEN_5920 = _T_432 | _T_434 | _T_431 ? _GEN_5273 : reservedFreeList4_17; // @[decode.scala 318:30 389:73]
  wire  _GEN_5921 = _T_432 | _T_434 | _T_431 ? _GEN_5274 : reservedFreeList4_18; // @[decode.scala 318:30 389:73]
  wire  _GEN_5922 = _T_432 | _T_434 | _T_431 ? _GEN_5275 : reservedFreeList4_19; // @[decode.scala 318:30 389:73]
  wire  _GEN_5923 = _T_432 | _T_434 | _T_431 ? _GEN_5276 : reservedFreeList4_20; // @[decode.scala 318:30 389:73]
  wire  _GEN_5924 = _T_432 | _T_434 | _T_431 ? _GEN_5277 : reservedFreeList4_21; // @[decode.scala 318:30 389:73]
  wire  _GEN_5925 = _T_432 | _T_434 | _T_431 ? _GEN_5278 : reservedFreeList4_22; // @[decode.scala 318:30 389:73]
  wire  _GEN_5926 = _T_432 | _T_434 | _T_431 ? _GEN_5279 : reservedFreeList4_23; // @[decode.scala 318:30 389:73]
  wire  _GEN_5927 = _T_432 | _T_434 | _T_431 ? _GEN_5280 : reservedFreeList4_24; // @[decode.scala 318:30 389:73]
  wire  _GEN_5928 = _T_432 | _T_434 | _T_431 ? _GEN_5281 : reservedFreeList4_25; // @[decode.scala 318:30 389:73]
  wire  _GEN_5929 = _T_432 | _T_434 | _T_431 ? _GEN_5282 : reservedFreeList4_26; // @[decode.scala 318:30 389:73]
  wire  _GEN_5930 = _T_432 | _T_434 | _T_431 ? _GEN_5283 : reservedFreeList4_27; // @[decode.scala 318:30 389:73]
  wire  _GEN_5931 = _T_432 | _T_434 | _T_431 ? _GEN_5284 : reservedFreeList4_28; // @[decode.scala 318:30 389:73]
  wire  _GEN_5932 = _T_432 | _T_434 | _T_431 ? _GEN_5285 : reservedFreeList4_29; // @[decode.scala 318:30 389:73]
  wire  _GEN_5933 = _T_432 | _T_434 | _T_431 ? _GEN_5286 : reservedFreeList4_30; // @[decode.scala 318:30 389:73]
  wire  _GEN_5934 = _T_432 | _T_434 | _T_431 ? _GEN_5287 : reservedFreeList4_31; // @[decode.scala 318:30 389:73]
  wire  _GEN_5935 = _T_432 | _T_434 | _T_431 ? _GEN_5288 : reservedFreeList4_32; // @[decode.scala 318:30 389:73]
  wire  _GEN_5936 = _T_432 | _T_434 | _T_431 ? _GEN_5289 : reservedFreeList4_33; // @[decode.scala 318:30 389:73]
  wire  _GEN_5937 = _T_432 | _T_434 | _T_431 ? _GEN_5290 : reservedFreeList4_34; // @[decode.scala 318:30 389:73]
  wire  _GEN_5938 = _T_432 | _T_434 | _T_431 ? _GEN_5291 : reservedFreeList4_35; // @[decode.scala 318:30 389:73]
  wire  _GEN_5939 = _T_432 | _T_434 | _T_431 ? _GEN_5292 : reservedFreeList4_36; // @[decode.scala 318:30 389:73]
  wire  _GEN_5940 = _T_432 | _T_434 | _T_431 ? _GEN_5293 : reservedFreeList4_37; // @[decode.scala 318:30 389:73]
  wire  _GEN_5941 = _T_432 | _T_434 | _T_431 ? _GEN_5294 : reservedFreeList4_38; // @[decode.scala 318:30 389:73]
  wire  _GEN_5942 = _T_432 | _T_434 | _T_431 ? _GEN_5295 : reservedFreeList4_39; // @[decode.scala 318:30 389:73]
  wire  _GEN_5943 = _T_432 | _T_434 | _T_431 ? _GEN_5296 : reservedFreeList4_40; // @[decode.scala 318:30 389:73]
  wire  _GEN_5944 = _T_432 | _T_434 | _T_431 ? _GEN_5297 : reservedFreeList4_41; // @[decode.scala 318:30 389:73]
  wire  _GEN_5945 = _T_432 | _T_434 | _T_431 ? _GEN_5298 : reservedFreeList4_42; // @[decode.scala 318:30 389:73]
  wire  _GEN_5946 = _T_432 | _T_434 | _T_431 ? _GEN_5299 : reservedFreeList4_43; // @[decode.scala 318:30 389:73]
  wire  _GEN_5947 = _T_432 | _T_434 | _T_431 ? _GEN_5300 : reservedFreeList4_44; // @[decode.scala 318:30 389:73]
  wire  _GEN_5948 = _T_432 | _T_434 | _T_431 ? _GEN_5301 : reservedFreeList4_45; // @[decode.scala 318:30 389:73]
  wire  _GEN_5949 = _T_432 | _T_434 | _T_431 ? _GEN_5302 : reservedFreeList4_46; // @[decode.scala 318:30 389:73]
  wire  _GEN_5950 = _T_432 | _T_434 | _T_431 ? _GEN_5303 : reservedFreeList4_47; // @[decode.scala 318:30 389:73]
  wire  _GEN_5951 = _T_432 | _T_434 | _T_431 ? _GEN_5304 : reservedFreeList4_48; // @[decode.scala 318:30 389:73]
  wire  _GEN_5952 = _T_432 | _T_434 | _T_431 ? _GEN_5305 : reservedFreeList4_49; // @[decode.scala 318:30 389:73]
  wire  _GEN_5953 = _T_432 | _T_434 | _T_431 ? _GEN_5306 : reservedFreeList4_50; // @[decode.scala 318:30 389:73]
  wire  _GEN_5954 = _T_432 | _T_434 | _T_431 ? _GEN_5307 : reservedFreeList4_51; // @[decode.scala 318:30 389:73]
  wire  _GEN_5955 = _T_432 | _T_434 | _T_431 ? _GEN_5308 : reservedFreeList4_52; // @[decode.scala 318:30 389:73]
  wire  _GEN_5956 = _T_432 | _T_434 | _T_431 ? _GEN_5309 : reservedFreeList4_53; // @[decode.scala 318:30 389:73]
  wire  _GEN_5957 = _T_432 | _T_434 | _T_431 ? _GEN_5310 : reservedFreeList4_54; // @[decode.scala 318:30 389:73]
  wire  _GEN_5958 = _T_432 | _T_434 | _T_431 ? _GEN_5311 : reservedFreeList4_55; // @[decode.scala 318:30 389:73]
  wire  _GEN_5959 = _T_432 | _T_434 | _T_431 ? _GEN_5312 : reservedFreeList4_56; // @[decode.scala 318:30 389:73]
  wire  _GEN_5960 = _T_432 | _T_434 | _T_431 ? _GEN_5313 : reservedFreeList4_57; // @[decode.scala 318:30 389:73]
  wire  _GEN_5961 = _T_432 | _T_434 | _T_431 ? _GEN_5314 : reservedFreeList4_58; // @[decode.scala 318:30 389:73]
  wire  _GEN_5962 = _T_432 | _T_434 | _T_431 ? _GEN_5315 : reservedFreeList4_59; // @[decode.scala 318:30 389:73]
  wire  _GEN_5963 = _T_432 | _T_434 | _T_431 ? _GEN_5316 : reservedFreeList4_60; // @[decode.scala 318:30 389:73]
  wire  _GEN_5964 = _T_432 | _T_434 | _T_431 ? _GEN_5317 : reservedFreeList4_61; // @[decode.scala 318:30 389:73]
  wire  _GEN_5965 = _T_432 | _T_434 | _T_431 ? _GEN_5318 : reservedFreeList4_62; // @[decode.scala 318:30 389:73]
  wire  _GEN_6071 = _T_3 ? _GEN_5423 : _GEN_2112; // @[decode.scala 388:41]
  wire  _GEN_6072 = _T_3 ? _GEN_5424 : _GEN_2113; // @[decode.scala 388:41]
  wire  _GEN_6073 = _T_3 ? _GEN_5425 : _GEN_2114; // @[decode.scala 388:41]
  wire  _GEN_6074 = _T_3 ? _GEN_5426 : _GEN_2115; // @[decode.scala 388:41]
  wire  _GEN_6075 = _T_3 ? _GEN_5427 : _GEN_2116; // @[decode.scala 388:41]
  wire  _GEN_6076 = _T_3 ? _GEN_5428 : _GEN_2117; // @[decode.scala 388:41]
  wire  _GEN_6077 = _T_3 ? _GEN_5429 : _GEN_2118; // @[decode.scala 388:41]
  wire  _GEN_6078 = _T_3 ? _GEN_5430 : _GEN_2119; // @[decode.scala 388:41]
  wire  _GEN_6079 = _T_3 ? _GEN_5431 : _GEN_2120; // @[decode.scala 388:41]
  wire  _GEN_6080 = _T_3 ? _GEN_5432 : _GEN_2121; // @[decode.scala 388:41]
  wire  _GEN_6081 = _T_3 ? _GEN_5433 : _GEN_2122; // @[decode.scala 388:41]
  wire  _GEN_6082 = _T_3 ? _GEN_5434 : _GEN_2123; // @[decode.scala 388:41]
  wire  _GEN_6083 = _T_3 ? _GEN_5435 : _GEN_2124; // @[decode.scala 388:41]
  wire  _GEN_6084 = _T_3 ? _GEN_5436 : _GEN_2125; // @[decode.scala 388:41]
  wire  _GEN_6085 = _T_3 ? _GEN_5437 : _GEN_2126; // @[decode.scala 388:41]
  wire  _GEN_6086 = _T_3 ? _GEN_5438 : _GEN_2127; // @[decode.scala 388:41]
  wire  _GEN_6087 = _T_3 ? _GEN_5439 : _GEN_2128; // @[decode.scala 388:41]
  wire  _GEN_6088 = _T_3 ? _GEN_5440 : _GEN_2129; // @[decode.scala 388:41]
  wire  _GEN_6089 = _T_3 ? _GEN_5441 : _GEN_2130; // @[decode.scala 388:41]
  wire  _GEN_6090 = _T_3 ? _GEN_5442 : _GEN_2131; // @[decode.scala 388:41]
  wire  _GEN_6091 = _T_3 ? _GEN_5443 : _GEN_2132; // @[decode.scala 388:41]
  wire  _GEN_6092 = _T_3 ? _GEN_5444 : _GEN_2133; // @[decode.scala 388:41]
  wire  _GEN_6093 = _T_3 ? _GEN_5445 : _GEN_2134; // @[decode.scala 388:41]
  wire  _GEN_6094 = _T_3 ? _GEN_5446 : _GEN_2135; // @[decode.scala 388:41]
  wire  _GEN_6095 = _T_3 ? _GEN_5447 : _GEN_2136; // @[decode.scala 388:41]
  wire  _GEN_6096 = _T_3 ? _GEN_5448 : _GEN_2137; // @[decode.scala 388:41]
  wire  _GEN_6097 = _T_3 ? _GEN_5449 : _GEN_2138; // @[decode.scala 388:41]
  wire  _GEN_6098 = _T_3 ? _GEN_5450 : _GEN_2139; // @[decode.scala 388:41]
  wire  _GEN_6099 = _T_3 ? _GEN_5451 : _GEN_2140; // @[decode.scala 388:41]
  wire  _GEN_6100 = _T_3 ? _GEN_5452 : _GEN_2141; // @[decode.scala 388:41]
  wire  _GEN_6101 = _T_3 ? _GEN_5453 : _GEN_2142; // @[decode.scala 388:41]
  wire  _GEN_6102 = _T_3 ? _GEN_5454 : _GEN_2143; // @[decode.scala 388:41]
  wire  _GEN_6103 = _T_3 ? _GEN_5455 : _GEN_2144; // @[decode.scala 388:41]
  wire  _GEN_6104 = _T_3 ? _GEN_5456 : _GEN_2145; // @[decode.scala 388:41]
  wire  _GEN_6105 = _T_3 ? _GEN_5457 : _GEN_2146; // @[decode.scala 388:41]
  wire  _GEN_6106 = _T_3 ? _GEN_5458 : _GEN_2147; // @[decode.scala 388:41]
  wire  _GEN_6107 = _T_3 ? _GEN_5459 : _GEN_2148; // @[decode.scala 388:41]
  wire  _GEN_6108 = _T_3 ? _GEN_5460 : _GEN_2149; // @[decode.scala 388:41]
  wire  _GEN_6109 = _T_3 ? _GEN_5461 : _GEN_2150; // @[decode.scala 388:41]
  wire  _GEN_6110 = _T_3 ? _GEN_5462 : _GEN_2151; // @[decode.scala 388:41]
  wire  _GEN_6111 = _T_3 ? _GEN_5463 : _GEN_2152; // @[decode.scala 388:41]
  wire  _GEN_6112 = _T_3 ? _GEN_5464 : _GEN_2153; // @[decode.scala 388:41]
  wire  _GEN_6113 = _T_3 ? _GEN_5465 : _GEN_2154; // @[decode.scala 388:41]
  wire  _GEN_6114 = _T_3 ? _GEN_5466 : _GEN_2155; // @[decode.scala 388:41]
  wire  _GEN_6115 = _T_3 ? _GEN_5467 : _GEN_2156; // @[decode.scala 388:41]
  wire  _GEN_6116 = _T_3 ? _GEN_5468 : _GEN_2157; // @[decode.scala 388:41]
  wire  _GEN_6117 = _T_3 ? _GEN_5469 : _GEN_2158; // @[decode.scala 388:41]
  wire  _GEN_6118 = _T_3 ? _GEN_5470 : _GEN_2159; // @[decode.scala 388:41]
  wire  _GEN_6119 = _T_3 ? _GEN_5471 : _GEN_2160; // @[decode.scala 388:41]
  wire  _GEN_6120 = _T_3 ? _GEN_5472 : _GEN_2161; // @[decode.scala 388:41]
  wire  _GEN_6121 = _T_3 ? _GEN_5473 : _GEN_2162; // @[decode.scala 388:41]
  wire  _GEN_6122 = _T_3 ? _GEN_5474 : _GEN_2163; // @[decode.scala 388:41]
  wire  _GEN_6123 = _T_3 ? _GEN_5475 : _GEN_2164; // @[decode.scala 388:41]
  wire  _GEN_6124 = _T_3 ? _GEN_5476 : _GEN_2165; // @[decode.scala 388:41]
  wire  _GEN_6125 = _T_3 ? _GEN_5477 : _GEN_2166; // @[decode.scala 388:41]
  wire  _GEN_6126 = _T_3 ? _GEN_5478 : _GEN_2167; // @[decode.scala 388:41]
  wire  _GEN_6127 = _T_3 ? _GEN_5479 : _GEN_2168; // @[decode.scala 388:41]
  wire  _GEN_6128 = _T_3 ? _GEN_5480 : _GEN_2169; // @[decode.scala 388:41]
  wire  _GEN_6129 = _T_3 ? _GEN_5481 : _GEN_2170; // @[decode.scala 388:41]
  wire  _GEN_6130 = _T_3 ? _GEN_5482 : _GEN_2171; // @[decode.scala 388:41]
  wire  _GEN_6131 = _T_3 ? _GEN_5483 : _GEN_2172; // @[decode.scala 388:41]
  wire  _GEN_6132 = _T_3 ? _GEN_5484 : _GEN_2173; // @[decode.scala 388:41]
  wire  _GEN_6133 = _T_3 ? _GEN_5485 : _GEN_2174; // @[decode.scala 388:41]
  wire  _GEN_6231 = _T_3 ? _GEN_5583 : _GEN_2176; // @[decode.scala 388:41]
  wire  _GEN_6232 = _T_3 ? _GEN_5584 : _GEN_2177; // @[decode.scala 388:41]
  wire  _GEN_6233 = _T_3 ? _GEN_5585 : _GEN_2178; // @[decode.scala 388:41]
  wire  _GEN_6234 = _T_3 ? _GEN_5586 : _GEN_2179; // @[decode.scala 388:41]
  wire  _GEN_6235 = _T_3 ? _GEN_5587 : _GEN_2180; // @[decode.scala 388:41]
  wire  _GEN_6236 = _T_3 ? _GEN_5588 : _GEN_2181; // @[decode.scala 388:41]
  wire  _GEN_6237 = _T_3 ? _GEN_5589 : _GEN_2182; // @[decode.scala 388:41]
  wire  _GEN_6238 = _T_3 ? _GEN_5590 : _GEN_2183; // @[decode.scala 388:41]
  wire  _GEN_6239 = _T_3 ? _GEN_5591 : _GEN_2184; // @[decode.scala 388:41]
  wire  _GEN_6240 = _T_3 ? _GEN_5592 : _GEN_2185; // @[decode.scala 388:41]
  wire  _GEN_6241 = _T_3 ? _GEN_5593 : _GEN_2186; // @[decode.scala 388:41]
  wire  _GEN_6242 = _T_3 ? _GEN_5594 : _GEN_2187; // @[decode.scala 388:41]
  wire  _GEN_6243 = _T_3 ? _GEN_5595 : _GEN_2188; // @[decode.scala 388:41]
  wire  _GEN_6244 = _T_3 ? _GEN_5596 : _GEN_2189; // @[decode.scala 388:41]
  wire  _GEN_6245 = _T_3 ? _GEN_5597 : _GEN_2190; // @[decode.scala 388:41]
  wire  _GEN_6246 = _T_3 ? _GEN_5598 : _GEN_2191; // @[decode.scala 388:41]
  wire  _GEN_6247 = _T_3 ? _GEN_5599 : _GEN_2192; // @[decode.scala 388:41]
  wire  _GEN_6248 = _T_3 ? _GEN_5600 : _GEN_2193; // @[decode.scala 388:41]
  wire  _GEN_6249 = _T_3 ? _GEN_5601 : _GEN_2194; // @[decode.scala 388:41]
  wire  _GEN_6250 = _T_3 ? _GEN_5602 : _GEN_2195; // @[decode.scala 388:41]
  wire  _GEN_6251 = _T_3 ? _GEN_5603 : _GEN_2196; // @[decode.scala 388:41]
  wire  _GEN_6252 = _T_3 ? _GEN_5604 : _GEN_2197; // @[decode.scala 388:41]
  wire  _GEN_6253 = _T_3 ? _GEN_5605 : _GEN_2198; // @[decode.scala 388:41]
  wire  _GEN_6254 = _T_3 ? _GEN_5606 : _GEN_2199; // @[decode.scala 388:41]
  wire  _GEN_6255 = _T_3 ? _GEN_5607 : _GEN_2200; // @[decode.scala 388:41]
  wire  _GEN_6256 = _T_3 ? _GEN_5608 : _GEN_2201; // @[decode.scala 388:41]
  wire  _GEN_6257 = _T_3 ? _GEN_5609 : _GEN_2202; // @[decode.scala 388:41]
  wire  _GEN_6258 = _T_3 ? _GEN_5610 : _GEN_2203; // @[decode.scala 388:41]
  wire  _GEN_6259 = _T_3 ? _GEN_5611 : _GEN_2204; // @[decode.scala 388:41]
  wire  _GEN_6260 = _T_3 ? _GEN_5612 : _GEN_2205; // @[decode.scala 388:41]
  wire  _GEN_6261 = _T_3 ? _GEN_5613 : _GEN_2206; // @[decode.scala 388:41]
  wire  _GEN_6262 = _T_3 ? _GEN_5614 : _GEN_2207; // @[decode.scala 388:41]
  wire  _GEN_6263 = _T_3 ? _GEN_5615 : _GEN_2208; // @[decode.scala 388:41]
  wire  _GEN_6264 = _T_3 ? _GEN_5616 : _GEN_2209; // @[decode.scala 388:41]
  wire  _GEN_6265 = _T_3 ? _GEN_5617 : _GEN_2210; // @[decode.scala 388:41]
  wire  _GEN_6266 = _T_3 ? _GEN_5618 : _GEN_2211; // @[decode.scala 388:41]
  wire  _GEN_6267 = _T_3 ? _GEN_5619 : _GEN_2212; // @[decode.scala 388:41]
  wire  _GEN_6268 = _T_3 ? _GEN_5620 : _GEN_2213; // @[decode.scala 388:41]
  wire  _GEN_6269 = _T_3 ? _GEN_5621 : _GEN_2214; // @[decode.scala 388:41]
  wire  _GEN_6270 = _T_3 ? _GEN_5622 : _GEN_2215; // @[decode.scala 388:41]
  wire  _GEN_6271 = _T_3 ? _GEN_5623 : _GEN_2216; // @[decode.scala 388:41]
  wire  _GEN_6272 = _T_3 ? _GEN_5624 : _GEN_2217; // @[decode.scala 388:41]
  wire  _GEN_6273 = _T_3 ? _GEN_5625 : _GEN_2218; // @[decode.scala 388:41]
  wire  _GEN_6274 = _T_3 ? _GEN_5626 : _GEN_2219; // @[decode.scala 388:41]
  wire  _GEN_6275 = _T_3 ? _GEN_5627 : _GEN_2220; // @[decode.scala 388:41]
  wire  _GEN_6276 = _T_3 ? _GEN_5628 : _GEN_2221; // @[decode.scala 388:41]
  wire  _GEN_6277 = _T_3 ? _GEN_5629 : _GEN_2222; // @[decode.scala 388:41]
  wire  _GEN_6278 = _T_3 ? _GEN_5630 : _GEN_2223; // @[decode.scala 388:41]
  wire  _GEN_6279 = _T_3 ? _GEN_5631 : _GEN_2224; // @[decode.scala 388:41]
  wire  _GEN_6280 = _T_3 ? _GEN_5632 : _GEN_2225; // @[decode.scala 388:41]
  wire  _GEN_6281 = _T_3 ? _GEN_5633 : _GEN_2226; // @[decode.scala 388:41]
  wire  _GEN_6282 = _T_3 ? _GEN_5634 : _GEN_2227; // @[decode.scala 388:41]
  wire  _GEN_6283 = _T_3 ? _GEN_5635 : _GEN_2228; // @[decode.scala 388:41]
  wire  _GEN_6284 = _T_3 ? _GEN_5636 : _GEN_2229; // @[decode.scala 388:41]
  wire  _GEN_6285 = _T_3 ? _GEN_5637 : _GEN_2230; // @[decode.scala 388:41]
  wire  _GEN_6286 = _T_3 ? _GEN_5638 : _GEN_2231; // @[decode.scala 388:41]
  wire  _GEN_6287 = _T_3 ? _GEN_5639 : _GEN_2232; // @[decode.scala 388:41]
  wire  _GEN_6288 = _T_3 ? _GEN_5640 : _GEN_2233; // @[decode.scala 388:41]
  wire  _GEN_6289 = _T_3 ? _GEN_5641 : _GEN_2234; // @[decode.scala 388:41]
  wire  _GEN_6290 = _T_3 ? _GEN_5642 : _GEN_2235; // @[decode.scala 388:41]
  wire  _GEN_6291 = _T_3 ? _GEN_5643 : _GEN_2236; // @[decode.scala 388:41]
  wire  _GEN_6292 = _T_3 ? _GEN_5644 : _GEN_2237; // @[decode.scala 388:41]
  wire  _GEN_6293 = _T_3 ? _GEN_5645 : _GEN_2238; // @[decode.scala 388:41]
  wire  _GEN_6391 = _T_3 ? _GEN_5743 : _GEN_2240; // @[decode.scala 388:41]
  wire  _GEN_6392 = _T_3 ? _GEN_5744 : _GEN_2241; // @[decode.scala 388:41]
  wire  _GEN_6393 = _T_3 ? _GEN_5745 : _GEN_2242; // @[decode.scala 388:41]
  wire  _GEN_6394 = _T_3 ? _GEN_5746 : _GEN_2243; // @[decode.scala 388:41]
  wire  _GEN_6395 = _T_3 ? _GEN_5747 : _GEN_2244; // @[decode.scala 388:41]
  wire  _GEN_6396 = _T_3 ? _GEN_5748 : _GEN_2245; // @[decode.scala 388:41]
  wire  _GEN_6397 = _T_3 ? _GEN_5749 : _GEN_2246; // @[decode.scala 388:41]
  wire  _GEN_6398 = _T_3 ? _GEN_5750 : _GEN_2247; // @[decode.scala 388:41]
  wire  _GEN_6399 = _T_3 ? _GEN_5751 : _GEN_2248; // @[decode.scala 388:41]
  wire  _GEN_6400 = _T_3 ? _GEN_5752 : _GEN_2249; // @[decode.scala 388:41]
  wire  _GEN_6401 = _T_3 ? _GEN_5753 : _GEN_2250; // @[decode.scala 388:41]
  wire  _GEN_6402 = _T_3 ? _GEN_5754 : _GEN_2251; // @[decode.scala 388:41]
  wire  _GEN_6403 = _T_3 ? _GEN_5755 : _GEN_2252; // @[decode.scala 388:41]
  wire  _GEN_6404 = _T_3 ? _GEN_5756 : _GEN_2253; // @[decode.scala 388:41]
  wire  _GEN_6405 = _T_3 ? _GEN_5757 : _GEN_2254; // @[decode.scala 388:41]
  wire  _GEN_6406 = _T_3 ? _GEN_5758 : _GEN_2255; // @[decode.scala 388:41]
  wire  _GEN_6407 = _T_3 ? _GEN_5759 : _GEN_2256; // @[decode.scala 388:41]
  wire  _GEN_6408 = _T_3 ? _GEN_5760 : _GEN_2257; // @[decode.scala 388:41]
  wire  _GEN_6409 = _T_3 ? _GEN_5761 : _GEN_2258; // @[decode.scala 388:41]
  wire  _GEN_6410 = _T_3 ? _GEN_5762 : _GEN_2259; // @[decode.scala 388:41]
  wire  _GEN_6411 = _T_3 ? _GEN_5763 : _GEN_2260; // @[decode.scala 388:41]
  wire  _GEN_6412 = _T_3 ? _GEN_5764 : _GEN_2261; // @[decode.scala 388:41]
  wire  _GEN_6413 = _T_3 ? _GEN_5765 : _GEN_2262; // @[decode.scala 388:41]
  wire  _GEN_6414 = _T_3 ? _GEN_5766 : _GEN_2263; // @[decode.scala 388:41]
  wire  _GEN_6415 = _T_3 ? _GEN_5767 : _GEN_2264; // @[decode.scala 388:41]
  wire  _GEN_6416 = _T_3 ? _GEN_5768 : _GEN_2265; // @[decode.scala 388:41]
  wire  _GEN_6417 = _T_3 ? _GEN_5769 : _GEN_2266; // @[decode.scala 388:41]
  wire  _GEN_6418 = _T_3 ? _GEN_5770 : _GEN_2267; // @[decode.scala 388:41]
  wire  _GEN_6419 = _T_3 ? _GEN_5771 : _GEN_2268; // @[decode.scala 388:41]
  wire  _GEN_6420 = _T_3 ? _GEN_5772 : _GEN_2269; // @[decode.scala 388:41]
  wire  _GEN_6421 = _T_3 ? _GEN_5773 : _GEN_2270; // @[decode.scala 388:41]
  wire  _GEN_6422 = _T_3 ? _GEN_5774 : _GEN_2271; // @[decode.scala 388:41]
  wire  _GEN_6423 = _T_3 ? _GEN_5775 : _GEN_2272; // @[decode.scala 388:41]
  wire  _GEN_6424 = _T_3 ? _GEN_5776 : _GEN_2273; // @[decode.scala 388:41]
  wire  _GEN_6425 = _T_3 ? _GEN_5777 : _GEN_2274; // @[decode.scala 388:41]
  wire  _GEN_6426 = _T_3 ? _GEN_5778 : _GEN_2275; // @[decode.scala 388:41]
  wire  _GEN_6427 = _T_3 ? _GEN_5779 : _GEN_2276; // @[decode.scala 388:41]
  wire  _GEN_6428 = _T_3 ? _GEN_5780 : _GEN_2277; // @[decode.scala 388:41]
  wire  _GEN_6429 = _T_3 ? _GEN_5781 : _GEN_2278; // @[decode.scala 388:41]
  wire  _GEN_6430 = _T_3 ? _GEN_5782 : _GEN_2279; // @[decode.scala 388:41]
  wire  _GEN_6431 = _T_3 ? _GEN_5783 : _GEN_2280; // @[decode.scala 388:41]
  wire  _GEN_6432 = _T_3 ? _GEN_5784 : _GEN_2281; // @[decode.scala 388:41]
  wire  _GEN_6433 = _T_3 ? _GEN_5785 : _GEN_2282; // @[decode.scala 388:41]
  wire  _GEN_6434 = _T_3 ? _GEN_5786 : _GEN_2283; // @[decode.scala 388:41]
  wire  _GEN_6435 = _T_3 ? _GEN_5787 : _GEN_2284; // @[decode.scala 388:41]
  wire  _GEN_6436 = _T_3 ? _GEN_5788 : _GEN_2285; // @[decode.scala 388:41]
  wire  _GEN_6437 = _T_3 ? _GEN_5789 : _GEN_2286; // @[decode.scala 388:41]
  wire  _GEN_6438 = _T_3 ? _GEN_5790 : _GEN_2287; // @[decode.scala 388:41]
  wire  _GEN_6439 = _T_3 ? _GEN_5791 : _GEN_2288; // @[decode.scala 388:41]
  wire  _GEN_6440 = _T_3 ? _GEN_5792 : _GEN_2289; // @[decode.scala 388:41]
  wire  _GEN_6441 = _T_3 ? _GEN_5793 : _GEN_2290; // @[decode.scala 388:41]
  wire  _GEN_6442 = _T_3 ? _GEN_5794 : _GEN_2291; // @[decode.scala 388:41]
  wire  _GEN_6443 = _T_3 ? _GEN_5795 : _GEN_2292; // @[decode.scala 388:41]
  wire  _GEN_6444 = _T_3 ? _GEN_5796 : _GEN_2293; // @[decode.scala 388:41]
  wire  _GEN_6445 = _T_3 ? _GEN_5797 : _GEN_2294; // @[decode.scala 388:41]
  wire  _GEN_6446 = _T_3 ? _GEN_5798 : _GEN_2295; // @[decode.scala 388:41]
  wire  _GEN_6447 = _T_3 ? _GEN_5799 : _GEN_2296; // @[decode.scala 388:41]
  wire  _GEN_6448 = _T_3 ? _GEN_5800 : _GEN_2297; // @[decode.scala 388:41]
  wire  _GEN_6449 = _T_3 ? _GEN_5801 : _GEN_2298; // @[decode.scala 388:41]
  wire  _GEN_6450 = _T_3 ? _GEN_5802 : _GEN_2299; // @[decode.scala 388:41]
  wire  _GEN_6451 = _T_3 ? _GEN_5803 : _GEN_2300; // @[decode.scala 388:41]
  wire  _GEN_6452 = _T_3 ? _GEN_5804 : _GEN_2301; // @[decode.scala 388:41]
  wire  _GEN_6453 = _T_3 ? _GEN_5805 : _GEN_2302; // @[decode.scala 388:41]
  wire  _GEN_6551 = _T_3 ? _GEN_5903 : reservedFreeList4_0; // @[decode.scala 318:30 388:41]
  wire  _GEN_6552 = _T_3 ? _GEN_5904 : reservedFreeList4_1; // @[decode.scala 318:30 388:41]
  wire  _GEN_6553 = _T_3 ? _GEN_5905 : reservedFreeList4_2; // @[decode.scala 318:30 388:41]
  wire  _GEN_6554 = _T_3 ? _GEN_5906 : reservedFreeList4_3; // @[decode.scala 318:30 388:41]
  wire  _GEN_6555 = _T_3 ? _GEN_5907 : reservedFreeList4_4; // @[decode.scala 318:30 388:41]
  wire  _GEN_6556 = _T_3 ? _GEN_5908 : reservedFreeList4_5; // @[decode.scala 318:30 388:41]
  wire  _GEN_6557 = _T_3 ? _GEN_5909 : reservedFreeList4_6; // @[decode.scala 318:30 388:41]
  wire  _GEN_6558 = _T_3 ? _GEN_5910 : reservedFreeList4_7; // @[decode.scala 318:30 388:41]
  wire  _GEN_6559 = _T_3 ? _GEN_5911 : reservedFreeList4_8; // @[decode.scala 318:30 388:41]
  wire  _GEN_6560 = _T_3 ? _GEN_5912 : reservedFreeList4_9; // @[decode.scala 318:30 388:41]
  wire  _GEN_6561 = _T_3 ? _GEN_5913 : reservedFreeList4_10; // @[decode.scala 318:30 388:41]
  wire  _GEN_6562 = _T_3 ? _GEN_5914 : reservedFreeList4_11; // @[decode.scala 318:30 388:41]
  wire  _GEN_6563 = _T_3 ? _GEN_5915 : reservedFreeList4_12; // @[decode.scala 318:30 388:41]
  wire  _GEN_6564 = _T_3 ? _GEN_5916 : reservedFreeList4_13; // @[decode.scala 318:30 388:41]
  wire  _GEN_6565 = _T_3 ? _GEN_5917 : reservedFreeList4_14; // @[decode.scala 318:30 388:41]
  wire  _GEN_6566 = _T_3 ? _GEN_5918 : reservedFreeList4_15; // @[decode.scala 318:30 388:41]
  wire  _GEN_6567 = _T_3 ? _GEN_5919 : reservedFreeList4_16; // @[decode.scala 318:30 388:41]
  wire  _GEN_6568 = _T_3 ? _GEN_5920 : reservedFreeList4_17; // @[decode.scala 318:30 388:41]
  wire  _GEN_6569 = _T_3 ? _GEN_5921 : reservedFreeList4_18; // @[decode.scala 318:30 388:41]
  wire  _GEN_6570 = _T_3 ? _GEN_5922 : reservedFreeList4_19; // @[decode.scala 318:30 388:41]
  wire  _GEN_6571 = _T_3 ? _GEN_5923 : reservedFreeList4_20; // @[decode.scala 318:30 388:41]
  wire  _GEN_6572 = _T_3 ? _GEN_5924 : reservedFreeList4_21; // @[decode.scala 318:30 388:41]
  wire  _GEN_6573 = _T_3 ? _GEN_5925 : reservedFreeList4_22; // @[decode.scala 318:30 388:41]
  wire  _GEN_6574 = _T_3 ? _GEN_5926 : reservedFreeList4_23; // @[decode.scala 318:30 388:41]
  wire  _GEN_6575 = _T_3 ? _GEN_5927 : reservedFreeList4_24; // @[decode.scala 318:30 388:41]
  wire  _GEN_6576 = _T_3 ? _GEN_5928 : reservedFreeList4_25; // @[decode.scala 318:30 388:41]
  wire  _GEN_6577 = _T_3 ? _GEN_5929 : reservedFreeList4_26; // @[decode.scala 318:30 388:41]
  wire  _GEN_6578 = _T_3 ? _GEN_5930 : reservedFreeList4_27; // @[decode.scala 318:30 388:41]
  wire  _GEN_6579 = _T_3 ? _GEN_5931 : reservedFreeList4_28; // @[decode.scala 318:30 388:41]
  wire  _GEN_6580 = _T_3 ? _GEN_5932 : reservedFreeList4_29; // @[decode.scala 318:30 388:41]
  wire  _GEN_6581 = _T_3 ? _GEN_5933 : reservedFreeList4_30; // @[decode.scala 318:30 388:41]
  wire  _GEN_6582 = _T_3 ? _GEN_5934 : reservedFreeList4_31; // @[decode.scala 318:30 388:41]
  wire  _GEN_6583 = _T_3 ? _GEN_5935 : reservedFreeList4_32; // @[decode.scala 318:30 388:41]
  wire  _GEN_6584 = _T_3 ? _GEN_5936 : reservedFreeList4_33; // @[decode.scala 318:30 388:41]
  wire  _GEN_6585 = _T_3 ? _GEN_5937 : reservedFreeList4_34; // @[decode.scala 318:30 388:41]
  wire  _GEN_6586 = _T_3 ? _GEN_5938 : reservedFreeList4_35; // @[decode.scala 318:30 388:41]
  wire  _GEN_6587 = _T_3 ? _GEN_5939 : reservedFreeList4_36; // @[decode.scala 318:30 388:41]
  wire  _GEN_6588 = _T_3 ? _GEN_5940 : reservedFreeList4_37; // @[decode.scala 318:30 388:41]
  wire  _GEN_6589 = _T_3 ? _GEN_5941 : reservedFreeList4_38; // @[decode.scala 318:30 388:41]
  wire  _GEN_6590 = _T_3 ? _GEN_5942 : reservedFreeList4_39; // @[decode.scala 318:30 388:41]
  wire  _GEN_6591 = _T_3 ? _GEN_5943 : reservedFreeList4_40; // @[decode.scala 318:30 388:41]
  wire  _GEN_6592 = _T_3 ? _GEN_5944 : reservedFreeList4_41; // @[decode.scala 318:30 388:41]
  wire  _GEN_6593 = _T_3 ? _GEN_5945 : reservedFreeList4_42; // @[decode.scala 318:30 388:41]
  wire  _GEN_6594 = _T_3 ? _GEN_5946 : reservedFreeList4_43; // @[decode.scala 318:30 388:41]
  wire  _GEN_6595 = _T_3 ? _GEN_5947 : reservedFreeList4_44; // @[decode.scala 318:30 388:41]
  wire  _GEN_6596 = _T_3 ? _GEN_5948 : reservedFreeList4_45; // @[decode.scala 318:30 388:41]
  wire  _GEN_6597 = _T_3 ? _GEN_5949 : reservedFreeList4_46; // @[decode.scala 318:30 388:41]
  wire  _GEN_6598 = _T_3 ? _GEN_5950 : reservedFreeList4_47; // @[decode.scala 318:30 388:41]
  wire  _GEN_6599 = _T_3 ? _GEN_5951 : reservedFreeList4_48; // @[decode.scala 318:30 388:41]
  wire  _GEN_6600 = _T_3 ? _GEN_5952 : reservedFreeList4_49; // @[decode.scala 318:30 388:41]
  wire  _GEN_6601 = _T_3 ? _GEN_5953 : reservedFreeList4_50; // @[decode.scala 318:30 388:41]
  wire  _GEN_6602 = _T_3 ? _GEN_5954 : reservedFreeList4_51; // @[decode.scala 318:30 388:41]
  wire  _GEN_6603 = _T_3 ? _GEN_5955 : reservedFreeList4_52; // @[decode.scala 318:30 388:41]
  wire  _GEN_6604 = _T_3 ? _GEN_5956 : reservedFreeList4_53; // @[decode.scala 318:30 388:41]
  wire  _GEN_6605 = _T_3 ? _GEN_5957 : reservedFreeList4_54; // @[decode.scala 318:30 388:41]
  wire  _GEN_6606 = _T_3 ? _GEN_5958 : reservedFreeList4_55; // @[decode.scala 318:30 388:41]
  wire  _GEN_6607 = _T_3 ? _GEN_5959 : reservedFreeList4_56; // @[decode.scala 318:30 388:41]
  wire  _GEN_6608 = _T_3 ? _GEN_5960 : reservedFreeList4_57; // @[decode.scala 318:30 388:41]
  wire  _GEN_6609 = _T_3 ? _GEN_5961 : reservedFreeList4_58; // @[decode.scala 318:30 388:41]
  wire  _GEN_6610 = _T_3 ? _GEN_5962 : reservedFreeList4_59; // @[decode.scala 318:30 388:41]
  wire  _GEN_6611 = _T_3 ? _GEN_5963 : reservedFreeList4_60; // @[decode.scala 318:30 388:41]
  wire  _GEN_6612 = _T_3 ? _GEN_5964 : reservedFreeList4_61; // @[decode.scala 318:30 388:41]
  wire  _GEN_6613 = _T_3 ? _GEN_5965 : reservedFreeList4_62; // @[decode.scala 318:30 388:41]
  wire  _T_212 = fromFetch_expected_pc == fromFetch_pc; // @[decode.scala 455:71]
  wire [63:0] _GEN_6681 = _fromFetch_expected_valid_T & fromFetch_fired & fromFetch_expected_pc == fromFetch_pc ? 64'h0
     : _GEN_1855; // @[decode.scala 455:89 456:16]
  wire  isCSR = csrIns & toExec_fired; // @[decode.scala 462:98]
  reg [63:0] ustatus; // @[decode.scala 464:28]
  reg [63:0] utvec; // @[decode.scala 465:28]
  reg [63:0] uepc; // @[decode.scala 466:28]
  reg [63:0] ucause; // @[decode.scala 467:28]
  reg [63:0] scounteren; // @[decode.scala 468:28]
  reg [63:0] satp; // @[decode.scala 469:28]
  reg [63:0] mstatus; // @[decode.scala 470:28]
  reg [63:0] misa; // @[decode.scala 471:28]
  reg [63:0] medeleg; // @[decode.scala 472:28]
  reg [63:0] mideleg; // @[decode.scala 473:28]
  reg [63:0] mie; // @[decode.scala 474:28]
  reg [63:0] mtvec; // @[decode.scala 475:28]
  reg [63:0] mcounteren; // @[decode.scala 476:28]
  reg [63:0] mscratch; // @[decode.scala 477:28]
  reg [63:0] mepc; // @[decode.scala 478:28]
  reg [63:0] mcause; // @[decode.scala 479:28]
  reg [63:0] mtval; // @[decode.scala 480:28]
  reg [63:0] mip; // @[decode.scala 481:28]
  reg [63:0] pmpcfg0; // @[decode.scala 482:28]
  reg [63:0] pmpaddr0; // @[decode.scala 483:28]
  reg [63:0] mvendorid; // @[decode.scala 484:28]
  reg [63:0] marchid; // @[decode.scala 485:28]
  reg [63:0] mimpid; // @[decode.scala 486:28]
  reg [63:0] mhartid; // @[decode.scala 487:28]
  wire [63:0] _mstatus_T = mstatus & 64'h1888; // @[decode.scala 489:23]
  wire [63:0] _mstatus_T_1 = _mstatus_T | 64'ha00000000; // @[decode.scala 489:48]
  wire [63:0] _GEN_6686 = isCSR ? outputBuffer_immediate : {{52'd0}, csrAddrReg}; // @[decode.scala 492:15 495:19 236:27]
  wire  _T_214 = opcode == 7'h73; // @[decode.scala 501:15]
  wire [63:0] _T_219 = immediate_immediate & 64'hfff; // @[decode.scala 502:22]
  wire [63:0] _GEN_6689 = 64'hf14 == _T_219 ? mhartid : csrReadDataReg; // @[decode.scala 234:31 502:34 526:37]
  wire [63:0] _GEN_6690 = 64'hf13 == _T_219 ? mimpid : _GEN_6689; // @[decode.scala 502:34 525:37]
  wire [63:0] _GEN_6691 = 64'hf12 == _T_219 ? marchid : _GEN_6690; // @[decode.scala 502:34 524:37]
  wire [63:0] _GEN_6692 = 64'hf11 == _T_219 ? mvendorid : _GEN_6691; // @[decode.scala 502:34 523:37]
  wire [63:0] _GEN_6693 = 64'h3b0 == _T_219 ? pmpaddr0 : _GEN_6692; // @[decode.scala 502:34 522:37]
  wire [63:0] _GEN_6694 = 64'h3a0 == _T_219 ? pmpcfg0 : _GEN_6693; // @[decode.scala 502:34 521:37]
  wire [63:0] _GEN_6695 = 64'h344 == _T_219 ? mip : _GEN_6694; // @[decode.scala 502:34 520:37]
  wire [63:0] _GEN_6696 = 64'h343 == _T_219 ? mtval : _GEN_6695; // @[decode.scala 502:34 519:37]
  wire [63:0] _GEN_6697 = 64'h342 == _T_219 ? mcause : _GEN_6696; // @[decode.scala 502:34 518:37]
  wire [63:0] _GEN_6698 = 64'h341 == _T_219 ? mepc : _GEN_6697; // @[decode.scala 502:34 517:37]
  wire [63:0] _GEN_6699 = 64'h340 == _T_219 ? mscratch : _GEN_6698; // @[decode.scala 502:34 516:37]
  wire [63:0] _GEN_6700 = 64'h306 == _T_219 ? mcounteren : _GEN_6699; // @[decode.scala 502:34 515:37]
  wire [63:0] _GEN_6701 = 64'h305 == _T_219 ? mtvec : _GEN_6700; // @[decode.scala 502:34 514:37]
  wire [63:0] _GEN_6702 = 64'h304 == _T_219 ? mie : _GEN_6701; // @[decode.scala 502:34 513:37]
  wire [63:0] _GEN_6703 = 64'h303 == _T_219 ? mideleg : _GEN_6702; // @[decode.scala 502:34 512:37]
  wire [63:0] _GEN_6704 = 64'h302 == _T_219 ? medeleg : _GEN_6703; // @[decode.scala 502:34 511:37]
  wire [63:0] _GEN_6705 = 64'h301 == _T_219 ? misa : _GEN_6704; // @[decode.scala 502:34 510:37]
  wire [63:0] _GEN_6706 = 64'h300 == _T_219 ? mstatus : _GEN_6705; // @[decode.scala 502:34 509:37]
  wire [63:0] _GEN_6707 = 64'h180 == _T_219 ? satp : _GEN_6706; // @[decode.scala 502:34 508:37]
  wire [63:0] _GEN_6708 = 64'h106 == _T_219 ? scounteren : _GEN_6707; // @[decode.scala 502:34 507:37]
  wire [63:0] _GEN_6709 = 64'h42 == _T_219 ? ucause : _GEN_6708; // @[decode.scala 502:34 506:37]
  wire [63:0] _GEN_6710 = 64'h41 == _T_219 ? uepc : _GEN_6709; // @[decode.scala 502:34 505:37]
  wire  _T_246 = writeBackResult_fired & writeBackResult_instruction[6:0] == 7'h73; // @[decode.scala 531:30]
  wire  _GEN_6714 = writeBackResult_fired & writeBackResult_instruction[6:0] == 7'h73 ? 1'h0 : _GEN_4; // @[decode.scala 531:80 532:14]
  wire  _T_256 = 12'h0 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_257 = 12'h5 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_258 = 12'h41 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_259 = 12'h42 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_260 = 12'h106 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_261 = 12'h180 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_262 = 12'h300 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_263 = 12'h301 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_264 = 12'h302 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_265 = 12'h303 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_266 = 12'h304 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_267 = 12'h305 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_268 = 12'h306 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_269 = 12'h340 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_270 = 12'h341 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_271 = 12'h342 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_272 = 12'h343 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_273 = 12'h344 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_274 = 12'h3a0 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_275 = 12'h3b0 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_276 = 12'hf11 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_277 = 12'hf12 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_278 = 12'hf13 == csrAddrReg; // @[decode.scala 540:39]
  wire  _T_279 = 12'hf14 == csrAddrReg; // @[decode.scala 540:39]
  wire [63:0] csrWriteData = _T_246 & writeBackResult_instruction[14:12] != 3'h0 ? writeBackResult_data : 64'h0; // @[decode.scala 535:126 537:18]
  wire [63:0] _GEN_6715 = 12'hf14 == csrAddrReg ? csrWriteData : mhartid; // @[decode.scala 487:28 540:39 564:37]
  wire [63:0] _GEN_6716 = 12'hf13 == csrAddrReg ? csrWriteData : mimpid; // @[decode.scala 486:28 540:39 563:37]
  wire [63:0] _GEN_6717 = 12'hf13 == csrAddrReg ? mhartid : _GEN_6715; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6718 = 12'hf12 == csrAddrReg ? csrWriteData : marchid; // @[decode.scala 485:28 540:39 562:37]
  wire [63:0] _GEN_6719 = 12'hf12 == csrAddrReg ? mimpid : _GEN_6716; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6720 = 12'hf12 == csrAddrReg ? mhartid : _GEN_6717; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6721 = 12'hf11 == csrAddrReg ? csrWriteData : mvendorid; // @[decode.scala 484:28 540:39 561:37]
  wire [63:0] _GEN_6722 = 12'hf11 == csrAddrReg ? marchid : _GEN_6718; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6723 = 12'hf11 == csrAddrReg ? mimpid : _GEN_6719; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6724 = 12'hf11 == csrAddrReg ? mhartid : _GEN_6720; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6725 = 12'h3b0 == csrAddrReg ? csrWriteData : pmpaddr0; // @[decode.scala 483:28 540:39 560:37]
  wire [63:0] _GEN_6726 = 12'h3b0 == csrAddrReg ? mvendorid : _GEN_6721; // @[decode.scala 484:28 540:39]
  wire [63:0] _GEN_6727 = 12'h3b0 == csrAddrReg ? marchid : _GEN_6722; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6728 = 12'h3b0 == csrAddrReg ? mimpid : _GEN_6723; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6729 = 12'h3b0 == csrAddrReg ? mhartid : _GEN_6724; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6730 = 12'h3a0 == csrAddrReg ? csrWriteData : pmpcfg0; // @[decode.scala 482:28 540:39 559:37]
  wire [63:0] _GEN_6731 = 12'h3a0 == csrAddrReg ? pmpaddr0 : _GEN_6725; // @[decode.scala 483:28 540:39]
  wire [63:0] _GEN_6732 = 12'h3a0 == csrAddrReg ? mvendorid : _GEN_6726; // @[decode.scala 484:28 540:39]
  wire [63:0] _GEN_6733 = 12'h3a0 == csrAddrReg ? marchid : _GEN_6727; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6734 = 12'h3a0 == csrAddrReg ? mimpid : _GEN_6728; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6735 = 12'h3a0 == csrAddrReg ? mhartid : _GEN_6729; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6736 = 12'h344 == csrAddrReg ? csrWriteData : mip; // @[decode.scala 481:28 540:39 558:37]
  wire [63:0] _GEN_6737 = 12'h344 == csrAddrReg ? pmpcfg0 : _GEN_6730; // @[decode.scala 482:28 540:39]
  wire [63:0] _GEN_6738 = 12'h344 == csrAddrReg ? pmpaddr0 : _GEN_6731; // @[decode.scala 483:28 540:39]
  wire [63:0] _GEN_6739 = 12'h344 == csrAddrReg ? mvendorid : _GEN_6732; // @[decode.scala 484:28 540:39]
  wire [63:0] _GEN_6740 = 12'h344 == csrAddrReg ? marchid : _GEN_6733; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6741 = 12'h344 == csrAddrReg ? mimpid : _GEN_6734; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6742 = 12'h344 == csrAddrReg ? mhartid : _GEN_6735; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6743 = 12'h343 == csrAddrReg ? csrWriteData : mtval; // @[decode.scala 480:28 540:39 557:37]
  wire [63:0] _GEN_6744 = 12'h343 == csrAddrReg ? mip : _GEN_6736; // @[decode.scala 481:28 540:39]
  wire [63:0] _GEN_6745 = 12'h343 == csrAddrReg ? pmpcfg0 : _GEN_6737; // @[decode.scala 482:28 540:39]
  wire [63:0] _GEN_6746 = 12'h343 == csrAddrReg ? pmpaddr0 : _GEN_6738; // @[decode.scala 483:28 540:39]
  wire [63:0] _GEN_6747 = 12'h343 == csrAddrReg ? mvendorid : _GEN_6739; // @[decode.scala 484:28 540:39]
  wire [63:0] _GEN_6748 = 12'h343 == csrAddrReg ? marchid : _GEN_6740; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6749 = 12'h343 == csrAddrReg ? mimpid : _GEN_6741; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6750 = 12'h343 == csrAddrReg ? mhartid : _GEN_6742; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6751 = 12'h342 == csrAddrReg ? csrWriteData : mcause; // @[decode.scala 479:28 540:39 556:37]
  wire [63:0] _GEN_6752 = 12'h342 == csrAddrReg ? mtval : _GEN_6743; // @[decode.scala 480:28 540:39]
  wire [63:0] _GEN_6753 = 12'h342 == csrAddrReg ? mip : _GEN_6744; // @[decode.scala 481:28 540:39]
  wire [63:0] _GEN_6754 = 12'h342 == csrAddrReg ? pmpcfg0 : _GEN_6745; // @[decode.scala 482:28 540:39]
  wire [63:0] _GEN_6755 = 12'h342 == csrAddrReg ? pmpaddr0 : _GEN_6746; // @[decode.scala 483:28 540:39]
  wire [63:0] _GEN_6756 = 12'h342 == csrAddrReg ? mvendorid : _GEN_6747; // @[decode.scala 484:28 540:39]
  wire [63:0] _GEN_6757 = 12'h342 == csrAddrReg ? marchid : _GEN_6748; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6758 = 12'h342 == csrAddrReg ? mimpid : _GEN_6749; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6759 = 12'h342 == csrAddrReg ? mhartid : _GEN_6750; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6760 = 12'h341 == csrAddrReg ? csrWriteData : mepc; // @[decode.scala 478:28 540:39 555:37]
  wire [63:0] _GEN_6761 = 12'h341 == csrAddrReg ? mcause : _GEN_6751; // @[decode.scala 479:28 540:39]
  wire [63:0] _GEN_6762 = 12'h341 == csrAddrReg ? mtval : _GEN_6752; // @[decode.scala 480:28 540:39]
  wire [63:0] _GEN_6763 = 12'h341 == csrAddrReg ? mip : _GEN_6753; // @[decode.scala 481:28 540:39]
  wire [63:0] _GEN_6764 = 12'h341 == csrAddrReg ? pmpcfg0 : _GEN_6754; // @[decode.scala 482:28 540:39]
  wire [63:0] _GEN_6765 = 12'h341 == csrAddrReg ? pmpaddr0 : _GEN_6755; // @[decode.scala 483:28 540:39]
  wire [63:0] _GEN_6766 = 12'h341 == csrAddrReg ? mvendorid : _GEN_6756; // @[decode.scala 484:28 540:39]
  wire [63:0] _GEN_6767 = 12'h341 == csrAddrReg ? marchid : _GEN_6757; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6768 = 12'h341 == csrAddrReg ? mimpid : _GEN_6758; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6769 = 12'h341 == csrAddrReg ? mhartid : _GEN_6759; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6770 = 12'h340 == csrAddrReg ? csrWriteData : mscratch; // @[decode.scala 477:28 540:39 554:37]
  wire [63:0] _GEN_6771 = 12'h340 == csrAddrReg ? mepc : _GEN_6760; // @[decode.scala 478:28 540:39]
  wire [63:0] _GEN_6772 = 12'h340 == csrAddrReg ? mcause : _GEN_6761; // @[decode.scala 479:28 540:39]
  wire [63:0] _GEN_6773 = 12'h340 == csrAddrReg ? mtval : _GEN_6762; // @[decode.scala 480:28 540:39]
  wire [63:0] _GEN_6774 = 12'h340 == csrAddrReg ? mip : _GEN_6763; // @[decode.scala 481:28 540:39]
  wire [63:0] _GEN_6775 = 12'h340 == csrAddrReg ? pmpcfg0 : _GEN_6764; // @[decode.scala 482:28 540:39]
  wire [63:0] _GEN_6776 = 12'h340 == csrAddrReg ? pmpaddr0 : _GEN_6765; // @[decode.scala 483:28 540:39]
  wire [63:0] _GEN_6777 = 12'h340 == csrAddrReg ? mvendorid : _GEN_6766; // @[decode.scala 484:28 540:39]
  wire [63:0] _GEN_6778 = 12'h340 == csrAddrReg ? marchid : _GEN_6767; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6779 = 12'h340 == csrAddrReg ? mimpid : _GEN_6768; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6780 = 12'h340 == csrAddrReg ? mhartid : _GEN_6769; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6781 = 12'h306 == csrAddrReg ? csrWriteData : mcounteren; // @[decode.scala 476:28 540:39 553:37]
  wire [63:0] _GEN_6782 = 12'h306 == csrAddrReg ? mscratch : _GEN_6770; // @[decode.scala 477:28 540:39]
  wire [63:0] _GEN_6783 = 12'h306 == csrAddrReg ? mepc : _GEN_6771; // @[decode.scala 478:28 540:39]
  wire [63:0] _GEN_6784 = 12'h306 == csrAddrReg ? mcause : _GEN_6772; // @[decode.scala 479:28 540:39]
  wire [63:0] _GEN_6785 = 12'h306 == csrAddrReg ? mtval : _GEN_6773; // @[decode.scala 480:28 540:39]
  wire [63:0] _GEN_6786 = 12'h306 == csrAddrReg ? mip : _GEN_6774; // @[decode.scala 481:28 540:39]
  wire [63:0] _GEN_6787 = 12'h306 == csrAddrReg ? pmpcfg0 : _GEN_6775; // @[decode.scala 482:28 540:39]
  wire [63:0] _GEN_6788 = 12'h306 == csrAddrReg ? pmpaddr0 : _GEN_6776; // @[decode.scala 483:28 540:39]
  wire [63:0] _GEN_6789 = 12'h306 == csrAddrReg ? mvendorid : _GEN_6777; // @[decode.scala 484:28 540:39]
  wire [63:0] _GEN_6790 = 12'h306 == csrAddrReg ? marchid : _GEN_6778; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6791 = 12'h306 == csrAddrReg ? mimpid : _GEN_6779; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6792 = 12'h306 == csrAddrReg ? mhartid : _GEN_6780; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6793 = 12'h305 == csrAddrReg ? csrWriteData : mtvec; // @[decode.scala 475:28 540:39 552:37]
  wire [63:0] _GEN_6794 = 12'h305 == csrAddrReg ? mcounteren : _GEN_6781; // @[decode.scala 476:28 540:39]
  wire [63:0] _GEN_6795 = 12'h305 == csrAddrReg ? mscratch : _GEN_6782; // @[decode.scala 477:28 540:39]
  wire [63:0] _GEN_6796 = 12'h305 == csrAddrReg ? mepc : _GEN_6783; // @[decode.scala 478:28 540:39]
  wire [63:0] _GEN_6797 = 12'h305 == csrAddrReg ? mcause : _GEN_6784; // @[decode.scala 479:28 540:39]
  wire [63:0] _GEN_6798 = 12'h305 == csrAddrReg ? mtval : _GEN_6785; // @[decode.scala 480:28 540:39]
  wire [63:0] _GEN_6799 = 12'h305 == csrAddrReg ? mip : _GEN_6786; // @[decode.scala 481:28 540:39]
  wire [63:0] _GEN_6800 = 12'h305 == csrAddrReg ? pmpcfg0 : _GEN_6787; // @[decode.scala 482:28 540:39]
  wire [63:0] _GEN_6801 = 12'h305 == csrAddrReg ? pmpaddr0 : _GEN_6788; // @[decode.scala 483:28 540:39]
  wire [63:0] _GEN_6802 = 12'h305 == csrAddrReg ? mvendorid : _GEN_6789; // @[decode.scala 484:28 540:39]
  wire [63:0] _GEN_6803 = 12'h305 == csrAddrReg ? marchid : _GEN_6790; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6804 = 12'h305 == csrAddrReg ? mimpid : _GEN_6791; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6805 = 12'h305 == csrAddrReg ? mhartid : _GEN_6792; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6806 = 12'h304 == csrAddrReg ? csrWriteData : mie; // @[decode.scala 474:28 540:39 551:37]
  wire [63:0] _GEN_6807 = 12'h304 == csrAddrReg ? mtvec : _GEN_6793; // @[decode.scala 475:28 540:39]
  wire [63:0] _GEN_6808 = 12'h304 == csrAddrReg ? mcounteren : _GEN_6794; // @[decode.scala 476:28 540:39]
  wire [63:0] _GEN_6809 = 12'h304 == csrAddrReg ? mscratch : _GEN_6795; // @[decode.scala 477:28 540:39]
  wire [63:0] _GEN_6810 = 12'h304 == csrAddrReg ? mepc : _GEN_6796; // @[decode.scala 478:28 540:39]
  wire [63:0] _GEN_6811 = 12'h304 == csrAddrReg ? mcause : _GEN_6797; // @[decode.scala 479:28 540:39]
  wire [63:0] _GEN_6812 = 12'h304 == csrAddrReg ? mtval : _GEN_6798; // @[decode.scala 480:28 540:39]
  wire [63:0] _GEN_6813 = 12'h304 == csrAddrReg ? mip : _GEN_6799; // @[decode.scala 481:28 540:39]
  wire [63:0] _GEN_6814 = 12'h304 == csrAddrReg ? pmpcfg0 : _GEN_6800; // @[decode.scala 482:28 540:39]
  wire [63:0] _GEN_6815 = 12'h304 == csrAddrReg ? pmpaddr0 : _GEN_6801; // @[decode.scala 483:28 540:39]
  wire [63:0] _GEN_6816 = 12'h304 == csrAddrReg ? mvendorid : _GEN_6802; // @[decode.scala 484:28 540:39]
  wire [63:0] _GEN_6817 = 12'h304 == csrAddrReg ? marchid : _GEN_6803; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6818 = 12'h304 == csrAddrReg ? mimpid : _GEN_6804; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6819 = 12'h304 == csrAddrReg ? mhartid : _GEN_6805; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6820 = 12'h303 == csrAddrReg ? csrWriteData : mideleg; // @[decode.scala 473:28 540:39 550:37]
  wire [63:0] _GEN_6821 = 12'h303 == csrAddrReg ? mie : _GEN_6806; // @[decode.scala 474:28 540:39]
  wire [63:0] _GEN_6822 = 12'h303 == csrAddrReg ? mtvec : _GEN_6807; // @[decode.scala 475:28 540:39]
  wire [63:0] _GEN_6823 = 12'h303 == csrAddrReg ? mcounteren : _GEN_6808; // @[decode.scala 476:28 540:39]
  wire [63:0] _GEN_6824 = 12'h303 == csrAddrReg ? mscratch : _GEN_6809; // @[decode.scala 477:28 540:39]
  wire [63:0] _GEN_6825 = 12'h303 == csrAddrReg ? mepc : _GEN_6810; // @[decode.scala 478:28 540:39]
  wire [63:0] _GEN_6826 = 12'h303 == csrAddrReg ? mcause : _GEN_6811; // @[decode.scala 479:28 540:39]
  wire [63:0] _GEN_6827 = 12'h303 == csrAddrReg ? mtval : _GEN_6812; // @[decode.scala 480:28 540:39]
  wire [63:0] _GEN_6828 = 12'h303 == csrAddrReg ? mip : _GEN_6813; // @[decode.scala 481:28 540:39]
  wire [63:0] _GEN_6829 = 12'h303 == csrAddrReg ? pmpcfg0 : _GEN_6814; // @[decode.scala 482:28 540:39]
  wire [63:0] _GEN_6830 = 12'h303 == csrAddrReg ? pmpaddr0 : _GEN_6815; // @[decode.scala 483:28 540:39]
  wire [63:0] _GEN_6831 = 12'h303 == csrAddrReg ? mvendorid : _GEN_6816; // @[decode.scala 484:28 540:39]
  wire [63:0] _GEN_6832 = 12'h303 == csrAddrReg ? marchid : _GEN_6817; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6833 = 12'h303 == csrAddrReg ? mimpid : _GEN_6818; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6834 = 12'h303 == csrAddrReg ? mhartid : _GEN_6819; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6835 = 12'h302 == csrAddrReg ? csrWriteData : medeleg; // @[decode.scala 472:28 540:39 549:37]
  wire [63:0] _GEN_6836 = 12'h302 == csrAddrReg ? mideleg : _GEN_6820; // @[decode.scala 473:28 540:39]
  wire [63:0] _GEN_6837 = 12'h302 == csrAddrReg ? mie : _GEN_6821; // @[decode.scala 474:28 540:39]
  wire [63:0] _GEN_6838 = 12'h302 == csrAddrReg ? mtvec : _GEN_6822; // @[decode.scala 475:28 540:39]
  wire [63:0] _GEN_6839 = 12'h302 == csrAddrReg ? mcounteren : _GEN_6823; // @[decode.scala 476:28 540:39]
  wire [63:0] _GEN_6840 = 12'h302 == csrAddrReg ? mscratch : _GEN_6824; // @[decode.scala 477:28 540:39]
  wire [63:0] _GEN_6841 = 12'h302 == csrAddrReg ? mepc : _GEN_6825; // @[decode.scala 478:28 540:39]
  wire [63:0] _GEN_6842 = 12'h302 == csrAddrReg ? mcause : _GEN_6826; // @[decode.scala 479:28 540:39]
  wire [63:0] _GEN_6843 = 12'h302 == csrAddrReg ? mtval : _GEN_6827; // @[decode.scala 480:28 540:39]
  wire [63:0] _GEN_6844 = 12'h302 == csrAddrReg ? mip : _GEN_6828; // @[decode.scala 481:28 540:39]
  wire [63:0] _GEN_6845 = 12'h302 == csrAddrReg ? pmpcfg0 : _GEN_6829; // @[decode.scala 482:28 540:39]
  wire [63:0] _GEN_6846 = 12'h302 == csrAddrReg ? pmpaddr0 : _GEN_6830; // @[decode.scala 483:28 540:39]
  wire [63:0] _GEN_6847 = 12'h302 == csrAddrReg ? mvendorid : _GEN_6831; // @[decode.scala 484:28 540:39]
  wire [63:0] _GEN_6848 = 12'h302 == csrAddrReg ? marchid : _GEN_6832; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6849 = 12'h302 == csrAddrReg ? mimpid : _GEN_6833; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6850 = 12'h302 == csrAddrReg ? mhartid : _GEN_6834; // @[decode.scala 487:28 540:39]
  wire [126:0] _GEN_6851 = 12'h301 == csrAddrReg ? {{63'd0}, csrWriteData} : 127'h8000000000101101; // @[decode.scala 540:39 548:37 490:8]
  wire [63:0] _GEN_6852 = 12'h301 == csrAddrReg ? medeleg : _GEN_6835; // @[decode.scala 472:28 540:39]
  wire [63:0] _GEN_6853 = 12'h301 == csrAddrReg ? mideleg : _GEN_6836; // @[decode.scala 473:28 540:39]
  wire [63:0] _GEN_6854 = 12'h301 == csrAddrReg ? mie : _GEN_6837; // @[decode.scala 474:28 540:39]
  wire [63:0] _GEN_6855 = 12'h301 == csrAddrReg ? mtvec : _GEN_6838; // @[decode.scala 475:28 540:39]
  wire [63:0] _GEN_6856 = 12'h301 == csrAddrReg ? mcounteren : _GEN_6839; // @[decode.scala 476:28 540:39]
  wire [63:0] _GEN_6857 = 12'h301 == csrAddrReg ? mscratch : _GEN_6840; // @[decode.scala 477:28 540:39]
  wire [63:0] _GEN_6858 = 12'h301 == csrAddrReg ? mepc : _GEN_6841; // @[decode.scala 478:28 540:39]
  wire [63:0] _GEN_6859 = 12'h301 == csrAddrReg ? mcause : _GEN_6842; // @[decode.scala 479:28 540:39]
  wire [63:0] _GEN_6860 = 12'h301 == csrAddrReg ? mtval : _GEN_6843; // @[decode.scala 480:28 540:39]
  wire [63:0] _GEN_6861 = 12'h301 == csrAddrReg ? mip : _GEN_6844; // @[decode.scala 481:28 540:39]
  wire [63:0] _GEN_6862 = 12'h301 == csrAddrReg ? pmpcfg0 : _GEN_6845; // @[decode.scala 482:28 540:39]
  wire [63:0] _GEN_6863 = 12'h301 == csrAddrReg ? pmpaddr0 : _GEN_6846; // @[decode.scala 483:28 540:39]
  wire [63:0] _GEN_6864 = 12'h301 == csrAddrReg ? mvendorid : _GEN_6847; // @[decode.scala 484:28 540:39]
  wire [63:0] _GEN_6865 = 12'h301 == csrAddrReg ? marchid : _GEN_6848; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6866 = 12'h301 == csrAddrReg ? mimpid : _GEN_6849; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6867 = 12'h301 == csrAddrReg ? mhartid : _GEN_6850; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6868 = 12'h300 == csrAddrReg ? csrWriteData : _mstatus_T_1; // @[decode.scala 489:11 540:39 547:37]
  wire [126:0] _GEN_6869 = 12'h300 == csrAddrReg ? 127'h8000000000101101 : _GEN_6851; // @[decode.scala 540:39 490:8]
  wire [63:0] _GEN_6870 = 12'h300 == csrAddrReg ? medeleg : _GEN_6852; // @[decode.scala 472:28 540:39]
  wire [63:0] _GEN_6871 = 12'h300 == csrAddrReg ? mideleg : _GEN_6853; // @[decode.scala 473:28 540:39]
  wire [63:0] _GEN_6872 = 12'h300 == csrAddrReg ? mie : _GEN_6854; // @[decode.scala 474:28 540:39]
  wire [63:0] _GEN_6873 = 12'h300 == csrAddrReg ? mtvec : _GEN_6855; // @[decode.scala 475:28 540:39]
  wire [63:0] _GEN_6874 = 12'h300 == csrAddrReg ? mcounteren : _GEN_6856; // @[decode.scala 476:28 540:39]
  wire [63:0] _GEN_6875 = 12'h300 == csrAddrReg ? mscratch : _GEN_6857; // @[decode.scala 477:28 540:39]
  wire [63:0] _GEN_6876 = 12'h300 == csrAddrReg ? mepc : _GEN_6858; // @[decode.scala 478:28 540:39]
  wire [63:0] _GEN_6877 = 12'h300 == csrAddrReg ? mcause : _GEN_6859; // @[decode.scala 479:28 540:39]
  wire [63:0] _GEN_6878 = 12'h300 == csrAddrReg ? mtval : _GEN_6860; // @[decode.scala 480:28 540:39]
  wire [63:0] _GEN_6879 = 12'h300 == csrAddrReg ? mip : _GEN_6861; // @[decode.scala 481:28 540:39]
  wire [63:0] _GEN_6880 = 12'h300 == csrAddrReg ? pmpcfg0 : _GEN_6862; // @[decode.scala 482:28 540:39]
  wire [63:0] _GEN_6881 = 12'h300 == csrAddrReg ? pmpaddr0 : _GEN_6863; // @[decode.scala 483:28 540:39]
  wire [63:0] _GEN_6882 = 12'h300 == csrAddrReg ? mvendorid : _GEN_6864; // @[decode.scala 484:28 540:39]
  wire [63:0] _GEN_6883 = 12'h300 == csrAddrReg ? marchid : _GEN_6865; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6884 = 12'h300 == csrAddrReg ? mimpid : _GEN_6866; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6885 = 12'h300 == csrAddrReg ? mhartid : _GEN_6867; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6886 = 12'h180 == csrAddrReg ? csrWriteData : satp; // @[decode.scala 469:28 540:39 546:37]
  wire [63:0] _GEN_6887 = 12'h180 == csrAddrReg ? _mstatus_T_1 : _GEN_6868; // @[decode.scala 489:11 540:39]
  wire [126:0] _GEN_6888 = 12'h180 == csrAddrReg ? 127'h8000000000101101 : _GEN_6869; // @[decode.scala 540:39 490:8]
  wire [63:0] _GEN_6889 = 12'h180 == csrAddrReg ? medeleg : _GEN_6870; // @[decode.scala 472:28 540:39]
  wire [63:0] _GEN_6890 = 12'h180 == csrAddrReg ? mideleg : _GEN_6871; // @[decode.scala 473:28 540:39]
  wire [63:0] _GEN_6891 = 12'h180 == csrAddrReg ? mie : _GEN_6872; // @[decode.scala 474:28 540:39]
  wire [63:0] _GEN_6892 = 12'h180 == csrAddrReg ? mtvec : _GEN_6873; // @[decode.scala 475:28 540:39]
  wire [63:0] _GEN_6893 = 12'h180 == csrAddrReg ? mcounteren : _GEN_6874; // @[decode.scala 476:28 540:39]
  wire [63:0] _GEN_6894 = 12'h180 == csrAddrReg ? mscratch : _GEN_6875; // @[decode.scala 477:28 540:39]
  wire [63:0] _GEN_6895 = 12'h180 == csrAddrReg ? mepc : _GEN_6876; // @[decode.scala 478:28 540:39]
  wire [63:0] _GEN_6896 = 12'h180 == csrAddrReg ? mcause : _GEN_6877; // @[decode.scala 479:28 540:39]
  wire [63:0] _GEN_6897 = 12'h180 == csrAddrReg ? mtval : _GEN_6878; // @[decode.scala 480:28 540:39]
  wire [63:0] _GEN_6898 = 12'h180 == csrAddrReg ? mip : _GEN_6879; // @[decode.scala 481:28 540:39]
  wire [63:0] _GEN_6899 = 12'h180 == csrAddrReg ? pmpcfg0 : _GEN_6880; // @[decode.scala 482:28 540:39]
  wire [63:0] _GEN_6900 = 12'h180 == csrAddrReg ? pmpaddr0 : _GEN_6881; // @[decode.scala 483:28 540:39]
  wire [63:0] _GEN_6901 = 12'h180 == csrAddrReg ? mvendorid : _GEN_6882; // @[decode.scala 484:28 540:39]
  wire [63:0] _GEN_6902 = 12'h180 == csrAddrReg ? marchid : _GEN_6883; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6903 = 12'h180 == csrAddrReg ? mimpid : _GEN_6884; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6904 = 12'h180 == csrAddrReg ? mhartid : _GEN_6885; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6905 = 12'h106 == csrAddrReg ? csrWriteData : scounteren; // @[decode.scala 468:28 540:39 545:37]
  wire [63:0] _GEN_6906 = 12'h106 == csrAddrReg ? satp : _GEN_6886; // @[decode.scala 469:28 540:39]
  wire [63:0] _GEN_6907 = 12'h106 == csrAddrReg ? _mstatus_T_1 : _GEN_6887; // @[decode.scala 489:11 540:39]
  wire [126:0] _GEN_6908 = 12'h106 == csrAddrReg ? 127'h8000000000101101 : _GEN_6888; // @[decode.scala 540:39 490:8]
  wire [63:0] _GEN_6909 = 12'h106 == csrAddrReg ? medeleg : _GEN_6889; // @[decode.scala 472:28 540:39]
  wire [63:0] _GEN_6910 = 12'h106 == csrAddrReg ? mideleg : _GEN_6890; // @[decode.scala 473:28 540:39]
  wire [63:0] _GEN_6911 = 12'h106 == csrAddrReg ? mie : _GEN_6891; // @[decode.scala 474:28 540:39]
  wire [63:0] _GEN_6912 = 12'h106 == csrAddrReg ? mtvec : _GEN_6892; // @[decode.scala 475:28 540:39]
  wire [63:0] _GEN_6913 = 12'h106 == csrAddrReg ? mcounteren : _GEN_6893; // @[decode.scala 476:28 540:39]
  wire [63:0] _GEN_6914 = 12'h106 == csrAddrReg ? mscratch : _GEN_6894; // @[decode.scala 477:28 540:39]
  wire [63:0] _GEN_6915 = 12'h106 == csrAddrReg ? mepc : _GEN_6895; // @[decode.scala 478:28 540:39]
  wire [63:0] _GEN_6916 = 12'h106 == csrAddrReg ? mcause : _GEN_6896; // @[decode.scala 479:28 540:39]
  wire [63:0] _GEN_6917 = 12'h106 == csrAddrReg ? mtval : _GEN_6897; // @[decode.scala 480:28 540:39]
  wire [63:0] _GEN_6918 = 12'h106 == csrAddrReg ? mip : _GEN_6898; // @[decode.scala 481:28 540:39]
  wire [63:0] _GEN_6919 = 12'h106 == csrAddrReg ? pmpcfg0 : _GEN_6899; // @[decode.scala 482:28 540:39]
  wire [63:0] _GEN_6920 = 12'h106 == csrAddrReg ? pmpaddr0 : _GEN_6900; // @[decode.scala 483:28 540:39]
  wire [63:0] _GEN_6921 = 12'h106 == csrAddrReg ? mvendorid : _GEN_6901; // @[decode.scala 484:28 540:39]
  wire [63:0] _GEN_6922 = 12'h106 == csrAddrReg ? marchid : _GEN_6902; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6923 = 12'h106 == csrAddrReg ? mimpid : _GEN_6903; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6924 = 12'h106 == csrAddrReg ? mhartid : _GEN_6904; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6925 = 12'h42 == csrAddrReg ? csrWriteData : ucause; // @[decode.scala 467:28 540:39 544:37]
  wire [63:0] _GEN_6926 = 12'h42 == csrAddrReg ? scounteren : _GEN_6905; // @[decode.scala 468:28 540:39]
  wire [63:0] _GEN_6927 = 12'h42 == csrAddrReg ? satp : _GEN_6906; // @[decode.scala 469:28 540:39]
  wire [63:0] _GEN_6928 = 12'h42 == csrAddrReg ? _mstatus_T_1 : _GEN_6907; // @[decode.scala 489:11 540:39]
  wire [126:0] _GEN_6929 = 12'h42 == csrAddrReg ? 127'h8000000000101101 : _GEN_6908; // @[decode.scala 540:39 490:8]
  wire [63:0] _GEN_6930 = 12'h42 == csrAddrReg ? medeleg : _GEN_6909; // @[decode.scala 472:28 540:39]
  wire [63:0] _GEN_6931 = 12'h42 == csrAddrReg ? mideleg : _GEN_6910; // @[decode.scala 473:28 540:39]
  wire [63:0] _GEN_6932 = 12'h42 == csrAddrReg ? mie : _GEN_6911; // @[decode.scala 474:28 540:39]
  wire [63:0] _GEN_6933 = 12'h42 == csrAddrReg ? mtvec : _GEN_6912; // @[decode.scala 475:28 540:39]
  wire [63:0] _GEN_6934 = 12'h42 == csrAddrReg ? mcounteren : _GEN_6913; // @[decode.scala 476:28 540:39]
  wire [63:0] _GEN_6935 = 12'h42 == csrAddrReg ? mscratch : _GEN_6914; // @[decode.scala 477:28 540:39]
  wire [63:0] _GEN_6936 = 12'h42 == csrAddrReg ? mepc : _GEN_6915; // @[decode.scala 478:28 540:39]
  wire [63:0] _GEN_6937 = 12'h42 == csrAddrReg ? mcause : _GEN_6916; // @[decode.scala 479:28 540:39]
  wire [63:0] _GEN_6938 = 12'h42 == csrAddrReg ? mtval : _GEN_6917; // @[decode.scala 480:28 540:39]
  wire [63:0] _GEN_6939 = 12'h42 == csrAddrReg ? mip : _GEN_6918; // @[decode.scala 481:28 540:39]
  wire [63:0] _GEN_6940 = 12'h42 == csrAddrReg ? pmpcfg0 : _GEN_6919; // @[decode.scala 482:28 540:39]
  wire [63:0] _GEN_6941 = 12'h42 == csrAddrReg ? pmpaddr0 : _GEN_6920; // @[decode.scala 483:28 540:39]
  wire [63:0] _GEN_6942 = 12'h42 == csrAddrReg ? mvendorid : _GEN_6921; // @[decode.scala 484:28 540:39]
  wire [63:0] _GEN_6943 = 12'h42 == csrAddrReg ? marchid : _GEN_6922; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6944 = 12'h42 == csrAddrReg ? mimpid : _GEN_6923; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6945 = 12'h42 == csrAddrReg ? mhartid : _GEN_6924; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6946 = 12'h41 == csrAddrReg ? csrWriteData : uepc; // @[decode.scala 466:28 540:39 543:37]
  wire [63:0] _GEN_6947 = 12'h41 == csrAddrReg ? ucause : _GEN_6925; // @[decode.scala 467:28 540:39]
  wire [63:0] _GEN_6948 = 12'h41 == csrAddrReg ? scounteren : _GEN_6926; // @[decode.scala 468:28 540:39]
  wire [63:0] _GEN_6949 = 12'h41 == csrAddrReg ? satp : _GEN_6927; // @[decode.scala 469:28 540:39]
  wire [63:0] _GEN_6950 = 12'h41 == csrAddrReg ? _mstatus_T_1 : _GEN_6928; // @[decode.scala 489:11 540:39]
  wire [126:0] _GEN_6951 = 12'h41 == csrAddrReg ? 127'h8000000000101101 : _GEN_6929; // @[decode.scala 540:39 490:8]
  wire [63:0] _GEN_6952 = 12'h41 == csrAddrReg ? medeleg : _GEN_6930; // @[decode.scala 472:28 540:39]
  wire [63:0] _GEN_6953 = 12'h41 == csrAddrReg ? mideleg : _GEN_6931; // @[decode.scala 473:28 540:39]
  wire [63:0] _GEN_6954 = 12'h41 == csrAddrReg ? mie : _GEN_6932; // @[decode.scala 474:28 540:39]
  wire [63:0] _GEN_6955 = 12'h41 == csrAddrReg ? mtvec : _GEN_6933; // @[decode.scala 475:28 540:39]
  wire [63:0] _GEN_6956 = 12'h41 == csrAddrReg ? mcounteren : _GEN_6934; // @[decode.scala 476:28 540:39]
  wire [63:0] _GEN_6957 = 12'h41 == csrAddrReg ? mscratch : _GEN_6935; // @[decode.scala 477:28 540:39]
  wire [63:0] _GEN_6958 = 12'h41 == csrAddrReg ? mepc : _GEN_6936; // @[decode.scala 478:28 540:39]
  wire [63:0] _GEN_6959 = 12'h41 == csrAddrReg ? mcause : _GEN_6937; // @[decode.scala 479:28 540:39]
  wire [63:0] _GEN_6960 = 12'h41 == csrAddrReg ? mtval : _GEN_6938; // @[decode.scala 480:28 540:39]
  wire [63:0] _GEN_6961 = 12'h41 == csrAddrReg ? mip : _GEN_6939; // @[decode.scala 481:28 540:39]
  wire [63:0] _GEN_6962 = 12'h41 == csrAddrReg ? pmpcfg0 : _GEN_6940; // @[decode.scala 482:28 540:39]
  wire [63:0] _GEN_6963 = 12'h41 == csrAddrReg ? pmpaddr0 : _GEN_6941; // @[decode.scala 483:28 540:39]
  wire [63:0] _GEN_6964 = 12'h41 == csrAddrReg ? mvendorid : _GEN_6942; // @[decode.scala 484:28 540:39]
  wire [63:0] _GEN_6965 = 12'h41 == csrAddrReg ? marchid : _GEN_6943; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6966 = 12'h41 == csrAddrReg ? mimpid : _GEN_6944; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6967 = 12'h41 == csrAddrReg ? mhartid : _GEN_6945; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6968 = 12'h5 == csrAddrReg ? csrWriteData : utvec; // @[decode.scala 465:28 540:39 542:37]
  wire [63:0] _GEN_6969 = 12'h5 == csrAddrReg ? uepc : _GEN_6946; // @[decode.scala 466:28 540:39]
  wire [63:0] _GEN_6970 = 12'h5 == csrAddrReg ? ucause : _GEN_6947; // @[decode.scala 467:28 540:39]
  wire [63:0] _GEN_6971 = 12'h5 == csrAddrReg ? scounteren : _GEN_6948; // @[decode.scala 468:28 540:39]
  wire [63:0] _GEN_6972 = 12'h5 == csrAddrReg ? satp : _GEN_6949; // @[decode.scala 469:28 540:39]
  wire [63:0] _GEN_6973 = 12'h5 == csrAddrReg ? _mstatus_T_1 : _GEN_6950; // @[decode.scala 489:11 540:39]
  wire [126:0] _GEN_6974 = 12'h5 == csrAddrReg ? 127'h8000000000101101 : _GEN_6951; // @[decode.scala 540:39 490:8]
  wire [63:0] _GEN_6975 = 12'h5 == csrAddrReg ? medeleg : _GEN_6952; // @[decode.scala 472:28 540:39]
  wire [63:0] _GEN_6976 = 12'h5 == csrAddrReg ? mideleg : _GEN_6953; // @[decode.scala 473:28 540:39]
  wire [63:0] _GEN_6977 = 12'h5 == csrAddrReg ? mie : _GEN_6954; // @[decode.scala 474:28 540:39]
  wire [63:0] _GEN_6978 = 12'h5 == csrAddrReg ? mtvec : _GEN_6955; // @[decode.scala 475:28 540:39]
  wire [63:0] _GEN_6979 = 12'h5 == csrAddrReg ? mcounteren : _GEN_6956; // @[decode.scala 476:28 540:39]
  wire [63:0] _GEN_6980 = 12'h5 == csrAddrReg ? mscratch : _GEN_6957; // @[decode.scala 477:28 540:39]
  wire [63:0] _GEN_6981 = 12'h5 == csrAddrReg ? mepc : _GEN_6958; // @[decode.scala 478:28 540:39]
  wire [63:0] _GEN_6982 = 12'h5 == csrAddrReg ? mcause : _GEN_6959; // @[decode.scala 479:28 540:39]
  wire [63:0] _GEN_6983 = 12'h5 == csrAddrReg ? mtval : _GEN_6960; // @[decode.scala 480:28 540:39]
  wire [63:0] _GEN_6984 = 12'h5 == csrAddrReg ? mip : _GEN_6961; // @[decode.scala 481:28 540:39]
  wire [63:0] _GEN_6985 = 12'h5 == csrAddrReg ? pmpcfg0 : _GEN_6962; // @[decode.scala 482:28 540:39]
  wire [63:0] _GEN_6986 = 12'h5 == csrAddrReg ? pmpaddr0 : _GEN_6963; // @[decode.scala 483:28 540:39]
  wire [63:0] _GEN_6987 = 12'h5 == csrAddrReg ? mvendorid : _GEN_6964; // @[decode.scala 484:28 540:39]
  wire [63:0] _GEN_6988 = 12'h5 == csrAddrReg ? marchid : _GEN_6965; // @[decode.scala 485:28 540:39]
  wire [63:0] _GEN_6989 = 12'h5 == csrAddrReg ? mimpid : _GEN_6966; // @[decode.scala 486:28 540:39]
  wire [63:0] _GEN_6990 = 12'h5 == csrAddrReg ? mhartid : _GEN_6967; // @[decode.scala 487:28 540:39]
  wire [63:0] _GEN_6997 = 12'h0 == csrAddrReg ? _mstatus_T_1 : _GEN_6973; // @[decode.scala 489:11 540:39]
  wire [126:0] _GEN_6998 = 12'h0 == csrAddrReg ? 127'h8000000000101101 : _GEN_6974; // @[decode.scala 540:39 490:8]
  wire [63:0] _GEN_7005 = 12'h0 == csrAddrReg ? mepc : _GEN_6981; // @[decode.scala 478:28 540:39]
  wire [63:0] _GEN_7006 = 12'h0 == csrAddrReg ? mcause : _GEN_6982; // @[decode.scala 479:28 540:39]
  wire [63:0] _ustatus_T = ustatus | csrWriteData; // @[decode.scala 569:49]
  wire [63:0] _utvec_T = utvec | csrWriteData; // @[decode.scala 570:47]
  wire [63:0] _uepc_T = uepc | csrWriteData; // @[decode.scala 571:46]
  wire [63:0] _ucause_T = ucause | csrWriteData; // @[decode.scala 572:48]
  wire [63:0] _scounteren_T = scounteren | csrWriteData; // @[decode.scala 573:52]
  wire [63:0] _satp_T = satp | csrWriteData; // @[decode.scala 574:46]
  wire [63:0] _mstatus_T_2 = mstatus | csrWriteData; // @[decode.scala 575:49]
  wire [63:0] _misa_T_2 = misa | csrWriteData; // @[decode.scala 576:46]
  wire [63:0] _medeleg_T = medeleg | csrWriteData; // @[decode.scala 577:49]
  wire [63:0] _mideleg_T = mideleg | csrWriteData; // @[decode.scala 578:49]
  wire [63:0] _mie_T = mie | csrWriteData; // @[decode.scala 579:46]
  wire [63:0] _mtvec_T = mtvec | csrWriteData; // @[decode.scala 580:47]
  wire [63:0] _mcounteren_T = mcounteren | csrWriteData; // @[decode.scala 581:52]
  wire [63:0] _mscratch_T = mscratch | csrWriteData; // @[decode.scala 582:50]
  wire [63:0] _mepc_T = mepc | csrWriteData; // @[decode.scala 583:46]
  wire [63:0] _mcause_T = mcause | csrWriteData; // @[decode.scala 584:48]
  wire [63:0] _mtval_T = mtval | csrWriteData; // @[decode.scala 585:47]
  wire [63:0] _mip_T = mip | csrWriteData; // @[decode.scala 586:45]
  wire [63:0] _pmpcfg0_T = pmpcfg0 | csrWriteData; // @[decode.scala 587:49]
  wire [63:0] _pmpaddr0_T = pmpaddr0 | csrWriteData; // @[decode.scala 588:50]
  wire [63:0] _mvendorid_T = mvendorid | csrWriteData; // @[decode.scala 589:51]
  wire [63:0] _marchid_T = marchid | csrWriteData; // @[decode.scala 590:49]
  wire [63:0] _mimpid_T = mimpid | csrWriteData; // @[decode.scala 591:48]
  wire [63:0] _mhartid_T = mhartid | csrWriteData; // @[decode.scala 592:49]
  wire [63:0] _GEN_7015 = _T_279 ? _mhartid_T : mhartid; // @[decode.scala 487:28 568:39 592:38]
  wire [63:0] _GEN_7016 = _T_278 ? _mimpid_T : mimpid; // @[decode.scala 486:28 568:39 591:38]
  wire [63:0] _GEN_7017 = _T_278 ? mhartid : _GEN_7015; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7018 = _T_277 ? _marchid_T : marchid; // @[decode.scala 485:28 568:39 590:38]
  wire [63:0] _GEN_7019 = _T_277 ? mimpid : _GEN_7016; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7020 = _T_277 ? mhartid : _GEN_7017; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7021 = _T_276 ? _mvendorid_T : mvendorid; // @[decode.scala 484:28 568:39 589:38]
  wire [63:0] _GEN_7022 = _T_276 ? marchid : _GEN_7018; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7023 = _T_276 ? mimpid : _GEN_7019; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7024 = _T_276 ? mhartid : _GEN_7020; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7025 = _T_275 ? _pmpaddr0_T : pmpaddr0; // @[decode.scala 483:28 568:39 588:38]
  wire [63:0] _GEN_7026 = _T_275 ? mvendorid : _GEN_7021; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7027 = _T_275 ? marchid : _GEN_7022; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7028 = _T_275 ? mimpid : _GEN_7023; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7029 = _T_275 ? mhartid : _GEN_7024; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7030 = _T_274 ? _pmpcfg0_T : pmpcfg0; // @[decode.scala 482:28 568:39 587:38]
  wire [63:0] _GEN_7031 = _T_274 ? pmpaddr0 : _GEN_7025; // @[decode.scala 483:28 568:39]
  wire [63:0] _GEN_7032 = _T_274 ? mvendorid : _GEN_7026; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7033 = _T_274 ? marchid : _GEN_7027; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7034 = _T_274 ? mimpid : _GEN_7028; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7035 = _T_274 ? mhartid : _GEN_7029; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7036 = _T_273 ? _mip_T : mip; // @[decode.scala 481:28 568:39 586:38]
  wire [63:0] _GEN_7037 = _T_273 ? pmpcfg0 : _GEN_7030; // @[decode.scala 482:28 568:39]
  wire [63:0] _GEN_7038 = _T_273 ? pmpaddr0 : _GEN_7031; // @[decode.scala 483:28 568:39]
  wire [63:0] _GEN_7039 = _T_273 ? mvendorid : _GEN_7032; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7040 = _T_273 ? marchid : _GEN_7033; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7041 = _T_273 ? mimpid : _GEN_7034; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7042 = _T_273 ? mhartid : _GEN_7035; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7043 = _T_272 ? _mtval_T : mtval; // @[decode.scala 480:28 568:39 585:38]
  wire [63:0] _GEN_7044 = _T_272 ? mip : _GEN_7036; // @[decode.scala 481:28 568:39]
  wire [63:0] _GEN_7045 = _T_272 ? pmpcfg0 : _GEN_7037; // @[decode.scala 482:28 568:39]
  wire [63:0] _GEN_7046 = _T_272 ? pmpaddr0 : _GEN_7038; // @[decode.scala 483:28 568:39]
  wire [63:0] _GEN_7047 = _T_272 ? mvendorid : _GEN_7039; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7048 = _T_272 ? marchid : _GEN_7040; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7049 = _T_272 ? mimpid : _GEN_7041; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7050 = _T_272 ? mhartid : _GEN_7042; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7051 = _T_271 ? _mcause_T : mcause; // @[decode.scala 479:28 568:39 584:38]
  wire [63:0] _GEN_7052 = _T_271 ? mtval : _GEN_7043; // @[decode.scala 480:28 568:39]
  wire [63:0] _GEN_7053 = _T_271 ? mip : _GEN_7044; // @[decode.scala 481:28 568:39]
  wire [63:0] _GEN_7054 = _T_271 ? pmpcfg0 : _GEN_7045; // @[decode.scala 482:28 568:39]
  wire [63:0] _GEN_7055 = _T_271 ? pmpaddr0 : _GEN_7046; // @[decode.scala 483:28 568:39]
  wire [63:0] _GEN_7056 = _T_271 ? mvendorid : _GEN_7047; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7057 = _T_271 ? marchid : _GEN_7048; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7058 = _T_271 ? mimpid : _GEN_7049; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7059 = _T_271 ? mhartid : _GEN_7050; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7060 = _T_270 ? _mepc_T : mepc; // @[decode.scala 478:28 568:39 583:38]
  wire [63:0] _GEN_7061 = _T_270 ? mcause : _GEN_7051; // @[decode.scala 479:28 568:39]
  wire [63:0] _GEN_7062 = _T_270 ? mtval : _GEN_7052; // @[decode.scala 480:28 568:39]
  wire [63:0] _GEN_7063 = _T_270 ? mip : _GEN_7053; // @[decode.scala 481:28 568:39]
  wire [63:0] _GEN_7064 = _T_270 ? pmpcfg0 : _GEN_7054; // @[decode.scala 482:28 568:39]
  wire [63:0] _GEN_7065 = _T_270 ? pmpaddr0 : _GEN_7055; // @[decode.scala 483:28 568:39]
  wire [63:0] _GEN_7066 = _T_270 ? mvendorid : _GEN_7056; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7067 = _T_270 ? marchid : _GEN_7057; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7068 = _T_270 ? mimpid : _GEN_7058; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7069 = _T_270 ? mhartid : _GEN_7059; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7070 = _T_269 ? _mscratch_T : mscratch; // @[decode.scala 477:28 568:39 582:38]
  wire [63:0] _GEN_7071 = _T_269 ? mepc : _GEN_7060; // @[decode.scala 478:28 568:39]
  wire [63:0] _GEN_7072 = _T_269 ? mcause : _GEN_7061; // @[decode.scala 479:28 568:39]
  wire [63:0] _GEN_7073 = _T_269 ? mtval : _GEN_7062; // @[decode.scala 480:28 568:39]
  wire [63:0] _GEN_7074 = _T_269 ? mip : _GEN_7063; // @[decode.scala 481:28 568:39]
  wire [63:0] _GEN_7075 = _T_269 ? pmpcfg0 : _GEN_7064; // @[decode.scala 482:28 568:39]
  wire [63:0] _GEN_7076 = _T_269 ? pmpaddr0 : _GEN_7065; // @[decode.scala 483:28 568:39]
  wire [63:0] _GEN_7077 = _T_269 ? mvendorid : _GEN_7066; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7078 = _T_269 ? marchid : _GEN_7067; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7079 = _T_269 ? mimpid : _GEN_7068; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7080 = _T_269 ? mhartid : _GEN_7069; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7081 = _T_268 ? _mcounteren_T : mcounteren; // @[decode.scala 476:28 568:39 581:38]
  wire [63:0] _GEN_7082 = _T_268 ? mscratch : _GEN_7070; // @[decode.scala 477:28 568:39]
  wire [63:0] _GEN_7083 = _T_268 ? mepc : _GEN_7071; // @[decode.scala 478:28 568:39]
  wire [63:0] _GEN_7084 = _T_268 ? mcause : _GEN_7072; // @[decode.scala 479:28 568:39]
  wire [63:0] _GEN_7085 = _T_268 ? mtval : _GEN_7073; // @[decode.scala 480:28 568:39]
  wire [63:0] _GEN_7086 = _T_268 ? mip : _GEN_7074; // @[decode.scala 481:28 568:39]
  wire [63:0] _GEN_7087 = _T_268 ? pmpcfg0 : _GEN_7075; // @[decode.scala 482:28 568:39]
  wire [63:0] _GEN_7088 = _T_268 ? pmpaddr0 : _GEN_7076; // @[decode.scala 483:28 568:39]
  wire [63:0] _GEN_7089 = _T_268 ? mvendorid : _GEN_7077; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7090 = _T_268 ? marchid : _GEN_7078; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7091 = _T_268 ? mimpid : _GEN_7079; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7092 = _T_268 ? mhartid : _GEN_7080; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7093 = _T_267 ? _mtvec_T : mtvec; // @[decode.scala 475:28 568:39 580:38]
  wire [63:0] _GEN_7094 = _T_267 ? mcounteren : _GEN_7081; // @[decode.scala 476:28 568:39]
  wire [63:0] _GEN_7095 = _T_267 ? mscratch : _GEN_7082; // @[decode.scala 477:28 568:39]
  wire [63:0] _GEN_7096 = _T_267 ? mepc : _GEN_7083; // @[decode.scala 478:28 568:39]
  wire [63:0] _GEN_7097 = _T_267 ? mcause : _GEN_7084; // @[decode.scala 479:28 568:39]
  wire [63:0] _GEN_7098 = _T_267 ? mtval : _GEN_7085; // @[decode.scala 480:28 568:39]
  wire [63:0] _GEN_7099 = _T_267 ? mip : _GEN_7086; // @[decode.scala 481:28 568:39]
  wire [63:0] _GEN_7100 = _T_267 ? pmpcfg0 : _GEN_7087; // @[decode.scala 482:28 568:39]
  wire [63:0] _GEN_7101 = _T_267 ? pmpaddr0 : _GEN_7088; // @[decode.scala 483:28 568:39]
  wire [63:0] _GEN_7102 = _T_267 ? mvendorid : _GEN_7089; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7103 = _T_267 ? marchid : _GEN_7090; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7104 = _T_267 ? mimpid : _GEN_7091; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7105 = _T_267 ? mhartid : _GEN_7092; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7106 = _T_266 ? _mie_T : mie; // @[decode.scala 474:28 568:39 579:38]
  wire [63:0] _GEN_7107 = _T_266 ? mtvec : _GEN_7093; // @[decode.scala 475:28 568:39]
  wire [63:0] _GEN_7108 = _T_266 ? mcounteren : _GEN_7094; // @[decode.scala 476:28 568:39]
  wire [63:0] _GEN_7109 = _T_266 ? mscratch : _GEN_7095; // @[decode.scala 477:28 568:39]
  wire [63:0] _GEN_7110 = _T_266 ? mepc : _GEN_7096; // @[decode.scala 478:28 568:39]
  wire [63:0] _GEN_7111 = _T_266 ? mcause : _GEN_7097; // @[decode.scala 479:28 568:39]
  wire [63:0] _GEN_7112 = _T_266 ? mtval : _GEN_7098; // @[decode.scala 480:28 568:39]
  wire [63:0] _GEN_7113 = _T_266 ? mip : _GEN_7099; // @[decode.scala 481:28 568:39]
  wire [63:0] _GEN_7114 = _T_266 ? pmpcfg0 : _GEN_7100; // @[decode.scala 482:28 568:39]
  wire [63:0] _GEN_7115 = _T_266 ? pmpaddr0 : _GEN_7101; // @[decode.scala 483:28 568:39]
  wire [63:0] _GEN_7116 = _T_266 ? mvendorid : _GEN_7102; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7117 = _T_266 ? marchid : _GEN_7103; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7118 = _T_266 ? mimpid : _GEN_7104; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7119 = _T_266 ? mhartid : _GEN_7105; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7120 = _T_265 ? _mideleg_T : mideleg; // @[decode.scala 473:28 568:39 578:38]
  wire [63:0] _GEN_7121 = _T_265 ? mie : _GEN_7106; // @[decode.scala 474:28 568:39]
  wire [63:0] _GEN_7122 = _T_265 ? mtvec : _GEN_7107; // @[decode.scala 475:28 568:39]
  wire [63:0] _GEN_7123 = _T_265 ? mcounteren : _GEN_7108; // @[decode.scala 476:28 568:39]
  wire [63:0] _GEN_7124 = _T_265 ? mscratch : _GEN_7109; // @[decode.scala 477:28 568:39]
  wire [63:0] _GEN_7125 = _T_265 ? mepc : _GEN_7110; // @[decode.scala 478:28 568:39]
  wire [63:0] _GEN_7126 = _T_265 ? mcause : _GEN_7111; // @[decode.scala 479:28 568:39]
  wire [63:0] _GEN_7127 = _T_265 ? mtval : _GEN_7112; // @[decode.scala 480:28 568:39]
  wire [63:0] _GEN_7128 = _T_265 ? mip : _GEN_7113; // @[decode.scala 481:28 568:39]
  wire [63:0] _GEN_7129 = _T_265 ? pmpcfg0 : _GEN_7114; // @[decode.scala 482:28 568:39]
  wire [63:0] _GEN_7130 = _T_265 ? pmpaddr0 : _GEN_7115; // @[decode.scala 483:28 568:39]
  wire [63:0] _GEN_7131 = _T_265 ? mvendorid : _GEN_7116; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7132 = _T_265 ? marchid : _GEN_7117; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7133 = _T_265 ? mimpid : _GEN_7118; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7134 = _T_265 ? mhartid : _GEN_7119; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7135 = _T_264 ? _medeleg_T : medeleg; // @[decode.scala 472:28 568:39 577:38]
  wire [63:0] _GEN_7136 = _T_264 ? mideleg : _GEN_7120; // @[decode.scala 473:28 568:39]
  wire [63:0] _GEN_7137 = _T_264 ? mie : _GEN_7121; // @[decode.scala 474:28 568:39]
  wire [63:0] _GEN_7138 = _T_264 ? mtvec : _GEN_7122; // @[decode.scala 475:28 568:39]
  wire [63:0] _GEN_7139 = _T_264 ? mcounteren : _GEN_7123; // @[decode.scala 476:28 568:39]
  wire [63:0] _GEN_7140 = _T_264 ? mscratch : _GEN_7124; // @[decode.scala 477:28 568:39]
  wire [63:0] _GEN_7141 = _T_264 ? mepc : _GEN_7125; // @[decode.scala 478:28 568:39]
  wire [63:0] _GEN_7142 = _T_264 ? mcause : _GEN_7126; // @[decode.scala 479:28 568:39]
  wire [63:0] _GEN_7143 = _T_264 ? mtval : _GEN_7127; // @[decode.scala 480:28 568:39]
  wire [63:0] _GEN_7144 = _T_264 ? mip : _GEN_7128; // @[decode.scala 481:28 568:39]
  wire [63:0] _GEN_7145 = _T_264 ? pmpcfg0 : _GEN_7129; // @[decode.scala 482:28 568:39]
  wire [63:0] _GEN_7146 = _T_264 ? pmpaddr0 : _GEN_7130; // @[decode.scala 483:28 568:39]
  wire [63:0] _GEN_7147 = _T_264 ? mvendorid : _GEN_7131; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7148 = _T_264 ? marchid : _GEN_7132; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7149 = _T_264 ? mimpid : _GEN_7133; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7150 = _T_264 ? mhartid : _GEN_7134; // @[decode.scala 487:28 568:39]
  wire [126:0] _GEN_7151 = _T_263 ? {{63'd0}, _misa_T_2} : 127'h8000000000101101; // @[decode.scala 568:39 576:38 490:8]
  wire [63:0] _GEN_7152 = _T_263 ? medeleg : _GEN_7135; // @[decode.scala 472:28 568:39]
  wire [63:0] _GEN_7153 = _T_263 ? mideleg : _GEN_7136; // @[decode.scala 473:28 568:39]
  wire [63:0] _GEN_7154 = _T_263 ? mie : _GEN_7137; // @[decode.scala 474:28 568:39]
  wire [63:0] _GEN_7155 = _T_263 ? mtvec : _GEN_7138; // @[decode.scala 475:28 568:39]
  wire [63:0] _GEN_7156 = _T_263 ? mcounteren : _GEN_7139; // @[decode.scala 476:28 568:39]
  wire [63:0] _GEN_7157 = _T_263 ? mscratch : _GEN_7140; // @[decode.scala 477:28 568:39]
  wire [63:0] _GEN_7158 = _T_263 ? mepc : _GEN_7141; // @[decode.scala 478:28 568:39]
  wire [63:0] _GEN_7159 = _T_263 ? mcause : _GEN_7142; // @[decode.scala 479:28 568:39]
  wire [63:0] _GEN_7160 = _T_263 ? mtval : _GEN_7143; // @[decode.scala 480:28 568:39]
  wire [63:0] _GEN_7161 = _T_263 ? mip : _GEN_7144; // @[decode.scala 481:28 568:39]
  wire [63:0] _GEN_7162 = _T_263 ? pmpcfg0 : _GEN_7145; // @[decode.scala 482:28 568:39]
  wire [63:0] _GEN_7163 = _T_263 ? pmpaddr0 : _GEN_7146; // @[decode.scala 483:28 568:39]
  wire [63:0] _GEN_7164 = _T_263 ? mvendorid : _GEN_7147; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7165 = _T_263 ? marchid : _GEN_7148; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7166 = _T_263 ? mimpid : _GEN_7149; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7167 = _T_263 ? mhartid : _GEN_7150; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7168 = _T_262 ? _mstatus_T_2 : _mstatus_T_1; // @[decode.scala 489:11 568:39 575:38]
  wire [126:0] _GEN_7169 = _T_262 ? 127'h8000000000101101 : _GEN_7151; // @[decode.scala 568:39 490:8]
  wire [63:0] _GEN_7170 = _T_262 ? medeleg : _GEN_7152; // @[decode.scala 472:28 568:39]
  wire [63:0] _GEN_7171 = _T_262 ? mideleg : _GEN_7153; // @[decode.scala 473:28 568:39]
  wire [63:0] _GEN_7172 = _T_262 ? mie : _GEN_7154; // @[decode.scala 474:28 568:39]
  wire [63:0] _GEN_7173 = _T_262 ? mtvec : _GEN_7155; // @[decode.scala 475:28 568:39]
  wire [63:0] _GEN_7174 = _T_262 ? mcounteren : _GEN_7156; // @[decode.scala 476:28 568:39]
  wire [63:0] _GEN_7175 = _T_262 ? mscratch : _GEN_7157; // @[decode.scala 477:28 568:39]
  wire [63:0] _GEN_7176 = _T_262 ? mepc : _GEN_7158; // @[decode.scala 478:28 568:39]
  wire [63:0] _GEN_7177 = _T_262 ? mcause : _GEN_7159; // @[decode.scala 479:28 568:39]
  wire [63:0] _GEN_7178 = _T_262 ? mtval : _GEN_7160; // @[decode.scala 480:28 568:39]
  wire [63:0] _GEN_7179 = _T_262 ? mip : _GEN_7161; // @[decode.scala 481:28 568:39]
  wire [63:0] _GEN_7180 = _T_262 ? pmpcfg0 : _GEN_7162; // @[decode.scala 482:28 568:39]
  wire [63:0] _GEN_7181 = _T_262 ? pmpaddr0 : _GEN_7163; // @[decode.scala 483:28 568:39]
  wire [63:0] _GEN_7182 = _T_262 ? mvendorid : _GEN_7164; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7183 = _T_262 ? marchid : _GEN_7165; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7184 = _T_262 ? mimpid : _GEN_7166; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7185 = _T_262 ? mhartid : _GEN_7167; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7186 = _T_261 ? _satp_T : satp; // @[decode.scala 469:28 568:39 574:38]
  wire [63:0] _GEN_7187 = _T_261 ? _mstatus_T_1 : _GEN_7168; // @[decode.scala 489:11 568:39]
  wire [126:0] _GEN_7188 = _T_261 ? 127'h8000000000101101 : _GEN_7169; // @[decode.scala 568:39 490:8]
  wire [63:0] _GEN_7189 = _T_261 ? medeleg : _GEN_7170; // @[decode.scala 472:28 568:39]
  wire [63:0] _GEN_7190 = _T_261 ? mideleg : _GEN_7171; // @[decode.scala 473:28 568:39]
  wire [63:0] _GEN_7191 = _T_261 ? mie : _GEN_7172; // @[decode.scala 474:28 568:39]
  wire [63:0] _GEN_7192 = _T_261 ? mtvec : _GEN_7173; // @[decode.scala 475:28 568:39]
  wire [63:0] _GEN_7193 = _T_261 ? mcounteren : _GEN_7174; // @[decode.scala 476:28 568:39]
  wire [63:0] _GEN_7194 = _T_261 ? mscratch : _GEN_7175; // @[decode.scala 477:28 568:39]
  wire [63:0] _GEN_7195 = _T_261 ? mepc : _GEN_7176; // @[decode.scala 478:28 568:39]
  wire [63:0] _GEN_7196 = _T_261 ? mcause : _GEN_7177; // @[decode.scala 479:28 568:39]
  wire [63:0] _GEN_7197 = _T_261 ? mtval : _GEN_7178; // @[decode.scala 480:28 568:39]
  wire [63:0] _GEN_7198 = _T_261 ? mip : _GEN_7179; // @[decode.scala 481:28 568:39]
  wire [63:0] _GEN_7199 = _T_261 ? pmpcfg0 : _GEN_7180; // @[decode.scala 482:28 568:39]
  wire [63:0] _GEN_7200 = _T_261 ? pmpaddr0 : _GEN_7181; // @[decode.scala 483:28 568:39]
  wire [63:0] _GEN_7201 = _T_261 ? mvendorid : _GEN_7182; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7202 = _T_261 ? marchid : _GEN_7183; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7203 = _T_261 ? mimpid : _GEN_7184; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7204 = _T_261 ? mhartid : _GEN_7185; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7205 = _T_260 ? _scounteren_T : scounteren; // @[decode.scala 468:28 568:39 573:38]
  wire [63:0] _GEN_7206 = _T_260 ? satp : _GEN_7186; // @[decode.scala 469:28 568:39]
  wire [63:0] _GEN_7207 = _T_260 ? _mstatus_T_1 : _GEN_7187; // @[decode.scala 489:11 568:39]
  wire [126:0] _GEN_7208 = _T_260 ? 127'h8000000000101101 : _GEN_7188; // @[decode.scala 568:39 490:8]
  wire [63:0] _GEN_7209 = _T_260 ? medeleg : _GEN_7189; // @[decode.scala 472:28 568:39]
  wire [63:0] _GEN_7210 = _T_260 ? mideleg : _GEN_7190; // @[decode.scala 473:28 568:39]
  wire [63:0] _GEN_7211 = _T_260 ? mie : _GEN_7191; // @[decode.scala 474:28 568:39]
  wire [63:0] _GEN_7212 = _T_260 ? mtvec : _GEN_7192; // @[decode.scala 475:28 568:39]
  wire [63:0] _GEN_7213 = _T_260 ? mcounteren : _GEN_7193; // @[decode.scala 476:28 568:39]
  wire [63:0] _GEN_7214 = _T_260 ? mscratch : _GEN_7194; // @[decode.scala 477:28 568:39]
  wire [63:0] _GEN_7215 = _T_260 ? mepc : _GEN_7195; // @[decode.scala 478:28 568:39]
  wire [63:0] _GEN_7216 = _T_260 ? mcause : _GEN_7196; // @[decode.scala 479:28 568:39]
  wire [63:0] _GEN_7217 = _T_260 ? mtval : _GEN_7197; // @[decode.scala 480:28 568:39]
  wire [63:0] _GEN_7218 = _T_260 ? mip : _GEN_7198; // @[decode.scala 481:28 568:39]
  wire [63:0] _GEN_7219 = _T_260 ? pmpcfg0 : _GEN_7199; // @[decode.scala 482:28 568:39]
  wire [63:0] _GEN_7220 = _T_260 ? pmpaddr0 : _GEN_7200; // @[decode.scala 483:28 568:39]
  wire [63:0] _GEN_7221 = _T_260 ? mvendorid : _GEN_7201; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7222 = _T_260 ? marchid : _GEN_7202; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7223 = _T_260 ? mimpid : _GEN_7203; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7224 = _T_260 ? mhartid : _GEN_7204; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7225 = _T_259 ? _ucause_T : ucause; // @[decode.scala 467:28 568:39 572:38]
  wire [63:0] _GEN_7226 = _T_259 ? scounteren : _GEN_7205; // @[decode.scala 468:28 568:39]
  wire [63:0] _GEN_7227 = _T_259 ? satp : _GEN_7206; // @[decode.scala 469:28 568:39]
  wire [63:0] _GEN_7228 = _T_259 ? _mstatus_T_1 : _GEN_7207; // @[decode.scala 489:11 568:39]
  wire [126:0] _GEN_7229 = _T_259 ? 127'h8000000000101101 : _GEN_7208; // @[decode.scala 568:39 490:8]
  wire [63:0] _GEN_7230 = _T_259 ? medeleg : _GEN_7209; // @[decode.scala 472:28 568:39]
  wire [63:0] _GEN_7231 = _T_259 ? mideleg : _GEN_7210; // @[decode.scala 473:28 568:39]
  wire [63:0] _GEN_7232 = _T_259 ? mie : _GEN_7211; // @[decode.scala 474:28 568:39]
  wire [63:0] _GEN_7233 = _T_259 ? mtvec : _GEN_7212; // @[decode.scala 475:28 568:39]
  wire [63:0] _GEN_7234 = _T_259 ? mcounteren : _GEN_7213; // @[decode.scala 476:28 568:39]
  wire [63:0] _GEN_7235 = _T_259 ? mscratch : _GEN_7214; // @[decode.scala 477:28 568:39]
  wire [63:0] _GEN_7236 = _T_259 ? mepc : _GEN_7215; // @[decode.scala 478:28 568:39]
  wire [63:0] _GEN_7237 = _T_259 ? mcause : _GEN_7216; // @[decode.scala 479:28 568:39]
  wire [63:0] _GEN_7238 = _T_259 ? mtval : _GEN_7217; // @[decode.scala 480:28 568:39]
  wire [63:0] _GEN_7239 = _T_259 ? mip : _GEN_7218; // @[decode.scala 481:28 568:39]
  wire [63:0] _GEN_7240 = _T_259 ? pmpcfg0 : _GEN_7219; // @[decode.scala 482:28 568:39]
  wire [63:0] _GEN_7241 = _T_259 ? pmpaddr0 : _GEN_7220; // @[decode.scala 483:28 568:39]
  wire [63:0] _GEN_7242 = _T_259 ? mvendorid : _GEN_7221; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7243 = _T_259 ? marchid : _GEN_7222; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7244 = _T_259 ? mimpid : _GEN_7223; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7245 = _T_259 ? mhartid : _GEN_7224; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7246 = _T_258 ? _uepc_T : uepc; // @[decode.scala 466:28 568:39 571:38]
  wire [63:0] _GEN_7247 = _T_258 ? ucause : _GEN_7225; // @[decode.scala 467:28 568:39]
  wire [63:0] _GEN_7248 = _T_258 ? scounteren : _GEN_7226; // @[decode.scala 468:28 568:39]
  wire [63:0] _GEN_7249 = _T_258 ? satp : _GEN_7227; // @[decode.scala 469:28 568:39]
  wire [63:0] _GEN_7250 = _T_258 ? _mstatus_T_1 : _GEN_7228; // @[decode.scala 489:11 568:39]
  wire [126:0] _GEN_7251 = _T_258 ? 127'h8000000000101101 : _GEN_7229; // @[decode.scala 568:39 490:8]
  wire [63:0] _GEN_7252 = _T_258 ? medeleg : _GEN_7230; // @[decode.scala 472:28 568:39]
  wire [63:0] _GEN_7253 = _T_258 ? mideleg : _GEN_7231; // @[decode.scala 473:28 568:39]
  wire [63:0] _GEN_7254 = _T_258 ? mie : _GEN_7232; // @[decode.scala 474:28 568:39]
  wire [63:0] _GEN_7255 = _T_258 ? mtvec : _GEN_7233; // @[decode.scala 475:28 568:39]
  wire [63:0] _GEN_7256 = _T_258 ? mcounteren : _GEN_7234; // @[decode.scala 476:28 568:39]
  wire [63:0] _GEN_7257 = _T_258 ? mscratch : _GEN_7235; // @[decode.scala 477:28 568:39]
  wire [63:0] _GEN_7258 = _T_258 ? mepc : _GEN_7236; // @[decode.scala 478:28 568:39]
  wire [63:0] _GEN_7259 = _T_258 ? mcause : _GEN_7237; // @[decode.scala 479:28 568:39]
  wire [63:0] _GEN_7260 = _T_258 ? mtval : _GEN_7238; // @[decode.scala 480:28 568:39]
  wire [63:0] _GEN_7261 = _T_258 ? mip : _GEN_7239; // @[decode.scala 481:28 568:39]
  wire [63:0] _GEN_7262 = _T_258 ? pmpcfg0 : _GEN_7240; // @[decode.scala 482:28 568:39]
  wire [63:0] _GEN_7263 = _T_258 ? pmpaddr0 : _GEN_7241; // @[decode.scala 483:28 568:39]
  wire [63:0] _GEN_7264 = _T_258 ? mvendorid : _GEN_7242; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7265 = _T_258 ? marchid : _GEN_7243; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7266 = _T_258 ? mimpid : _GEN_7244; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7267 = _T_258 ? mhartid : _GEN_7245; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7268 = _T_257 ? _utvec_T : utvec; // @[decode.scala 465:28 568:39 570:38]
  wire [63:0] _GEN_7269 = _T_257 ? uepc : _GEN_7246; // @[decode.scala 466:28 568:39]
  wire [63:0] _GEN_7270 = _T_257 ? ucause : _GEN_7247; // @[decode.scala 467:28 568:39]
  wire [63:0] _GEN_7271 = _T_257 ? scounteren : _GEN_7248; // @[decode.scala 468:28 568:39]
  wire [63:0] _GEN_7272 = _T_257 ? satp : _GEN_7249; // @[decode.scala 469:28 568:39]
  wire [63:0] _GEN_7273 = _T_257 ? _mstatus_T_1 : _GEN_7250; // @[decode.scala 489:11 568:39]
  wire [126:0] _GEN_7274 = _T_257 ? 127'h8000000000101101 : _GEN_7251; // @[decode.scala 568:39 490:8]
  wire [63:0] _GEN_7275 = _T_257 ? medeleg : _GEN_7252; // @[decode.scala 472:28 568:39]
  wire [63:0] _GEN_7276 = _T_257 ? mideleg : _GEN_7253; // @[decode.scala 473:28 568:39]
  wire [63:0] _GEN_7277 = _T_257 ? mie : _GEN_7254; // @[decode.scala 474:28 568:39]
  wire [63:0] _GEN_7278 = _T_257 ? mtvec : _GEN_7255; // @[decode.scala 475:28 568:39]
  wire [63:0] _GEN_7279 = _T_257 ? mcounteren : _GEN_7256; // @[decode.scala 476:28 568:39]
  wire [63:0] _GEN_7280 = _T_257 ? mscratch : _GEN_7257; // @[decode.scala 477:28 568:39]
  wire [63:0] _GEN_7281 = _T_257 ? mepc : _GEN_7258; // @[decode.scala 478:28 568:39]
  wire [63:0] _GEN_7282 = _T_257 ? mcause : _GEN_7259; // @[decode.scala 479:28 568:39]
  wire [63:0] _GEN_7283 = _T_257 ? mtval : _GEN_7260; // @[decode.scala 480:28 568:39]
  wire [63:0] _GEN_7284 = _T_257 ? mip : _GEN_7261; // @[decode.scala 481:28 568:39]
  wire [63:0] _GEN_7285 = _T_257 ? pmpcfg0 : _GEN_7262; // @[decode.scala 482:28 568:39]
  wire [63:0] _GEN_7286 = _T_257 ? pmpaddr0 : _GEN_7263; // @[decode.scala 483:28 568:39]
  wire [63:0] _GEN_7287 = _T_257 ? mvendorid : _GEN_7264; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7288 = _T_257 ? marchid : _GEN_7265; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7289 = _T_257 ? mimpid : _GEN_7266; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7290 = _T_257 ? mhartid : _GEN_7267; // @[decode.scala 487:28 568:39]
  wire [63:0] _GEN_7291 = _T_256 ? _ustatus_T : ustatus; // @[decode.scala 464:28 568:39 569:38]
  wire [63:0] _GEN_7292 = _T_256 ? utvec : _GEN_7268; // @[decode.scala 465:28 568:39]
  wire [63:0] _GEN_7293 = _T_256 ? uepc : _GEN_7269; // @[decode.scala 466:28 568:39]
  wire [63:0] _GEN_7294 = _T_256 ? ucause : _GEN_7270; // @[decode.scala 467:28 568:39]
  wire [63:0] _GEN_7295 = _T_256 ? scounteren : _GEN_7271; // @[decode.scala 468:28 568:39]
  wire [63:0] _GEN_7296 = _T_256 ? satp : _GEN_7272; // @[decode.scala 469:28 568:39]
  wire [63:0] _GEN_7297 = _T_256 ? _mstatus_T_1 : _GEN_7273; // @[decode.scala 489:11 568:39]
  wire [126:0] _GEN_7298 = _T_256 ? 127'h8000000000101101 : _GEN_7274; // @[decode.scala 568:39 490:8]
  wire [63:0] _GEN_7299 = _T_256 ? medeleg : _GEN_7275; // @[decode.scala 472:28 568:39]
  wire [63:0] _GEN_7300 = _T_256 ? mideleg : _GEN_7276; // @[decode.scala 473:28 568:39]
  wire [63:0] _GEN_7301 = _T_256 ? mie : _GEN_7277; // @[decode.scala 474:28 568:39]
  wire [63:0] _GEN_7302 = _T_256 ? mtvec : _GEN_7278; // @[decode.scala 475:28 568:39]
  wire [63:0] _GEN_7303 = _T_256 ? mcounteren : _GEN_7279; // @[decode.scala 476:28 568:39]
  wire [63:0] _GEN_7304 = _T_256 ? mscratch : _GEN_7280; // @[decode.scala 477:28 568:39]
  wire [63:0] _GEN_7305 = _T_256 ? mepc : _GEN_7281; // @[decode.scala 478:28 568:39]
  wire [63:0] _GEN_7306 = _T_256 ? mcause : _GEN_7282; // @[decode.scala 479:28 568:39]
  wire [63:0] _GEN_7307 = _T_256 ? mtval : _GEN_7283; // @[decode.scala 480:28 568:39]
  wire [63:0] _GEN_7308 = _T_256 ? mip : _GEN_7284; // @[decode.scala 481:28 568:39]
  wire [63:0] _GEN_7309 = _T_256 ? pmpcfg0 : _GEN_7285; // @[decode.scala 482:28 568:39]
  wire [63:0] _GEN_7310 = _T_256 ? pmpaddr0 : _GEN_7286; // @[decode.scala 483:28 568:39]
  wire [63:0] _GEN_7311 = _T_256 ? mvendorid : _GEN_7287; // @[decode.scala 484:28 568:39]
  wire [63:0] _GEN_7312 = _T_256 ? marchid : _GEN_7288; // @[decode.scala 485:28 568:39]
  wire [63:0] _GEN_7313 = _T_256 ? mimpid : _GEN_7289; // @[decode.scala 486:28 568:39]
  wire [63:0] _GEN_7314 = _T_256 ? mhartid : _GEN_7290; // @[decode.scala 487:28 568:39]
  wire [63:0] _ustatus_T_1 = ~csrWriteData; // @[decode.scala 597:51]
  wire [63:0] _ustatus_T_2 = ustatus & _ustatus_T_1; // @[decode.scala 597:49]
  wire [63:0] _utvec_T_2 = mtvec & _ustatus_T_1; // @[decode.scala 598:47]
  wire [63:0] _uepc_T_2 = uepc & _ustatus_T_1; // @[decode.scala 599:46]
  wire [63:0] _ucause_T_2 = ucause & _ustatus_T_1; // @[decode.scala 600:48]
  wire [63:0] _scounteren_T_2 = scounteren & _ustatus_T_1; // @[decode.scala 601:52]
  wire [63:0] _satp_T_2 = satp & _ustatus_T_1; // @[decode.scala 602:46]
  wire [63:0] _mstatus_T_4 = mstatus & _ustatus_T_1; // @[decode.scala 603:49]
  wire [63:0] _misa_T_4 = misa & _ustatus_T_1; // @[decode.scala 604:46]
  wire [63:0] _medeleg_T_2 = medeleg & _ustatus_T_1; // @[decode.scala 605:49]
  wire [63:0] _mideleg_T_2 = mideleg & _ustatus_T_1; // @[decode.scala 606:49]
  wire [63:0] _mie_T_2 = mie & _ustatus_T_1; // @[decode.scala 607:45]
  wire [63:0] _mcounteren_T_2 = mcounteren & _ustatus_T_1; // @[decode.scala 609:52]
  wire [63:0] _mscratch_T_2 = mscratch & _ustatus_T_1; // @[decode.scala 610:50]
  wire [63:0] _mepc_T_2 = mepc & _ustatus_T_1; // @[decode.scala 611:46]
  wire [63:0] _mcause_T_2 = mcause & _ustatus_T_1; // @[decode.scala 612:48]
  wire [63:0] _mtval_T_2 = mtval & _ustatus_T_1; // @[decode.scala 613:47]
  wire [63:0] _mip_T_2 = mip & _ustatus_T_1; // @[decode.scala 614:45]
  wire [63:0] _pmpcfg0_T_2 = pmpcfg0 & _ustatus_T_1; // @[decode.scala 615:49]
  wire [63:0] _pmpaddr0_T_2 = pmpaddr0 & _ustatus_T_1; // @[decode.scala 616:50]
  wire [63:0] _mvendorid_T_2 = mvendorid & _ustatus_T_1; // @[decode.scala 617:51]
  wire [63:0] _marchid_T_2 = marchid & _ustatus_T_1; // @[decode.scala 618:49]
  wire [63:0] _mimpid_T_2 = mimpid & _ustatus_T_1; // @[decode.scala 619:48]
  wire [63:0] _mhartid_T_2 = mhartid & _ustatus_T_1; // @[decode.scala 620:49]
  wire [63:0] _GEN_7315 = _T_279 ? _mhartid_T_2 : mhartid; // @[decode.scala 487:28 596:39 620:38]
  wire [63:0] _GEN_7316 = _T_278 ? _mimpid_T_2 : mimpid; // @[decode.scala 486:28 596:39 619:38]
  wire [63:0] _GEN_7317 = _T_278 ? mhartid : _GEN_7315; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7318 = _T_277 ? _marchid_T_2 : marchid; // @[decode.scala 485:28 596:39 618:38]
  wire [63:0] _GEN_7319 = _T_277 ? mimpid : _GEN_7316; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7320 = _T_277 ? mhartid : _GEN_7317; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7321 = _T_276 ? _mvendorid_T_2 : mvendorid; // @[decode.scala 484:28 596:39 617:38]
  wire [63:0] _GEN_7322 = _T_276 ? marchid : _GEN_7318; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7323 = _T_276 ? mimpid : _GEN_7319; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7324 = _T_276 ? mhartid : _GEN_7320; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7325 = _T_275 ? _pmpaddr0_T_2 : pmpaddr0; // @[decode.scala 483:28 596:39 616:38]
  wire [63:0] _GEN_7326 = _T_275 ? mvendorid : _GEN_7321; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7327 = _T_275 ? marchid : _GEN_7322; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7328 = _T_275 ? mimpid : _GEN_7323; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7329 = _T_275 ? mhartid : _GEN_7324; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7330 = _T_274 ? _pmpcfg0_T_2 : pmpcfg0; // @[decode.scala 482:28 596:39 615:38]
  wire [63:0] _GEN_7331 = _T_274 ? pmpaddr0 : _GEN_7325; // @[decode.scala 483:28 596:39]
  wire [63:0] _GEN_7332 = _T_274 ? mvendorid : _GEN_7326; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7333 = _T_274 ? marchid : _GEN_7327; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7334 = _T_274 ? mimpid : _GEN_7328; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7335 = _T_274 ? mhartid : _GEN_7329; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7336 = _T_273 ? _mip_T_2 : mip; // @[decode.scala 481:28 596:39 614:38]
  wire [63:0] _GEN_7337 = _T_273 ? pmpcfg0 : _GEN_7330; // @[decode.scala 482:28 596:39]
  wire [63:0] _GEN_7338 = _T_273 ? pmpaddr0 : _GEN_7331; // @[decode.scala 483:28 596:39]
  wire [63:0] _GEN_7339 = _T_273 ? mvendorid : _GEN_7332; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7340 = _T_273 ? marchid : _GEN_7333; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7341 = _T_273 ? mimpid : _GEN_7334; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7342 = _T_273 ? mhartid : _GEN_7335; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7343 = _T_272 ? _mtval_T_2 : mtval; // @[decode.scala 480:28 596:39 613:38]
  wire [63:0] _GEN_7344 = _T_272 ? mip : _GEN_7336; // @[decode.scala 481:28 596:39]
  wire [63:0] _GEN_7345 = _T_272 ? pmpcfg0 : _GEN_7337; // @[decode.scala 482:28 596:39]
  wire [63:0] _GEN_7346 = _T_272 ? pmpaddr0 : _GEN_7338; // @[decode.scala 483:28 596:39]
  wire [63:0] _GEN_7347 = _T_272 ? mvendorid : _GEN_7339; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7348 = _T_272 ? marchid : _GEN_7340; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7349 = _T_272 ? mimpid : _GEN_7341; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7350 = _T_272 ? mhartid : _GEN_7342; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7351 = _T_271 ? _mcause_T_2 : mcause; // @[decode.scala 479:28 596:39 612:38]
  wire [63:0] _GEN_7352 = _T_271 ? mtval : _GEN_7343; // @[decode.scala 480:28 596:39]
  wire [63:0] _GEN_7353 = _T_271 ? mip : _GEN_7344; // @[decode.scala 481:28 596:39]
  wire [63:0] _GEN_7354 = _T_271 ? pmpcfg0 : _GEN_7345; // @[decode.scala 482:28 596:39]
  wire [63:0] _GEN_7355 = _T_271 ? pmpaddr0 : _GEN_7346; // @[decode.scala 483:28 596:39]
  wire [63:0] _GEN_7356 = _T_271 ? mvendorid : _GEN_7347; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7357 = _T_271 ? marchid : _GEN_7348; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7358 = _T_271 ? mimpid : _GEN_7349; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7359 = _T_271 ? mhartid : _GEN_7350; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7360 = _T_270 ? _mepc_T_2 : mepc; // @[decode.scala 478:28 596:39 611:38]
  wire [63:0] _GEN_7361 = _T_270 ? mcause : _GEN_7351; // @[decode.scala 479:28 596:39]
  wire [63:0] _GEN_7362 = _T_270 ? mtval : _GEN_7352; // @[decode.scala 480:28 596:39]
  wire [63:0] _GEN_7363 = _T_270 ? mip : _GEN_7353; // @[decode.scala 481:28 596:39]
  wire [63:0] _GEN_7364 = _T_270 ? pmpcfg0 : _GEN_7354; // @[decode.scala 482:28 596:39]
  wire [63:0] _GEN_7365 = _T_270 ? pmpaddr0 : _GEN_7355; // @[decode.scala 483:28 596:39]
  wire [63:0] _GEN_7366 = _T_270 ? mvendorid : _GEN_7356; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7367 = _T_270 ? marchid : _GEN_7357; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7368 = _T_270 ? mimpid : _GEN_7358; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7369 = _T_270 ? mhartid : _GEN_7359; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7370 = _T_269 ? _mscratch_T_2 : mscratch; // @[decode.scala 477:28 596:39 610:38]
  wire [63:0] _GEN_7371 = _T_269 ? mepc : _GEN_7360; // @[decode.scala 478:28 596:39]
  wire [63:0] _GEN_7372 = _T_269 ? mcause : _GEN_7361; // @[decode.scala 479:28 596:39]
  wire [63:0] _GEN_7373 = _T_269 ? mtval : _GEN_7362; // @[decode.scala 480:28 596:39]
  wire [63:0] _GEN_7374 = _T_269 ? mip : _GEN_7363; // @[decode.scala 481:28 596:39]
  wire [63:0] _GEN_7375 = _T_269 ? pmpcfg0 : _GEN_7364; // @[decode.scala 482:28 596:39]
  wire [63:0] _GEN_7376 = _T_269 ? pmpaddr0 : _GEN_7365; // @[decode.scala 483:28 596:39]
  wire [63:0] _GEN_7377 = _T_269 ? mvendorid : _GEN_7366; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7378 = _T_269 ? marchid : _GEN_7367; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7379 = _T_269 ? mimpid : _GEN_7368; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7380 = _T_269 ? mhartid : _GEN_7369; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7381 = _T_268 ? _mcounteren_T_2 : mcounteren; // @[decode.scala 476:28 596:39 609:38]
  wire [63:0] _GEN_7382 = _T_268 ? mscratch : _GEN_7370; // @[decode.scala 477:28 596:39]
  wire [63:0] _GEN_7383 = _T_268 ? mepc : _GEN_7371; // @[decode.scala 478:28 596:39]
  wire [63:0] _GEN_7384 = _T_268 ? mcause : _GEN_7372; // @[decode.scala 479:28 596:39]
  wire [63:0] _GEN_7385 = _T_268 ? mtval : _GEN_7373; // @[decode.scala 480:28 596:39]
  wire [63:0] _GEN_7386 = _T_268 ? mip : _GEN_7374; // @[decode.scala 481:28 596:39]
  wire [63:0] _GEN_7387 = _T_268 ? pmpcfg0 : _GEN_7375; // @[decode.scala 482:28 596:39]
  wire [63:0] _GEN_7388 = _T_268 ? pmpaddr0 : _GEN_7376; // @[decode.scala 483:28 596:39]
  wire [63:0] _GEN_7389 = _T_268 ? mvendorid : _GEN_7377; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7390 = _T_268 ? marchid : _GEN_7378; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7391 = _T_268 ? mimpid : _GEN_7379; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7392 = _T_268 ? mhartid : _GEN_7380; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7393 = _T_267 ? _utvec_T_2 : mtvec; // @[decode.scala 475:28 596:39 608:38]
  wire [63:0] _GEN_7394 = _T_267 ? mcounteren : _GEN_7381; // @[decode.scala 476:28 596:39]
  wire [63:0] _GEN_7395 = _T_267 ? mscratch : _GEN_7382; // @[decode.scala 477:28 596:39]
  wire [63:0] _GEN_7396 = _T_267 ? mepc : _GEN_7383; // @[decode.scala 478:28 596:39]
  wire [63:0] _GEN_7397 = _T_267 ? mcause : _GEN_7384; // @[decode.scala 479:28 596:39]
  wire [63:0] _GEN_7398 = _T_267 ? mtval : _GEN_7385; // @[decode.scala 480:28 596:39]
  wire [63:0] _GEN_7399 = _T_267 ? mip : _GEN_7386; // @[decode.scala 481:28 596:39]
  wire [63:0] _GEN_7400 = _T_267 ? pmpcfg0 : _GEN_7387; // @[decode.scala 482:28 596:39]
  wire [63:0] _GEN_7401 = _T_267 ? pmpaddr0 : _GEN_7388; // @[decode.scala 483:28 596:39]
  wire [63:0] _GEN_7402 = _T_267 ? mvendorid : _GEN_7389; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7403 = _T_267 ? marchid : _GEN_7390; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7404 = _T_267 ? mimpid : _GEN_7391; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7405 = _T_267 ? mhartid : _GEN_7392; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7406 = _T_266 ? _mie_T_2 : mie; // @[decode.scala 474:28 596:39 607:38]
  wire [63:0] _GEN_7407 = _T_266 ? mtvec : _GEN_7393; // @[decode.scala 475:28 596:39]
  wire [63:0] _GEN_7408 = _T_266 ? mcounteren : _GEN_7394; // @[decode.scala 476:28 596:39]
  wire [63:0] _GEN_7409 = _T_266 ? mscratch : _GEN_7395; // @[decode.scala 477:28 596:39]
  wire [63:0] _GEN_7410 = _T_266 ? mepc : _GEN_7396; // @[decode.scala 478:28 596:39]
  wire [63:0] _GEN_7411 = _T_266 ? mcause : _GEN_7397; // @[decode.scala 479:28 596:39]
  wire [63:0] _GEN_7412 = _T_266 ? mtval : _GEN_7398; // @[decode.scala 480:28 596:39]
  wire [63:0] _GEN_7413 = _T_266 ? mip : _GEN_7399; // @[decode.scala 481:28 596:39]
  wire [63:0] _GEN_7414 = _T_266 ? pmpcfg0 : _GEN_7400; // @[decode.scala 482:28 596:39]
  wire [63:0] _GEN_7415 = _T_266 ? pmpaddr0 : _GEN_7401; // @[decode.scala 483:28 596:39]
  wire [63:0] _GEN_7416 = _T_266 ? mvendorid : _GEN_7402; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7417 = _T_266 ? marchid : _GEN_7403; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7418 = _T_266 ? mimpid : _GEN_7404; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7419 = _T_266 ? mhartid : _GEN_7405; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7420 = _T_265 ? _mideleg_T_2 : mideleg; // @[decode.scala 473:28 596:39 606:38]
  wire [63:0] _GEN_7421 = _T_265 ? mie : _GEN_7406; // @[decode.scala 474:28 596:39]
  wire [63:0] _GEN_7422 = _T_265 ? mtvec : _GEN_7407; // @[decode.scala 475:28 596:39]
  wire [63:0] _GEN_7423 = _T_265 ? mcounteren : _GEN_7408; // @[decode.scala 476:28 596:39]
  wire [63:0] _GEN_7424 = _T_265 ? mscratch : _GEN_7409; // @[decode.scala 477:28 596:39]
  wire [63:0] _GEN_7425 = _T_265 ? mepc : _GEN_7410; // @[decode.scala 478:28 596:39]
  wire [63:0] _GEN_7426 = _T_265 ? mcause : _GEN_7411; // @[decode.scala 479:28 596:39]
  wire [63:0] _GEN_7427 = _T_265 ? mtval : _GEN_7412; // @[decode.scala 480:28 596:39]
  wire [63:0] _GEN_7428 = _T_265 ? mip : _GEN_7413; // @[decode.scala 481:28 596:39]
  wire [63:0] _GEN_7429 = _T_265 ? pmpcfg0 : _GEN_7414; // @[decode.scala 482:28 596:39]
  wire [63:0] _GEN_7430 = _T_265 ? pmpaddr0 : _GEN_7415; // @[decode.scala 483:28 596:39]
  wire [63:0] _GEN_7431 = _T_265 ? mvendorid : _GEN_7416; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7432 = _T_265 ? marchid : _GEN_7417; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7433 = _T_265 ? mimpid : _GEN_7418; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7434 = _T_265 ? mhartid : _GEN_7419; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7435 = _T_264 ? _medeleg_T_2 : medeleg; // @[decode.scala 472:28 596:39 605:38]
  wire [63:0] _GEN_7436 = _T_264 ? mideleg : _GEN_7420; // @[decode.scala 473:28 596:39]
  wire [63:0] _GEN_7437 = _T_264 ? mie : _GEN_7421; // @[decode.scala 474:28 596:39]
  wire [63:0] _GEN_7438 = _T_264 ? mtvec : _GEN_7422; // @[decode.scala 475:28 596:39]
  wire [63:0] _GEN_7439 = _T_264 ? mcounteren : _GEN_7423; // @[decode.scala 476:28 596:39]
  wire [63:0] _GEN_7440 = _T_264 ? mscratch : _GEN_7424; // @[decode.scala 477:28 596:39]
  wire [63:0] _GEN_7441 = _T_264 ? mepc : _GEN_7425; // @[decode.scala 478:28 596:39]
  wire [63:0] _GEN_7442 = _T_264 ? mcause : _GEN_7426; // @[decode.scala 479:28 596:39]
  wire [63:0] _GEN_7443 = _T_264 ? mtval : _GEN_7427; // @[decode.scala 480:28 596:39]
  wire [63:0] _GEN_7444 = _T_264 ? mip : _GEN_7428; // @[decode.scala 481:28 596:39]
  wire [63:0] _GEN_7445 = _T_264 ? pmpcfg0 : _GEN_7429; // @[decode.scala 482:28 596:39]
  wire [63:0] _GEN_7446 = _T_264 ? pmpaddr0 : _GEN_7430; // @[decode.scala 483:28 596:39]
  wire [63:0] _GEN_7447 = _T_264 ? mvendorid : _GEN_7431; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7448 = _T_264 ? marchid : _GEN_7432; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7449 = _T_264 ? mimpid : _GEN_7433; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7450 = _T_264 ? mhartid : _GEN_7434; // @[decode.scala 487:28 596:39]
  wire [126:0] _GEN_7451 = _T_263 ? {{63'd0}, _misa_T_4} : 127'h8000000000101101; // @[decode.scala 596:39 604:38 490:8]
  wire [63:0] _GEN_7452 = _T_263 ? medeleg : _GEN_7435; // @[decode.scala 472:28 596:39]
  wire [63:0] _GEN_7453 = _T_263 ? mideleg : _GEN_7436; // @[decode.scala 473:28 596:39]
  wire [63:0] _GEN_7454 = _T_263 ? mie : _GEN_7437; // @[decode.scala 474:28 596:39]
  wire [63:0] _GEN_7455 = _T_263 ? mtvec : _GEN_7438; // @[decode.scala 475:28 596:39]
  wire [63:0] _GEN_7456 = _T_263 ? mcounteren : _GEN_7439; // @[decode.scala 476:28 596:39]
  wire [63:0] _GEN_7457 = _T_263 ? mscratch : _GEN_7440; // @[decode.scala 477:28 596:39]
  wire [63:0] _GEN_7458 = _T_263 ? mepc : _GEN_7441; // @[decode.scala 478:28 596:39]
  wire [63:0] _GEN_7459 = _T_263 ? mcause : _GEN_7442; // @[decode.scala 479:28 596:39]
  wire [63:0] _GEN_7460 = _T_263 ? mtval : _GEN_7443; // @[decode.scala 480:28 596:39]
  wire [63:0] _GEN_7461 = _T_263 ? mip : _GEN_7444; // @[decode.scala 481:28 596:39]
  wire [63:0] _GEN_7462 = _T_263 ? pmpcfg0 : _GEN_7445; // @[decode.scala 482:28 596:39]
  wire [63:0] _GEN_7463 = _T_263 ? pmpaddr0 : _GEN_7446; // @[decode.scala 483:28 596:39]
  wire [63:0] _GEN_7464 = _T_263 ? mvendorid : _GEN_7447; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7465 = _T_263 ? marchid : _GEN_7448; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7466 = _T_263 ? mimpid : _GEN_7449; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7467 = _T_263 ? mhartid : _GEN_7450; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7468 = _T_262 ? _mstatus_T_4 : _mstatus_T_1; // @[decode.scala 489:11 596:39 603:38]
  wire [126:0] _GEN_7469 = _T_262 ? 127'h8000000000101101 : _GEN_7451; // @[decode.scala 596:39 490:8]
  wire [63:0] _GEN_7470 = _T_262 ? medeleg : _GEN_7452; // @[decode.scala 472:28 596:39]
  wire [63:0] _GEN_7471 = _T_262 ? mideleg : _GEN_7453; // @[decode.scala 473:28 596:39]
  wire [63:0] _GEN_7472 = _T_262 ? mie : _GEN_7454; // @[decode.scala 474:28 596:39]
  wire [63:0] _GEN_7473 = _T_262 ? mtvec : _GEN_7455; // @[decode.scala 475:28 596:39]
  wire [63:0] _GEN_7474 = _T_262 ? mcounteren : _GEN_7456; // @[decode.scala 476:28 596:39]
  wire [63:0] _GEN_7475 = _T_262 ? mscratch : _GEN_7457; // @[decode.scala 477:28 596:39]
  wire [63:0] _GEN_7476 = _T_262 ? mepc : _GEN_7458; // @[decode.scala 478:28 596:39]
  wire [63:0] _GEN_7477 = _T_262 ? mcause : _GEN_7459; // @[decode.scala 479:28 596:39]
  wire [63:0] _GEN_7478 = _T_262 ? mtval : _GEN_7460; // @[decode.scala 480:28 596:39]
  wire [63:0] _GEN_7479 = _T_262 ? mip : _GEN_7461; // @[decode.scala 481:28 596:39]
  wire [63:0] _GEN_7480 = _T_262 ? pmpcfg0 : _GEN_7462; // @[decode.scala 482:28 596:39]
  wire [63:0] _GEN_7481 = _T_262 ? pmpaddr0 : _GEN_7463; // @[decode.scala 483:28 596:39]
  wire [63:0] _GEN_7482 = _T_262 ? mvendorid : _GEN_7464; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7483 = _T_262 ? marchid : _GEN_7465; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7484 = _T_262 ? mimpid : _GEN_7466; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7485 = _T_262 ? mhartid : _GEN_7467; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7486 = _T_261 ? _satp_T_2 : satp; // @[decode.scala 469:28 596:39 602:38]
  wire [63:0] _GEN_7487 = _T_261 ? _mstatus_T_1 : _GEN_7468; // @[decode.scala 489:11 596:39]
  wire [126:0] _GEN_7488 = _T_261 ? 127'h8000000000101101 : _GEN_7469; // @[decode.scala 596:39 490:8]
  wire [63:0] _GEN_7489 = _T_261 ? medeleg : _GEN_7470; // @[decode.scala 472:28 596:39]
  wire [63:0] _GEN_7490 = _T_261 ? mideleg : _GEN_7471; // @[decode.scala 473:28 596:39]
  wire [63:0] _GEN_7491 = _T_261 ? mie : _GEN_7472; // @[decode.scala 474:28 596:39]
  wire [63:0] _GEN_7492 = _T_261 ? mtvec : _GEN_7473; // @[decode.scala 475:28 596:39]
  wire [63:0] _GEN_7493 = _T_261 ? mcounteren : _GEN_7474; // @[decode.scala 476:28 596:39]
  wire [63:0] _GEN_7494 = _T_261 ? mscratch : _GEN_7475; // @[decode.scala 477:28 596:39]
  wire [63:0] _GEN_7495 = _T_261 ? mepc : _GEN_7476; // @[decode.scala 478:28 596:39]
  wire [63:0] _GEN_7496 = _T_261 ? mcause : _GEN_7477; // @[decode.scala 479:28 596:39]
  wire [63:0] _GEN_7497 = _T_261 ? mtval : _GEN_7478; // @[decode.scala 480:28 596:39]
  wire [63:0] _GEN_7498 = _T_261 ? mip : _GEN_7479; // @[decode.scala 481:28 596:39]
  wire [63:0] _GEN_7499 = _T_261 ? pmpcfg0 : _GEN_7480; // @[decode.scala 482:28 596:39]
  wire [63:0] _GEN_7500 = _T_261 ? pmpaddr0 : _GEN_7481; // @[decode.scala 483:28 596:39]
  wire [63:0] _GEN_7501 = _T_261 ? mvendorid : _GEN_7482; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7502 = _T_261 ? marchid : _GEN_7483; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7503 = _T_261 ? mimpid : _GEN_7484; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7504 = _T_261 ? mhartid : _GEN_7485; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7505 = _T_260 ? _scounteren_T_2 : scounteren; // @[decode.scala 468:28 596:39 601:38]
  wire [63:0] _GEN_7506 = _T_260 ? satp : _GEN_7486; // @[decode.scala 469:28 596:39]
  wire [63:0] _GEN_7507 = _T_260 ? _mstatus_T_1 : _GEN_7487; // @[decode.scala 489:11 596:39]
  wire [126:0] _GEN_7508 = _T_260 ? 127'h8000000000101101 : _GEN_7488; // @[decode.scala 596:39 490:8]
  wire [63:0] _GEN_7509 = _T_260 ? medeleg : _GEN_7489; // @[decode.scala 472:28 596:39]
  wire [63:0] _GEN_7510 = _T_260 ? mideleg : _GEN_7490; // @[decode.scala 473:28 596:39]
  wire [63:0] _GEN_7511 = _T_260 ? mie : _GEN_7491; // @[decode.scala 474:28 596:39]
  wire [63:0] _GEN_7512 = _T_260 ? mtvec : _GEN_7492; // @[decode.scala 475:28 596:39]
  wire [63:0] _GEN_7513 = _T_260 ? mcounteren : _GEN_7493; // @[decode.scala 476:28 596:39]
  wire [63:0] _GEN_7514 = _T_260 ? mscratch : _GEN_7494; // @[decode.scala 477:28 596:39]
  wire [63:0] _GEN_7515 = _T_260 ? mepc : _GEN_7495; // @[decode.scala 478:28 596:39]
  wire [63:0] _GEN_7516 = _T_260 ? mcause : _GEN_7496; // @[decode.scala 479:28 596:39]
  wire [63:0] _GEN_7517 = _T_260 ? mtval : _GEN_7497; // @[decode.scala 480:28 596:39]
  wire [63:0] _GEN_7518 = _T_260 ? mip : _GEN_7498; // @[decode.scala 481:28 596:39]
  wire [63:0] _GEN_7519 = _T_260 ? pmpcfg0 : _GEN_7499; // @[decode.scala 482:28 596:39]
  wire [63:0] _GEN_7520 = _T_260 ? pmpaddr0 : _GEN_7500; // @[decode.scala 483:28 596:39]
  wire [63:0] _GEN_7521 = _T_260 ? mvendorid : _GEN_7501; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7522 = _T_260 ? marchid : _GEN_7502; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7523 = _T_260 ? mimpid : _GEN_7503; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7524 = _T_260 ? mhartid : _GEN_7504; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7525 = _T_259 ? _ucause_T_2 : ucause; // @[decode.scala 467:28 596:39 600:38]
  wire [63:0] _GEN_7526 = _T_259 ? scounteren : _GEN_7505; // @[decode.scala 468:28 596:39]
  wire [63:0] _GEN_7527 = _T_259 ? satp : _GEN_7506; // @[decode.scala 469:28 596:39]
  wire [63:0] _GEN_7528 = _T_259 ? _mstatus_T_1 : _GEN_7507; // @[decode.scala 489:11 596:39]
  wire [126:0] _GEN_7529 = _T_259 ? 127'h8000000000101101 : _GEN_7508; // @[decode.scala 596:39 490:8]
  wire [63:0] _GEN_7530 = _T_259 ? medeleg : _GEN_7509; // @[decode.scala 472:28 596:39]
  wire [63:0] _GEN_7531 = _T_259 ? mideleg : _GEN_7510; // @[decode.scala 473:28 596:39]
  wire [63:0] _GEN_7532 = _T_259 ? mie : _GEN_7511; // @[decode.scala 474:28 596:39]
  wire [63:0] _GEN_7533 = _T_259 ? mtvec : _GEN_7512; // @[decode.scala 475:28 596:39]
  wire [63:0] _GEN_7534 = _T_259 ? mcounteren : _GEN_7513; // @[decode.scala 476:28 596:39]
  wire [63:0] _GEN_7535 = _T_259 ? mscratch : _GEN_7514; // @[decode.scala 477:28 596:39]
  wire [63:0] _GEN_7536 = _T_259 ? mepc : _GEN_7515; // @[decode.scala 478:28 596:39]
  wire [63:0] _GEN_7537 = _T_259 ? mcause : _GEN_7516; // @[decode.scala 479:28 596:39]
  wire [63:0] _GEN_7538 = _T_259 ? mtval : _GEN_7517; // @[decode.scala 480:28 596:39]
  wire [63:0] _GEN_7539 = _T_259 ? mip : _GEN_7518; // @[decode.scala 481:28 596:39]
  wire [63:0] _GEN_7540 = _T_259 ? pmpcfg0 : _GEN_7519; // @[decode.scala 482:28 596:39]
  wire [63:0] _GEN_7541 = _T_259 ? pmpaddr0 : _GEN_7520; // @[decode.scala 483:28 596:39]
  wire [63:0] _GEN_7542 = _T_259 ? mvendorid : _GEN_7521; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7543 = _T_259 ? marchid : _GEN_7522; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7544 = _T_259 ? mimpid : _GEN_7523; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7545 = _T_259 ? mhartid : _GEN_7524; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7546 = _T_258 ? _uepc_T_2 : uepc; // @[decode.scala 466:28 596:39 599:38]
  wire [63:0] _GEN_7547 = _T_258 ? ucause : _GEN_7525; // @[decode.scala 467:28 596:39]
  wire [63:0] _GEN_7548 = _T_258 ? scounteren : _GEN_7526; // @[decode.scala 468:28 596:39]
  wire [63:0] _GEN_7549 = _T_258 ? satp : _GEN_7527; // @[decode.scala 469:28 596:39]
  wire [63:0] _GEN_7550 = _T_258 ? _mstatus_T_1 : _GEN_7528; // @[decode.scala 489:11 596:39]
  wire [126:0] _GEN_7551 = _T_258 ? 127'h8000000000101101 : _GEN_7529; // @[decode.scala 596:39 490:8]
  wire [63:0] _GEN_7552 = _T_258 ? medeleg : _GEN_7530; // @[decode.scala 472:28 596:39]
  wire [63:0] _GEN_7553 = _T_258 ? mideleg : _GEN_7531; // @[decode.scala 473:28 596:39]
  wire [63:0] _GEN_7554 = _T_258 ? mie : _GEN_7532; // @[decode.scala 474:28 596:39]
  wire [63:0] _GEN_7555 = _T_258 ? mtvec : _GEN_7533; // @[decode.scala 475:28 596:39]
  wire [63:0] _GEN_7556 = _T_258 ? mcounteren : _GEN_7534; // @[decode.scala 476:28 596:39]
  wire [63:0] _GEN_7557 = _T_258 ? mscratch : _GEN_7535; // @[decode.scala 477:28 596:39]
  wire [63:0] _GEN_7558 = _T_258 ? mepc : _GEN_7536; // @[decode.scala 478:28 596:39]
  wire [63:0] _GEN_7559 = _T_258 ? mcause : _GEN_7537; // @[decode.scala 479:28 596:39]
  wire [63:0] _GEN_7560 = _T_258 ? mtval : _GEN_7538; // @[decode.scala 480:28 596:39]
  wire [63:0] _GEN_7561 = _T_258 ? mip : _GEN_7539; // @[decode.scala 481:28 596:39]
  wire [63:0] _GEN_7562 = _T_258 ? pmpcfg0 : _GEN_7540; // @[decode.scala 482:28 596:39]
  wire [63:0] _GEN_7563 = _T_258 ? pmpaddr0 : _GEN_7541; // @[decode.scala 483:28 596:39]
  wire [63:0] _GEN_7564 = _T_258 ? mvendorid : _GEN_7542; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7565 = _T_258 ? marchid : _GEN_7543; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7566 = _T_258 ? mimpid : _GEN_7544; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7567 = _T_258 ? mhartid : _GEN_7545; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7568 = _T_257 ? _utvec_T_2 : utvec; // @[decode.scala 465:28 596:39 598:38]
  wire [63:0] _GEN_7569 = _T_257 ? uepc : _GEN_7546; // @[decode.scala 466:28 596:39]
  wire [63:0] _GEN_7570 = _T_257 ? ucause : _GEN_7547; // @[decode.scala 467:28 596:39]
  wire [63:0] _GEN_7571 = _T_257 ? scounteren : _GEN_7548; // @[decode.scala 468:28 596:39]
  wire [63:0] _GEN_7572 = _T_257 ? satp : _GEN_7549; // @[decode.scala 469:28 596:39]
  wire [63:0] _GEN_7573 = _T_257 ? _mstatus_T_1 : _GEN_7550; // @[decode.scala 489:11 596:39]
  wire [126:0] _GEN_7574 = _T_257 ? 127'h8000000000101101 : _GEN_7551; // @[decode.scala 596:39 490:8]
  wire [63:0] _GEN_7575 = _T_257 ? medeleg : _GEN_7552; // @[decode.scala 472:28 596:39]
  wire [63:0] _GEN_7576 = _T_257 ? mideleg : _GEN_7553; // @[decode.scala 473:28 596:39]
  wire [63:0] _GEN_7577 = _T_257 ? mie : _GEN_7554; // @[decode.scala 474:28 596:39]
  wire [63:0] _GEN_7578 = _T_257 ? mtvec : _GEN_7555; // @[decode.scala 475:28 596:39]
  wire [63:0] _GEN_7579 = _T_257 ? mcounteren : _GEN_7556; // @[decode.scala 476:28 596:39]
  wire [63:0] _GEN_7580 = _T_257 ? mscratch : _GEN_7557; // @[decode.scala 477:28 596:39]
  wire [63:0] _GEN_7581 = _T_257 ? mepc : _GEN_7558; // @[decode.scala 478:28 596:39]
  wire [63:0] _GEN_7582 = _T_257 ? mcause : _GEN_7559; // @[decode.scala 479:28 596:39]
  wire [63:0] _GEN_7583 = _T_257 ? mtval : _GEN_7560; // @[decode.scala 480:28 596:39]
  wire [63:0] _GEN_7584 = _T_257 ? mip : _GEN_7561; // @[decode.scala 481:28 596:39]
  wire [63:0] _GEN_7585 = _T_257 ? pmpcfg0 : _GEN_7562; // @[decode.scala 482:28 596:39]
  wire [63:0] _GEN_7586 = _T_257 ? pmpaddr0 : _GEN_7563; // @[decode.scala 483:28 596:39]
  wire [63:0] _GEN_7587 = _T_257 ? mvendorid : _GEN_7564; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7588 = _T_257 ? marchid : _GEN_7565; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7589 = _T_257 ? mimpid : _GEN_7566; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7590 = _T_257 ? mhartid : _GEN_7567; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7591 = _T_256 ? _ustatus_T_2 : ustatus; // @[decode.scala 464:28 596:39 597:38]
  wire [63:0] _GEN_7592 = _T_256 ? utvec : _GEN_7568; // @[decode.scala 465:28 596:39]
  wire [63:0] _GEN_7593 = _T_256 ? uepc : _GEN_7569; // @[decode.scala 466:28 596:39]
  wire [63:0] _GEN_7594 = _T_256 ? ucause : _GEN_7570; // @[decode.scala 467:28 596:39]
  wire [63:0] _GEN_7595 = _T_256 ? scounteren : _GEN_7571; // @[decode.scala 468:28 596:39]
  wire [63:0] _GEN_7596 = _T_256 ? satp : _GEN_7572; // @[decode.scala 469:28 596:39]
  wire [63:0] _GEN_7597 = _T_256 ? _mstatus_T_1 : _GEN_7573; // @[decode.scala 489:11 596:39]
  wire [126:0] _GEN_7598 = _T_256 ? 127'h8000000000101101 : _GEN_7574; // @[decode.scala 596:39 490:8]
  wire [63:0] _GEN_7599 = _T_256 ? medeleg : _GEN_7575; // @[decode.scala 472:28 596:39]
  wire [63:0] _GEN_7600 = _T_256 ? mideleg : _GEN_7576; // @[decode.scala 473:28 596:39]
  wire [63:0] _GEN_7601 = _T_256 ? mie : _GEN_7577; // @[decode.scala 474:28 596:39]
  wire [63:0] _GEN_7602 = _T_256 ? mtvec : _GEN_7578; // @[decode.scala 475:28 596:39]
  wire [63:0] _GEN_7603 = _T_256 ? mcounteren : _GEN_7579; // @[decode.scala 476:28 596:39]
  wire [63:0] _GEN_7604 = _T_256 ? mscratch : _GEN_7580; // @[decode.scala 477:28 596:39]
  wire [63:0] _GEN_7605 = _T_256 ? mepc : _GEN_7581; // @[decode.scala 478:28 596:39]
  wire [63:0] _GEN_7606 = _T_256 ? mcause : _GEN_7582; // @[decode.scala 479:28 596:39]
  wire [63:0] _GEN_7607 = _T_256 ? mtval : _GEN_7583; // @[decode.scala 480:28 596:39]
  wire [63:0] _GEN_7608 = _T_256 ? mip : _GEN_7584; // @[decode.scala 481:28 596:39]
  wire [63:0] _GEN_7609 = _T_256 ? pmpcfg0 : _GEN_7585; // @[decode.scala 482:28 596:39]
  wire [63:0] _GEN_7610 = _T_256 ? pmpaddr0 : _GEN_7586; // @[decode.scala 483:28 596:39]
  wire [63:0] _GEN_7611 = _T_256 ? mvendorid : _GEN_7587; // @[decode.scala 484:28 596:39]
  wire [63:0] _GEN_7612 = _T_256 ? marchid : _GEN_7588; // @[decode.scala 485:28 596:39]
  wire [63:0] _GEN_7613 = _T_256 ? mimpid : _GEN_7589; // @[decode.scala 486:28 596:39]
  wire [63:0] _GEN_7614 = _T_256 ? mhartid : _GEN_7590; // @[decode.scala 487:28 596:39]
  wire [63:0] _GEN_7615 = _T_279 ? csrImmReg : mhartid; // @[decode.scala 487:28 624:39 648:38]
  wire [63:0] _GEN_7616 = _T_278 ? csrImmReg : mimpid; // @[decode.scala 486:28 624:39 647:38]
  wire [63:0] _GEN_7617 = _T_278 ? mhartid : _GEN_7615; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7618 = _T_277 ? csrImmReg : marchid; // @[decode.scala 485:28 624:39 646:38]
  wire [63:0] _GEN_7619 = _T_277 ? mimpid : _GEN_7616; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7620 = _T_277 ? mhartid : _GEN_7617; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7621 = _T_276 ? csrImmReg : mvendorid; // @[decode.scala 484:28 624:39 645:38]
  wire [63:0] _GEN_7622 = _T_276 ? marchid : _GEN_7618; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7623 = _T_276 ? mimpid : _GEN_7619; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7624 = _T_276 ? mhartid : _GEN_7620; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7625 = _T_275 ? csrImmReg : pmpaddr0; // @[decode.scala 483:28 624:39 644:38]
  wire [63:0] _GEN_7626 = _T_275 ? mvendorid : _GEN_7621; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7627 = _T_275 ? marchid : _GEN_7622; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7628 = _T_275 ? mimpid : _GEN_7623; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7629 = _T_275 ? mhartid : _GEN_7624; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7630 = _T_274 ? csrImmReg : pmpcfg0; // @[decode.scala 482:28 624:39 643:38]
  wire [63:0] _GEN_7631 = _T_274 ? pmpaddr0 : _GEN_7625; // @[decode.scala 483:28 624:39]
  wire [63:0] _GEN_7632 = _T_274 ? mvendorid : _GEN_7626; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7633 = _T_274 ? marchid : _GEN_7627; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7634 = _T_274 ? mimpid : _GEN_7628; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7635 = _T_274 ? mhartid : _GEN_7629; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7636 = _T_273 ? csrImmReg : mip; // @[decode.scala 481:28 624:39 642:38]
  wire [63:0] _GEN_7637 = _T_273 ? pmpcfg0 : _GEN_7630; // @[decode.scala 482:28 624:39]
  wire [63:0] _GEN_7638 = _T_273 ? pmpaddr0 : _GEN_7631; // @[decode.scala 483:28 624:39]
  wire [63:0] _GEN_7639 = _T_273 ? mvendorid : _GEN_7632; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7640 = _T_273 ? marchid : _GEN_7633; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7641 = _T_273 ? mimpid : _GEN_7634; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7642 = _T_273 ? mhartid : _GEN_7635; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7643 = _T_272 ? csrImmReg : mtval; // @[decode.scala 480:28 624:39 641:38]
  wire [63:0] _GEN_7644 = _T_272 ? mip : _GEN_7636; // @[decode.scala 481:28 624:39]
  wire [63:0] _GEN_7645 = _T_272 ? pmpcfg0 : _GEN_7637; // @[decode.scala 482:28 624:39]
  wire [63:0] _GEN_7646 = _T_272 ? pmpaddr0 : _GEN_7638; // @[decode.scala 483:28 624:39]
  wire [63:0] _GEN_7647 = _T_272 ? mvendorid : _GEN_7639; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7648 = _T_272 ? marchid : _GEN_7640; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7649 = _T_272 ? mimpid : _GEN_7641; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7650 = _T_272 ? mhartid : _GEN_7642; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7651 = _T_271 ? csrImmReg : mcause; // @[decode.scala 479:28 624:39 640:38]
  wire [63:0] _GEN_7652 = _T_271 ? mtval : _GEN_7643; // @[decode.scala 480:28 624:39]
  wire [63:0] _GEN_7653 = _T_271 ? mip : _GEN_7644; // @[decode.scala 481:28 624:39]
  wire [63:0] _GEN_7654 = _T_271 ? pmpcfg0 : _GEN_7645; // @[decode.scala 482:28 624:39]
  wire [63:0] _GEN_7655 = _T_271 ? pmpaddr0 : _GEN_7646; // @[decode.scala 483:28 624:39]
  wire [63:0] _GEN_7656 = _T_271 ? mvendorid : _GEN_7647; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7657 = _T_271 ? marchid : _GEN_7648; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7658 = _T_271 ? mimpid : _GEN_7649; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7659 = _T_271 ? mhartid : _GEN_7650; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7660 = _T_270 ? csrImmReg : mepc; // @[decode.scala 478:28 624:39 639:38]
  wire [63:0] _GEN_7661 = _T_270 ? mcause : _GEN_7651; // @[decode.scala 479:28 624:39]
  wire [63:0] _GEN_7662 = _T_270 ? mtval : _GEN_7652; // @[decode.scala 480:28 624:39]
  wire [63:0] _GEN_7663 = _T_270 ? mip : _GEN_7653; // @[decode.scala 481:28 624:39]
  wire [63:0] _GEN_7664 = _T_270 ? pmpcfg0 : _GEN_7654; // @[decode.scala 482:28 624:39]
  wire [63:0] _GEN_7665 = _T_270 ? pmpaddr0 : _GEN_7655; // @[decode.scala 483:28 624:39]
  wire [63:0] _GEN_7666 = _T_270 ? mvendorid : _GEN_7656; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7667 = _T_270 ? marchid : _GEN_7657; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7668 = _T_270 ? mimpid : _GEN_7658; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7669 = _T_270 ? mhartid : _GEN_7659; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7670 = _T_269 ? csrImmReg : mscratch; // @[decode.scala 477:28 624:39 638:38]
  wire [63:0] _GEN_7671 = _T_269 ? mepc : _GEN_7660; // @[decode.scala 478:28 624:39]
  wire [63:0] _GEN_7672 = _T_269 ? mcause : _GEN_7661; // @[decode.scala 479:28 624:39]
  wire [63:0] _GEN_7673 = _T_269 ? mtval : _GEN_7662; // @[decode.scala 480:28 624:39]
  wire [63:0] _GEN_7674 = _T_269 ? mip : _GEN_7663; // @[decode.scala 481:28 624:39]
  wire [63:0] _GEN_7675 = _T_269 ? pmpcfg0 : _GEN_7664; // @[decode.scala 482:28 624:39]
  wire [63:0] _GEN_7676 = _T_269 ? pmpaddr0 : _GEN_7665; // @[decode.scala 483:28 624:39]
  wire [63:0] _GEN_7677 = _T_269 ? mvendorid : _GEN_7666; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7678 = _T_269 ? marchid : _GEN_7667; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7679 = _T_269 ? mimpid : _GEN_7668; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7680 = _T_269 ? mhartid : _GEN_7669; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7681 = _T_268 ? csrImmReg : mcounteren; // @[decode.scala 476:28 624:39 637:38]
  wire [63:0] _GEN_7682 = _T_268 ? mscratch : _GEN_7670; // @[decode.scala 477:28 624:39]
  wire [63:0] _GEN_7683 = _T_268 ? mepc : _GEN_7671; // @[decode.scala 478:28 624:39]
  wire [63:0] _GEN_7684 = _T_268 ? mcause : _GEN_7672; // @[decode.scala 479:28 624:39]
  wire [63:0] _GEN_7685 = _T_268 ? mtval : _GEN_7673; // @[decode.scala 480:28 624:39]
  wire [63:0] _GEN_7686 = _T_268 ? mip : _GEN_7674; // @[decode.scala 481:28 624:39]
  wire [63:0] _GEN_7687 = _T_268 ? pmpcfg0 : _GEN_7675; // @[decode.scala 482:28 624:39]
  wire [63:0] _GEN_7688 = _T_268 ? pmpaddr0 : _GEN_7676; // @[decode.scala 483:28 624:39]
  wire [63:0] _GEN_7689 = _T_268 ? mvendorid : _GEN_7677; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7690 = _T_268 ? marchid : _GEN_7678; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7691 = _T_268 ? mimpid : _GEN_7679; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7692 = _T_268 ? mhartid : _GEN_7680; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7693 = _T_267 ? csrImmReg : mtvec; // @[decode.scala 475:28 624:39 636:38]
  wire [63:0] _GEN_7694 = _T_267 ? mcounteren : _GEN_7681; // @[decode.scala 476:28 624:39]
  wire [63:0] _GEN_7695 = _T_267 ? mscratch : _GEN_7682; // @[decode.scala 477:28 624:39]
  wire [63:0] _GEN_7696 = _T_267 ? mepc : _GEN_7683; // @[decode.scala 478:28 624:39]
  wire [63:0] _GEN_7697 = _T_267 ? mcause : _GEN_7684; // @[decode.scala 479:28 624:39]
  wire [63:0] _GEN_7698 = _T_267 ? mtval : _GEN_7685; // @[decode.scala 480:28 624:39]
  wire [63:0] _GEN_7699 = _T_267 ? mip : _GEN_7686; // @[decode.scala 481:28 624:39]
  wire [63:0] _GEN_7700 = _T_267 ? pmpcfg0 : _GEN_7687; // @[decode.scala 482:28 624:39]
  wire [63:0] _GEN_7701 = _T_267 ? pmpaddr0 : _GEN_7688; // @[decode.scala 483:28 624:39]
  wire [63:0] _GEN_7702 = _T_267 ? mvendorid : _GEN_7689; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7703 = _T_267 ? marchid : _GEN_7690; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7704 = _T_267 ? mimpid : _GEN_7691; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7705 = _T_267 ? mhartid : _GEN_7692; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7706 = _T_266 ? csrImmReg : mie; // @[decode.scala 474:28 624:39 635:38]
  wire [63:0] _GEN_7707 = _T_266 ? mtvec : _GEN_7693; // @[decode.scala 475:28 624:39]
  wire [63:0] _GEN_7708 = _T_266 ? mcounteren : _GEN_7694; // @[decode.scala 476:28 624:39]
  wire [63:0] _GEN_7709 = _T_266 ? mscratch : _GEN_7695; // @[decode.scala 477:28 624:39]
  wire [63:0] _GEN_7710 = _T_266 ? mepc : _GEN_7696; // @[decode.scala 478:28 624:39]
  wire [63:0] _GEN_7711 = _T_266 ? mcause : _GEN_7697; // @[decode.scala 479:28 624:39]
  wire [63:0] _GEN_7712 = _T_266 ? mtval : _GEN_7698; // @[decode.scala 480:28 624:39]
  wire [63:0] _GEN_7713 = _T_266 ? mip : _GEN_7699; // @[decode.scala 481:28 624:39]
  wire [63:0] _GEN_7714 = _T_266 ? pmpcfg0 : _GEN_7700; // @[decode.scala 482:28 624:39]
  wire [63:0] _GEN_7715 = _T_266 ? pmpaddr0 : _GEN_7701; // @[decode.scala 483:28 624:39]
  wire [63:0] _GEN_7716 = _T_266 ? mvendorid : _GEN_7702; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7717 = _T_266 ? marchid : _GEN_7703; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7718 = _T_266 ? mimpid : _GEN_7704; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7719 = _T_266 ? mhartid : _GEN_7705; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7720 = _T_265 ? csrImmReg : mideleg; // @[decode.scala 473:28 624:39 634:38]
  wire [63:0] _GEN_7721 = _T_265 ? mie : _GEN_7706; // @[decode.scala 474:28 624:39]
  wire [63:0] _GEN_7722 = _T_265 ? mtvec : _GEN_7707; // @[decode.scala 475:28 624:39]
  wire [63:0] _GEN_7723 = _T_265 ? mcounteren : _GEN_7708; // @[decode.scala 476:28 624:39]
  wire [63:0] _GEN_7724 = _T_265 ? mscratch : _GEN_7709; // @[decode.scala 477:28 624:39]
  wire [63:0] _GEN_7725 = _T_265 ? mepc : _GEN_7710; // @[decode.scala 478:28 624:39]
  wire [63:0] _GEN_7726 = _T_265 ? mcause : _GEN_7711; // @[decode.scala 479:28 624:39]
  wire [63:0] _GEN_7727 = _T_265 ? mtval : _GEN_7712; // @[decode.scala 480:28 624:39]
  wire [63:0] _GEN_7728 = _T_265 ? mip : _GEN_7713; // @[decode.scala 481:28 624:39]
  wire [63:0] _GEN_7729 = _T_265 ? pmpcfg0 : _GEN_7714; // @[decode.scala 482:28 624:39]
  wire [63:0] _GEN_7730 = _T_265 ? pmpaddr0 : _GEN_7715; // @[decode.scala 483:28 624:39]
  wire [63:0] _GEN_7731 = _T_265 ? mvendorid : _GEN_7716; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7732 = _T_265 ? marchid : _GEN_7717; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7733 = _T_265 ? mimpid : _GEN_7718; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7734 = _T_265 ? mhartid : _GEN_7719; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7735 = _T_264 ? csrImmReg : medeleg; // @[decode.scala 472:28 624:39 633:38]
  wire [63:0] _GEN_7736 = _T_264 ? mideleg : _GEN_7720; // @[decode.scala 473:28 624:39]
  wire [63:0] _GEN_7737 = _T_264 ? mie : _GEN_7721; // @[decode.scala 474:28 624:39]
  wire [63:0] _GEN_7738 = _T_264 ? mtvec : _GEN_7722; // @[decode.scala 475:28 624:39]
  wire [63:0] _GEN_7739 = _T_264 ? mcounteren : _GEN_7723; // @[decode.scala 476:28 624:39]
  wire [63:0] _GEN_7740 = _T_264 ? mscratch : _GEN_7724; // @[decode.scala 477:28 624:39]
  wire [63:0] _GEN_7741 = _T_264 ? mepc : _GEN_7725; // @[decode.scala 478:28 624:39]
  wire [63:0] _GEN_7742 = _T_264 ? mcause : _GEN_7726; // @[decode.scala 479:28 624:39]
  wire [63:0] _GEN_7743 = _T_264 ? mtval : _GEN_7727; // @[decode.scala 480:28 624:39]
  wire [63:0] _GEN_7744 = _T_264 ? mip : _GEN_7728; // @[decode.scala 481:28 624:39]
  wire [63:0] _GEN_7745 = _T_264 ? pmpcfg0 : _GEN_7729; // @[decode.scala 482:28 624:39]
  wire [63:0] _GEN_7746 = _T_264 ? pmpaddr0 : _GEN_7730; // @[decode.scala 483:28 624:39]
  wire [63:0] _GEN_7747 = _T_264 ? mvendorid : _GEN_7731; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7748 = _T_264 ? marchid : _GEN_7732; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7749 = _T_264 ? mimpid : _GEN_7733; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7750 = _T_264 ? mhartid : _GEN_7734; // @[decode.scala 487:28 624:39]
  wire [126:0] _GEN_7751 = _T_263 ? {{63'd0}, csrImmReg} : 127'h8000000000101101; // @[decode.scala 624:39 632:38 490:8]
  wire [63:0] _GEN_7752 = _T_263 ? medeleg : _GEN_7735; // @[decode.scala 472:28 624:39]
  wire [63:0] _GEN_7753 = _T_263 ? mideleg : _GEN_7736; // @[decode.scala 473:28 624:39]
  wire [63:0] _GEN_7754 = _T_263 ? mie : _GEN_7737; // @[decode.scala 474:28 624:39]
  wire [63:0] _GEN_7755 = _T_263 ? mtvec : _GEN_7738; // @[decode.scala 475:28 624:39]
  wire [63:0] _GEN_7756 = _T_263 ? mcounteren : _GEN_7739; // @[decode.scala 476:28 624:39]
  wire [63:0] _GEN_7757 = _T_263 ? mscratch : _GEN_7740; // @[decode.scala 477:28 624:39]
  wire [63:0] _GEN_7758 = _T_263 ? mepc : _GEN_7741; // @[decode.scala 478:28 624:39]
  wire [63:0] _GEN_7759 = _T_263 ? mcause : _GEN_7742; // @[decode.scala 479:28 624:39]
  wire [63:0] _GEN_7760 = _T_263 ? mtval : _GEN_7743; // @[decode.scala 480:28 624:39]
  wire [63:0] _GEN_7761 = _T_263 ? mip : _GEN_7744; // @[decode.scala 481:28 624:39]
  wire [63:0] _GEN_7762 = _T_263 ? pmpcfg0 : _GEN_7745; // @[decode.scala 482:28 624:39]
  wire [63:0] _GEN_7763 = _T_263 ? pmpaddr0 : _GEN_7746; // @[decode.scala 483:28 624:39]
  wire [63:0] _GEN_7764 = _T_263 ? mvendorid : _GEN_7747; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7765 = _T_263 ? marchid : _GEN_7748; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7766 = _T_263 ? mimpid : _GEN_7749; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7767 = _T_263 ? mhartid : _GEN_7750; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7768 = _T_262 ? csrImmReg : _mstatus_T_1; // @[decode.scala 489:11 624:39 631:38]
  wire [126:0] _GEN_7769 = _T_262 ? 127'h8000000000101101 : _GEN_7751; // @[decode.scala 624:39 490:8]
  wire [63:0] _GEN_7770 = _T_262 ? medeleg : _GEN_7752; // @[decode.scala 472:28 624:39]
  wire [63:0] _GEN_7771 = _T_262 ? mideleg : _GEN_7753; // @[decode.scala 473:28 624:39]
  wire [63:0] _GEN_7772 = _T_262 ? mie : _GEN_7754; // @[decode.scala 474:28 624:39]
  wire [63:0] _GEN_7773 = _T_262 ? mtvec : _GEN_7755; // @[decode.scala 475:28 624:39]
  wire [63:0] _GEN_7774 = _T_262 ? mcounteren : _GEN_7756; // @[decode.scala 476:28 624:39]
  wire [63:0] _GEN_7775 = _T_262 ? mscratch : _GEN_7757; // @[decode.scala 477:28 624:39]
  wire [63:0] _GEN_7776 = _T_262 ? mepc : _GEN_7758; // @[decode.scala 478:28 624:39]
  wire [63:0] _GEN_7777 = _T_262 ? mcause : _GEN_7759; // @[decode.scala 479:28 624:39]
  wire [63:0] _GEN_7778 = _T_262 ? mtval : _GEN_7760; // @[decode.scala 480:28 624:39]
  wire [63:0] _GEN_7779 = _T_262 ? mip : _GEN_7761; // @[decode.scala 481:28 624:39]
  wire [63:0] _GEN_7780 = _T_262 ? pmpcfg0 : _GEN_7762; // @[decode.scala 482:28 624:39]
  wire [63:0] _GEN_7781 = _T_262 ? pmpaddr0 : _GEN_7763; // @[decode.scala 483:28 624:39]
  wire [63:0] _GEN_7782 = _T_262 ? mvendorid : _GEN_7764; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7783 = _T_262 ? marchid : _GEN_7765; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7784 = _T_262 ? mimpid : _GEN_7766; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7785 = _T_262 ? mhartid : _GEN_7767; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7786 = _T_261 ? csrImmReg : satp; // @[decode.scala 469:28 624:39 630:38]
  wire [63:0] _GEN_7787 = _T_261 ? _mstatus_T_1 : _GEN_7768; // @[decode.scala 489:11 624:39]
  wire [126:0] _GEN_7788 = _T_261 ? 127'h8000000000101101 : _GEN_7769; // @[decode.scala 624:39 490:8]
  wire [63:0] _GEN_7789 = _T_261 ? medeleg : _GEN_7770; // @[decode.scala 472:28 624:39]
  wire [63:0] _GEN_7790 = _T_261 ? mideleg : _GEN_7771; // @[decode.scala 473:28 624:39]
  wire [63:0] _GEN_7791 = _T_261 ? mie : _GEN_7772; // @[decode.scala 474:28 624:39]
  wire [63:0] _GEN_7792 = _T_261 ? mtvec : _GEN_7773; // @[decode.scala 475:28 624:39]
  wire [63:0] _GEN_7793 = _T_261 ? mcounteren : _GEN_7774; // @[decode.scala 476:28 624:39]
  wire [63:0] _GEN_7794 = _T_261 ? mscratch : _GEN_7775; // @[decode.scala 477:28 624:39]
  wire [63:0] _GEN_7795 = _T_261 ? mepc : _GEN_7776; // @[decode.scala 478:28 624:39]
  wire [63:0] _GEN_7796 = _T_261 ? mcause : _GEN_7777; // @[decode.scala 479:28 624:39]
  wire [63:0] _GEN_7797 = _T_261 ? mtval : _GEN_7778; // @[decode.scala 480:28 624:39]
  wire [63:0] _GEN_7798 = _T_261 ? mip : _GEN_7779; // @[decode.scala 481:28 624:39]
  wire [63:0] _GEN_7799 = _T_261 ? pmpcfg0 : _GEN_7780; // @[decode.scala 482:28 624:39]
  wire [63:0] _GEN_7800 = _T_261 ? pmpaddr0 : _GEN_7781; // @[decode.scala 483:28 624:39]
  wire [63:0] _GEN_7801 = _T_261 ? mvendorid : _GEN_7782; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7802 = _T_261 ? marchid : _GEN_7783; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7803 = _T_261 ? mimpid : _GEN_7784; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7804 = _T_261 ? mhartid : _GEN_7785; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7805 = _T_260 ? csrImmReg : scounteren; // @[decode.scala 468:28 624:39 629:38]
  wire [63:0] _GEN_7806 = _T_260 ? satp : _GEN_7786; // @[decode.scala 469:28 624:39]
  wire [63:0] _GEN_7807 = _T_260 ? _mstatus_T_1 : _GEN_7787; // @[decode.scala 489:11 624:39]
  wire [126:0] _GEN_7808 = _T_260 ? 127'h8000000000101101 : _GEN_7788; // @[decode.scala 624:39 490:8]
  wire [63:0] _GEN_7809 = _T_260 ? medeleg : _GEN_7789; // @[decode.scala 472:28 624:39]
  wire [63:0] _GEN_7810 = _T_260 ? mideleg : _GEN_7790; // @[decode.scala 473:28 624:39]
  wire [63:0] _GEN_7811 = _T_260 ? mie : _GEN_7791; // @[decode.scala 474:28 624:39]
  wire [63:0] _GEN_7812 = _T_260 ? mtvec : _GEN_7792; // @[decode.scala 475:28 624:39]
  wire [63:0] _GEN_7813 = _T_260 ? mcounteren : _GEN_7793; // @[decode.scala 476:28 624:39]
  wire [63:0] _GEN_7814 = _T_260 ? mscratch : _GEN_7794; // @[decode.scala 477:28 624:39]
  wire [63:0] _GEN_7815 = _T_260 ? mepc : _GEN_7795; // @[decode.scala 478:28 624:39]
  wire [63:0] _GEN_7816 = _T_260 ? mcause : _GEN_7796; // @[decode.scala 479:28 624:39]
  wire [63:0] _GEN_7817 = _T_260 ? mtval : _GEN_7797; // @[decode.scala 480:28 624:39]
  wire [63:0] _GEN_7818 = _T_260 ? mip : _GEN_7798; // @[decode.scala 481:28 624:39]
  wire [63:0] _GEN_7819 = _T_260 ? pmpcfg0 : _GEN_7799; // @[decode.scala 482:28 624:39]
  wire [63:0] _GEN_7820 = _T_260 ? pmpaddr0 : _GEN_7800; // @[decode.scala 483:28 624:39]
  wire [63:0] _GEN_7821 = _T_260 ? mvendorid : _GEN_7801; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7822 = _T_260 ? marchid : _GEN_7802; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7823 = _T_260 ? mimpid : _GEN_7803; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7824 = _T_260 ? mhartid : _GEN_7804; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7825 = _T_259 ? csrImmReg : ucause; // @[decode.scala 467:28 624:39 628:38]
  wire [63:0] _GEN_7826 = _T_259 ? scounteren : _GEN_7805; // @[decode.scala 468:28 624:39]
  wire [63:0] _GEN_7827 = _T_259 ? satp : _GEN_7806; // @[decode.scala 469:28 624:39]
  wire [63:0] _GEN_7828 = _T_259 ? _mstatus_T_1 : _GEN_7807; // @[decode.scala 489:11 624:39]
  wire [126:0] _GEN_7829 = _T_259 ? 127'h8000000000101101 : _GEN_7808; // @[decode.scala 624:39 490:8]
  wire [63:0] _GEN_7830 = _T_259 ? medeleg : _GEN_7809; // @[decode.scala 472:28 624:39]
  wire [63:0] _GEN_7831 = _T_259 ? mideleg : _GEN_7810; // @[decode.scala 473:28 624:39]
  wire [63:0] _GEN_7832 = _T_259 ? mie : _GEN_7811; // @[decode.scala 474:28 624:39]
  wire [63:0] _GEN_7833 = _T_259 ? mtvec : _GEN_7812; // @[decode.scala 475:28 624:39]
  wire [63:0] _GEN_7834 = _T_259 ? mcounteren : _GEN_7813; // @[decode.scala 476:28 624:39]
  wire [63:0] _GEN_7835 = _T_259 ? mscratch : _GEN_7814; // @[decode.scala 477:28 624:39]
  wire [63:0] _GEN_7836 = _T_259 ? mepc : _GEN_7815; // @[decode.scala 478:28 624:39]
  wire [63:0] _GEN_7837 = _T_259 ? mcause : _GEN_7816; // @[decode.scala 479:28 624:39]
  wire [63:0] _GEN_7838 = _T_259 ? mtval : _GEN_7817; // @[decode.scala 480:28 624:39]
  wire [63:0] _GEN_7839 = _T_259 ? mip : _GEN_7818; // @[decode.scala 481:28 624:39]
  wire [63:0] _GEN_7840 = _T_259 ? pmpcfg0 : _GEN_7819; // @[decode.scala 482:28 624:39]
  wire [63:0] _GEN_7841 = _T_259 ? pmpaddr0 : _GEN_7820; // @[decode.scala 483:28 624:39]
  wire [63:0] _GEN_7842 = _T_259 ? mvendorid : _GEN_7821; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7843 = _T_259 ? marchid : _GEN_7822; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7844 = _T_259 ? mimpid : _GEN_7823; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7845 = _T_259 ? mhartid : _GEN_7824; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7846 = _T_258 ? csrImmReg : uepc; // @[decode.scala 466:28 624:39 627:38]
  wire [63:0] _GEN_7847 = _T_258 ? ucause : _GEN_7825; // @[decode.scala 467:28 624:39]
  wire [63:0] _GEN_7848 = _T_258 ? scounteren : _GEN_7826; // @[decode.scala 468:28 624:39]
  wire [63:0] _GEN_7849 = _T_258 ? satp : _GEN_7827; // @[decode.scala 469:28 624:39]
  wire [63:0] _GEN_7850 = _T_258 ? _mstatus_T_1 : _GEN_7828; // @[decode.scala 489:11 624:39]
  wire [126:0] _GEN_7851 = _T_258 ? 127'h8000000000101101 : _GEN_7829; // @[decode.scala 624:39 490:8]
  wire [63:0] _GEN_7852 = _T_258 ? medeleg : _GEN_7830; // @[decode.scala 472:28 624:39]
  wire [63:0] _GEN_7853 = _T_258 ? mideleg : _GEN_7831; // @[decode.scala 473:28 624:39]
  wire [63:0] _GEN_7854 = _T_258 ? mie : _GEN_7832; // @[decode.scala 474:28 624:39]
  wire [63:0] _GEN_7855 = _T_258 ? mtvec : _GEN_7833; // @[decode.scala 475:28 624:39]
  wire [63:0] _GEN_7856 = _T_258 ? mcounteren : _GEN_7834; // @[decode.scala 476:28 624:39]
  wire [63:0] _GEN_7857 = _T_258 ? mscratch : _GEN_7835; // @[decode.scala 477:28 624:39]
  wire [63:0] _GEN_7858 = _T_258 ? mepc : _GEN_7836; // @[decode.scala 478:28 624:39]
  wire [63:0] _GEN_7859 = _T_258 ? mcause : _GEN_7837; // @[decode.scala 479:28 624:39]
  wire [63:0] _GEN_7860 = _T_258 ? mtval : _GEN_7838; // @[decode.scala 480:28 624:39]
  wire [63:0] _GEN_7861 = _T_258 ? mip : _GEN_7839; // @[decode.scala 481:28 624:39]
  wire [63:0] _GEN_7862 = _T_258 ? pmpcfg0 : _GEN_7840; // @[decode.scala 482:28 624:39]
  wire [63:0] _GEN_7863 = _T_258 ? pmpaddr0 : _GEN_7841; // @[decode.scala 483:28 624:39]
  wire [63:0] _GEN_7864 = _T_258 ? mvendorid : _GEN_7842; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7865 = _T_258 ? marchid : _GEN_7843; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7866 = _T_258 ? mimpid : _GEN_7844; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7867 = _T_258 ? mhartid : _GEN_7845; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7868 = _T_257 ? csrImmReg : utvec; // @[decode.scala 465:28 624:39 626:38]
  wire [63:0] _GEN_7869 = _T_257 ? uepc : _GEN_7846; // @[decode.scala 466:28 624:39]
  wire [63:0] _GEN_7870 = _T_257 ? ucause : _GEN_7847; // @[decode.scala 467:28 624:39]
  wire [63:0] _GEN_7871 = _T_257 ? scounteren : _GEN_7848; // @[decode.scala 468:28 624:39]
  wire [63:0] _GEN_7872 = _T_257 ? satp : _GEN_7849; // @[decode.scala 469:28 624:39]
  wire [63:0] _GEN_7873 = _T_257 ? _mstatus_T_1 : _GEN_7850; // @[decode.scala 489:11 624:39]
  wire [126:0] _GEN_7874 = _T_257 ? 127'h8000000000101101 : _GEN_7851; // @[decode.scala 624:39 490:8]
  wire [63:0] _GEN_7875 = _T_257 ? medeleg : _GEN_7852; // @[decode.scala 472:28 624:39]
  wire [63:0] _GEN_7876 = _T_257 ? mideleg : _GEN_7853; // @[decode.scala 473:28 624:39]
  wire [63:0] _GEN_7877 = _T_257 ? mie : _GEN_7854; // @[decode.scala 474:28 624:39]
  wire [63:0] _GEN_7878 = _T_257 ? mtvec : _GEN_7855; // @[decode.scala 475:28 624:39]
  wire [63:0] _GEN_7879 = _T_257 ? mcounteren : _GEN_7856; // @[decode.scala 476:28 624:39]
  wire [63:0] _GEN_7880 = _T_257 ? mscratch : _GEN_7857; // @[decode.scala 477:28 624:39]
  wire [63:0] _GEN_7881 = _T_257 ? mepc : _GEN_7858; // @[decode.scala 478:28 624:39]
  wire [63:0] _GEN_7882 = _T_257 ? mcause : _GEN_7859; // @[decode.scala 479:28 624:39]
  wire [63:0] _GEN_7883 = _T_257 ? mtval : _GEN_7860; // @[decode.scala 480:28 624:39]
  wire [63:0] _GEN_7884 = _T_257 ? mip : _GEN_7861; // @[decode.scala 481:28 624:39]
  wire [63:0] _GEN_7885 = _T_257 ? pmpcfg0 : _GEN_7862; // @[decode.scala 482:28 624:39]
  wire [63:0] _GEN_7886 = _T_257 ? pmpaddr0 : _GEN_7863; // @[decode.scala 483:28 624:39]
  wire [63:0] _GEN_7887 = _T_257 ? mvendorid : _GEN_7864; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7888 = _T_257 ? marchid : _GEN_7865; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7889 = _T_257 ? mimpid : _GEN_7866; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7890 = _T_257 ? mhartid : _GEN_7867; // @[decode.scala 487:28 624:39]
  wire [63:0] _GEN_7891 = _T_256 ? csrImmReg : ustatus; // @[decode.scala 464:28 624:39 625:38]
  wire [63:0] _GEN_7892 = _T_256 ? utvec : _GEN_7868; // @[decode.scala 465:28 624:39]
  wire [63:0] _GEN_7893 = _T_256 ? uepc : _GEN_7869; // @[decode.scala 466:28 624:39]
  wire [63:0] _GEN_7894 = _T_256 ? ucause : _GEN_7870; // @[decode.scala 467:28 624:39]
  wire [63:0] _GEN_7895 = _T_256 ? scounteren : _GEN_7871; // @[decode.scala 468:28 624:39]
  wire [63:0] _GEN_7896 = _T_256 ? satp : _GEN_7872; // @[decode.scala 469:28 624:39]
  wire [63:0] _GEN_7897 = _T_256 ? _mstatus_T_1 : _GEN_7873; // @[decode.scala 489:11 624:39]
  wire [126:0] _GEN_7898 = _T_256 ? 127'h8000000000101101 : _GEN_7874; // @[decode.scala 624:39 490:8]
  wire [63:0] _GEN_7899 = _T_256 ? medeleg : _GEN_7875; // @[decode.scala 472:28 624:39]
  wire [63:0] _GEN_7900 = _T_256 ? mideleg : _GEN_7876; // @[decode.scala 473:28 624:39]
  wire [63:0] _GEN_7901 = _T_256 ? mie : _GEN_7877; // @[decode.scala 474:28 624:39]
  wire [63:0] _GEN_7902 = _T_256 ? mtvec : _GEN_7878; // @[decode.scala 475:28 624:39]
  wire [63:0] _GEN_7903 = _T_256 ? mcounteren : _GEN_7879; // @[decode.scala 476:28 624:39]
  wire [63:0] _GEN_7904 = _T_256 ? mscratch : _GEN_7880; // @[decode.scala 477:28 624:39]
  wire [63:0] _GEN_7905 = _T_256 ? mepc : _GEN_7881; // @[decode.scala 478:28 624:39]
  wire [63:0] _GEN_7906 = _T_256 ? mcause : _GEN_7882; // @[decode.scala 479:28 624:39]
  wire [63:0] _GEN_7907 = _T_256 ? mtval : _GEN_7883; // @[decode.scala 480:28 624:39]
  wire [63:0] _GEN_7908 = _T_256 ? mip : _GEN_7884; // @[decode.scala 481:28 624:39]
  wire [63:0] _GEN_7909 = _T_256 ? pmpcfg0 : _GEN_7885; // @[decode.scala 482:28 624:39]
  wire [63:0] _GEN_7910 = _T_256 ? pmpaddr0 : _GEN_7886; // @[decode.scala 483:28 624:39]
  wire [63:0] _GEN_7911 = _T_256 ? mvendorid : _GEN_7887; // @[decode.scala 484:28 624:39]
  wire [63:0] _GEN_7912 = _T_256 ? marchid : _GEN_7888; // @[decode.scala 485:28 624:39]
  wire [63:0] _GEN_7913 = _T_256 ? mimpid : _GEN_7889; // @[decode.scala 486:28 624:39]
  wire [63:0] _GEN_7914 = _T_256 ? mhartid : _GEN_7890; // @[decode.scala 487:28 624:39]
  wire [63:0] _ustatus_T_3 = ustatus | csrImmReg; // @[decode.scala 653:49]
  wire [63:0] _utvec_T_3 = utvec | csrImmReg; // @[decode.scala 654:47]
  wire [63:0] _uepc_T_3 = uepc | csrImmReg; // @[decode.scala 655:46]
  wire [63:0] _ucause_T_3 = ucause | csrImmReg; // @[decode.scala 656:48]
  wire [63:0] _scounteren_T_3 = scounteren | csrImmReg; // @[decode.scala 657:52]
  wire [63:0] _satp_T_3 = satp | csrImmReg; // @[decode.scala 658:46]
  wire [63:0] _mstatus_T_5 = mstatus | csrImmReg; // @[decode.scala 659:49]
  wire [63:0] _misa_T_5 = misa | csrImmReg; // @[decode.scala 660:46]
  wire [63:0] _medeleg_T_3 = medeleg | csrImmReg; // @[decode.scala 661:49]
  wire [63:0] _mideleg_T_3 = mideleg | csrImmReg; // @[decode.scala 662:49]
  wire [63:0] _mie_T_3 = mie | csrImmReg; // @[decode.scala 663:45]
  wire [63:0] _mtvec_T_3 = mtvec | csrImmReg; // @[decode.scala 664:47]
  wire [63:0] _mcounteren_T_3 = mcounteren | csrImmReg; // @[decode.scala 665:52]
  wire [63:0] _mscratch_T_3 = mscratch | csrImmReg; // @[decode.scala 666:50]
  wire [63:0] _mepc_T_3 = mepc | csrImmReg; // @[decode.scala 667:46]
  wire [63:0] _mcause_T_3 = mcause | csrImmReg; // @[decode.scala 668:48]
  wire [63:0] _mtval_T_3 = mtval | csrImmReg; // @[decode.scala 669:47]
  wire [63:0] _mip_T_3 = mip | csrImmReg; // @[decode.scala 670:45]
  wire [63:0] _pmpcfg0_T_3 = pmpcfg0 | csrImmReg; // @[decode.scala 671:49]
  wire [63:0] _pmpaddr0_T_3 = pmpaddr0 | csrImmReg; // @[decode.scala 672:50]
  wire [63:0] _mvendorid_T_3 = mvendorid | csrImmReg; // @[decode.scala 673:51]
  wire [63:0] _marchid_T_3 = marchid | csrImmReg; // @[decode.scala 674:49]
  wire [63:0] _mimpid_T_3 = mimpid | csrImmReg; // @[decode.scala 675:48]
  wire [63:0] _mhartid_T_3 = mhartid | csrImmReg; // @[decode.scala 676:49]
  wire [63:0] _GEN_7915 = _T_279 ? _mhartid_T_3 : mhartid; // @[decode.scala 487:28 652:39 676:38]
  wire [63:0] _GEN_7916 = _T_278 ? _mimpid_T_3 : mimpid; // @[decode.scala 486:28 652:39 675:38]
  wire [63:0] _GEN_7917 = _T_278 ? mhartid : _GEN_7915; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_7918 = _T_277 ? _marchid_T_3 : marchid; // @[decode.scala 485:28 652:39 674:38]
  wire [63:0] _GEN_7919 = _T_277 ? mimpid : _GEN_7916; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_7920 = _T_277 ? mhartid : _GEN_7917; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_7921 = _T_276 ? _mvendorid_T_3 : mvendorid; // @[decode.scala 484:28 652:39 673:38]
  wire [63:0] _GEN_7922 = _T_276 ? marchid : _GEN_7918; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_7923 = _T_276 ? mimpid : _GEN_7919; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_7924 = _T_276 ? mhartid : _GEN_7920; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_7925 = _T_275 ? _pmpaddr0_T_3 : pmpaddr0; // @[decode.scala 483:28 652:39 672:38]
  wire [63:0] _GEN_7926 = _T_275 ? mvendorid : _GEN_7921; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_7927 = _T_275 ? marchid : _GEN_7922; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_7928 = _T_275 ? mimpid : _GEN_7923; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_7929 = _T_275 ? mhartid : _GEN_7924; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_7930 = _T_274 ? _pmpcfg0_T_3 : pmpcfg0; // @[decode.scala 482:28 652:39 671:38]
  wire [63:0] _GEN_7931 = _T_274 ? pmpaddr0 : _GEN_7925; // @[decode.scala 483:28 652:39]
  wire [63:0] _GEN_7932 = _T_274 ? mvendorid : _GEN_7926; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_7933 = _T_274 ? marchid : _GEN_7927; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_7934 = _T_274 ? mimpid : _GEN_7928; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_7935 = _T_274 ? mhartid : _GEN_7929; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_7936 = _T_273 ? _mip_T_3 : mip; // @[decode.scala 481:28 652:39 670:38]
  wire [63:0] _GEN_7937 = _T_273 ? pmpcfg0 : _GEN_7930; // @[decode.scala 482:28 652:39]
  wire [63:0] _GEN_7938 = _T_273 ? pmpaddr0 : _GEN_7931; // @[decode.scala 483:28 652:39]
  wire [63:0] _GEN_7939 = _T_273 ? mvendorid : _GEN_7932; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_7940 = _T_273 ? marchid : _GEN_7933; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_7941 = _T_273 ? mimpid : _GEN_7934; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_7942 = _T_273 ? mhartid : _GEN_7935; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_7943 = _T_272 ? _mtval_T_3 : mtval; // @[decode.scala 480:28 652:39 669:38]
  wire [63:0] _GEN_7944 = _T_272 ? mip : _GEN_7936; // @[decode.scala 481:28 652:39]
  wire [63:0] _GEN_7945 = _T_272 ? pmpcfg0 : _GEN_7937; // @[decode.scala 482:28 652:39]
  wire [63:0] _GEN_7946 = _T_272 ? pmpaddr0 : _GEN_7938; // @[decode.scala 483:28 652:39]
  wire [63:0] _GEN_7947 = _T_272 ? mvendorid : _GEN_7939; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_7948 = _T_272 ? marchid : _GEN_7940; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_7949 = _T_272 ? mimpid : _GEN_7941; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_7950 = _T_272 ? mhartid : _GEN_7942; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_7951 = _T_271 ? _mcause_T_3 : mcause; // @[decode.scala 479:28 652:39 668:38]
  wire [63:0] _GEN_7952 = _T_271 ? mtval : _GEN_7943; // @[decode.scala 480:28 652:39]
  wire [63:0] _GEN_7953 = _T_271 ? mip : _GEN_7944; // @[decode.scala 481:28 652:39]
  wire [63:0] _GEN_7954 = _T_271 ? pmpcfg0 : _GEN_7945; // @[decode.scala 482:28 652:39]
  wire [63:0] _GEN_7955 = _T_271 ? pmpaddr0 : _GEN_7946; // @[decode.scala 483:28 652:39]
  wire [63:0] _GEN_7956 = _T_271 ? mvendorid : _GEN_7947; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_7957 = _T_271 ? marchid : _GEN_7948; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_7958 = _T_271 ? mimpid : _GEN_7949; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_7959 = _T_271 ? mhartid : _GEN_7950; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_7960 = _T_270 ? _mepc_T_3 : mepc; // @[decode.scala 478:28 652:39 667:38]
  wire [63:0] _GEN_7961 = _T_270 ? mcause : _GEN_7951; // @[decode.scala 479:28 652:39]
  wire [63:0] _GEN_7962 = _T_270 ? mtval : _GEN_7952; // @[decode.scala 480:28 652:39]
  wire [63:0] _GEN_7963 = _T_270 ? mip : _GEN_7953; // @[decode.scala 481:28 652:39]
  wire [63:0] _GEN_7964 = _T_270 ? pmpcfg0 : _GEN_7954; // @[decode.scala 482:28 652:39]
  wire [63:0] _GEN_7965 = _T_270 ? pmpaddr0 : _GEN_7955; // @[decode.scala 483:28 652:39]
  wire [63:0] _GEN_7966 = _T_270 ? mvendorid : _GEN_7956; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_7967 = _T_270 ? marchid : _GEN_7957; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_7968 = _T_270 ? mimpid : _GEN_7958; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_7969 = _T_270 ? mhartid : _GEN_7959; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_7970 = _T_269 ? _mscratch_T_3 : mscratch; // @[decode.scala 477:28 652:39 666:38]
  wire [63:0] _GEN_7971 = _T_269 ? mepc : _GEN_7960; // @[decode.scala 478:28 652:39]
  wire [63:0] _GEN_7972 = _T_269 ? mcause : _GEN_7961; // @[decode.scala 479:28 652:39]
  wire [63:0] _GEN_7973 = _T_269 ? mtval : _GEN_7962; // @[decode.scala 480:28 652:39]
  wire [63:0] _GEN_7974 = _T_269 ? mip : _GEN_7963; // @[decode.scala 481:28 652:39]
  wire [63:0] _GEN_7975 = _T_269 ? pmpcfg0 : _GEN_7964; // @[decode.scala 482:28 652:39]
  wire [63:0] _GEN_7976 = _T_269 ? pmpaddr0 : _GEN_7965; // @[decode.scala 483:28 652:39]
  wire [63:0] _GEN_7977 = _T_269 ? mvendorid : _GEN_7966; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_7978 = _T_269 ? marchid : _GEN_7967; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_7979 = _T_269 ? mimpid : _GEN_7968; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_7980 = _T_269 ? mhartid : _GEN_7969; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_7981 = _T_268 ? _mcounteren_T_3 : mcounteren; // @[decode.scala 476:28 652:39 665:38]
  wire [63:0] _GEN_7982 = _T_268 ? mscratch : _GEN_7970; // @[decode.scala 477:28 652:39]
  wire [63:0] _GEN_7983 = _T_268 ? mepc : _GEN_7971; // @[decode.scala 478:28 652:39]
  wire [63:0] _GEN_7984 = _T_268 ? mcause : _GEN_7972; // @[decode.scala 479:28 652:39]
  wire [63:0] _GEN_7985 = _T_268 ? mtval : _GEN_7973; // @[decode.scala 480:28 652:39]
  wire [63:0] _GEN_7986 = _T_268 ? mip : _GEN_7974; // @[decode.scala 481:28 652:39]
  wire [63:0] _GEN_7987 = _T_268 ? pmpcfg0 : _GEN_7975; // @[decode.scala 482:28 652:39]
  wire [63:0] _GEN_7988 = _T_268 ? pmpaddr0 : _GEN_7976; // @[decode.scala 483:28 652:39]
  wire [63:0] _GEN_7989 = _T_268 ? mvendorid : _GEN_7977; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_7990 = _T_268 ? marchid : _GEN_7978; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_7991 = _T_268 ? mimpid : _GEN_7979; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_7992 = _T_268 ? mhartid : _GEN_7980; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_7993 = _T_267 ? _mtvec_T_3 : mtvec; // @[decode.scala 475:28 652:39 664:38]
  wire [63:0] _GEN_7994 = _T_267 ? mcounteren : _GEN_7981; // @[decode.scala 476:28 652:39]
  wire [63:0] _GEN_7995 = _T_267 ? mscratch : _GEN_7982; // @[decode.scala 477:28 652:39]
  wire [63:0] _GEN_7996 = _T_267 ? mepc : _GEN_7983; // @[decode.scala 478:28 652:39]
  wire [63:0] _GEN_7997 = _T_267 ? mcause : _GEN_7984; // @[decode.scala 479:28 652:39]
  wire [63:0] _GEN_7998 = _T_267 ? mtval : _GEN_7985; // @[decode.scala 480:28 652:39]
  wire [63:0] _GEN_7999 = _T_267 ? mip : _GEN_7986; // @[decode.scala 481:28 652:39]
  wire [63:0] _GEN_8000 = _T_267 ? pmpcfg0 : _GEN_7987; // @[decode.scala 482:28 652:39]
  wire [63:0] _GEN_8001 = _T_267 ? pmpaddr0 : _GEN_7988; // @[decode.scala 483:28 652:39]
  wire [63:0] _GEN_8002 = _T_267 ? mvendorid : _GEN_7989; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_8003 = _T_267 ? marchid : _GEN_7990; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_8004 = _T_267 ? mimpid : _GEN_7991; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_8005 = _T_267 ? mhartid : _GEN_7992; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_8006 = _T_266 ? _mie_T_3 : mie; // @[decode.scala 474:28 652:39 663:38]
  wire [63:0] _GEN_8007 = _T_266 ? mtvec : _GEN_7993; // @[decode.scala 475:28 652:39]
  wire [63:0] _GEN_8008 = _T_266 ? mcounteren : _GEN_7994; // @[decode.scala 476:28 652:39]
  wire [63:0] _GEN_8009 = _T_266 ? mscratch : _GEN_7995; // @[decode.scala 477:28 652:39]
  wire [63:0] _GEN_8010 = _T_266 ? mepc : _GEN_7996; // @[decode.scala 478:28 652:39]
  wire [63:0] _GEN_8011 = _T_266 ? mcause : _GEN_7997; // @[decode.scala 479:28 652:39]
  wire [63:0] _GEN_8012 = _T_266 ? mtval : _GEN_7998; // @[decode.scala 480:28 652:39]
  wire [63:0] _GEN_8013 = _T_266 ? mip : _GEN_7999; // @[decode.scala 481:28 652:39]
  wire [63:0] _GEN_8014 = _T_266 ? pmpcfg0 : _GEN_8000; // @[decode.scala 482:28 652:39]
  wire [63:0] _GEN_8015 = _T_266 ? pmpaddr0 : _GEN_8001; // @[decode.scala 483:28 652:39]
  wire [63:0] _GEN_8016 = _T_266 ? mvendorid : _GEN_8002; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_8017 = _T_266 ? marchid : _GEN_8003; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_8018 = _T_266 ? mimpid : _GEN_8004; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_8019 = _T_266 ? mhartid : _GEN_8005; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_8020 = _T_265 ? _mideleg_T_3 : mideleg; // @[decode.scala 473:28 652:39 662:38]
  wire [63:0] _GEN_8021 = _T_265 ? mie : _GEN_8006; // @[decode.scala 474:28 652:39]
  wire [63:0] _GEN_8022 = _T_265 ? mtvec : _GEN_8007; // @[decode.scala 475:28 652:39]
  wire [63:0] _GEN_8023 = _T_265 ? mcounteren : _GEN_8008; // @[decode.scala 476:28 652:39]
  wire [63:0] _GEN_8024 = _T_265 ? mscratch : _GEN_8009; // @[decode.scala 477:28 652:39]
  wire [63:0] _GEN_8025 = _T_265 ? mepc : _GEN_8010; // @[decode.scala 478:28 652:39]
  wire [63:0] _GEN_8026 = _T_265 ? mcause : _GEN_8011; // @[decode.scala 479:28 652:39]
  wire [63:0] _GEN_8027 = _T_265 ? mtval : _GEN_8012; // @[decode.scala 480:28 652:39]
  wire [63:0] _GEN_8028 = _T_265 ? mip : _GEN_8013; // @[decode.scala 481:28 652:39]
  wire [63:0] _GEN_8029 = _T_265 ? pmpcfg0 : _GEN_8014; // @[decode.scala 482:28 652:39]
  wire [63:0] _GEN_8030 = _T_265 ? pmpaddr0 : _GEN_8015; // @[decode.scala 483:28 652:39]
  wire [63:0] _GEN_8031 = _T_265 ? mvendorid : _GEN_8016; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_8032 = _T_265 ? marchid : _GEN_8017; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_8033 = _T_265 ? mimpid : _GEN_8018; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_8034 = _T_265 ? mhartid : _GEN_8019; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_8035 = _T_264 ? _medeleg_T_3 : medeleg; // @[decode.scala 472:28 652:39 661:38]
  wire [63:0] _GEN_8036 = _T_264 ? mideleg : _GEN_8020; // @[decode.scala 473:28 652:39]
  wire [63:0] _GEN_8037 = _T_264 ? mie : _GEN_8021; // @[decode.scala 474:28 652:39]
  wire [63:0] _GEN_8038 = _T_264 ? mtvec : _GEN_8022; // @[decode.scala 475:28 652:39]
  wire [63:0] _GEN_8039 = _T_264 ? mcounteren : _GEN_8023; // @[decode.scala 476:28 652:39]
  wire [63:0] _GEN_8040 = _T_264 ? mscratch : _GEN_8024; // @[decode.scala 477:28 652:39]
  wire [63:0] _GEN_8041 = _T_264 ? mepc : _GEN_8025; // @[decode.scala 478:28 652:39]
  wire [63:0] _GEN_8042 = _T_264 ? mcause : _GEN_8026; // @[decode.scala 479:28 652:39]
  wire [63:0] _GEN_8043 = _T_264 ? mtval : _GEN_8027; // @[decode.scala 480:28 652:39]
  wire [63:0] _GEN_8044 = _T_264 ? mip : _GEN_8028; // @[decode.scala 481:28 652:39]
  wire [63:0] _GEN_8045 = _T_264 ? pmpcfg0 : _GEN_8029; // @[decode.scala 482:28 652:39]
  wire [63:0] _GEN_8046 = _T_264 ? pmpaddr0 : _GEN_8030; // @[decode.scala 483:28 652:39]
  wire [63:0] _GEN_8047 = _T_264 ? mvendorid : _GEN_8031; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_8048 = _T_264 ? marchid : _GEN_8032; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_8049 = _T_264 ? mimpid : _GEN_8033; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_8050 = _T_264 ? mhartid : _GEN_8034; // @[decode.scala 487:28 652:39]
  wire [126:0] _GEN_8051 = _T_263 ? {{63'd0}, _misa_T_5} : 127'h8000000000101101; // @[decode.scala 652:39 660:38 490:8]
  wire [63:0] _GEN_8052 = _T_263 ? medeleg : _GEN_8035; // @[decode.scala 472:28 652:39]
  wire [63:0] _GEN_8053 = _T_263 ? mideleg : _GEN_8036; // @[decode.scala 473:28 652:39]
  wire [63:0] _GEN_8054 = _T_263 ? mie : _GEN_8037; // @[decode.scala 474:28 652:39]
  wire [63:0] _GEN_8055 = _T_263 ? mtvec : _GEN_8038; // @[decode.scala 475:28 652:39]
  wire [63:0] _GEN_8056 = _T_263 ? mcounteren : _GEN_8039; // @[decode.scala 476:28 652:39]
  wire [63:0] _GEN_8057 = _T_263 ? mscratch : _GEN_8040; // @[decode.scala 477:28 652:39]
  wire [63:0] _GEN_8058 = _T_263 ? mepc : _GEN_8041; // @[decode.scala 478:28 652:39]
  wire [63:0] _GEN_8059 = _T_263 ? mcause : _GEN_8042; // @[decode.scala 479:28 652:39]
  wire [63:0] _GEN_8060 = _T_263 ? mtval : _GEN_8043; // @[decode.scala 480:28 652:39]
  wire [63:0] _GEN_8061 = _T_263 ? mip : _GEN_8044; // @[decode.scala 481:28 652:39]
  wire [63:0] _GEN_8062 = _T_263 ? pmpcfg0 : _GEN_8045; // @[decode.scala 482:28 652:39]
  wire [63:0] _GEN_8063 = _T_263 ? pmpaddr0 : _GEN_8046; // @[decode.scala 483:28 652:39]
  wire [63:0] _GEN_8064 = _T_263 ? mvendorid : _GEN_8047; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_8065 = _T_263 ? marchid : _GEN_8048; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_8066 = _T_263 ? mimpid : _GEN_8049; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_8067 = _T_263 ? mhartid : _GEN_8050; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_8068 = _T_262 ? _mstatus_T_5 : _mstatus_T_1; // @[decode.scala 489:11 652:39 659:38]
  wire [126:0] _GEN_8069 = _T_262 ? 127'h8000000000101101 : _GEN_8051; // @[decode.scala 652:39 490:8]
  wire [63:0] _GEN_8070 = _T_262 ? medeleg : _GEN_8052; // @[decode.scala 472:28 652:39]
  wire [63:0] _GEN_8071 = _T_262 ? mideleg : _GEN_8053; // @[decode.scala 473:28 652:39]
  wire [63:0] _GEN_8072 = _T_262 ? mie : _GEN_8054; // @[decode.scala 474:28 652:39]
  wire [63:0] _GEN_8073 = _T_262 ? mtvec : _GEN_8055; // @[decode.scala 475:28 652:39]
  wire [63:0] _GEN_8074 = _T_262 ? mcounteren : _GEN_8056; // @[decode.scala 476:28 652:39]
  wire [63:0] _GEN_8075 = _T_262 ? mscratch : _GEN_8057; // @[decode.scala 477:28 652:39]
  wire [63:0] _GEN_8076 = _T_262 ? mepc : _GEN_8058; // @[decode.scala 478:28 652:39]
  wire [63:0] _GEN_8077 = _T_262 ? mcause : _GEN_8059; // @[decode.scala 479:28 652:39]
  wire [63:0] _GEN_8078 = _T_262 ? mtval : _GEN_8060; // @[decode.scala 480:28 652:39]
  wire [63:0] _GEN_8079 = _T_262 ? mip : _GEN_8061; // @[decode.scala 481:28 652:39]
  wire [63:0] _GEN_8080 = _T_262 ? pmpcfg0 : _GEN_8062; // @[decode.scala 482:28 652:39]
  wire [63:0] _GEN_8081 = _T_262 ? pmpaddr0 : _GEN_8063; // @[decode.scala 483:28 652:39]
  wire [63:0] _GEN_8082 = _T_262 ? mvendorid : _GEN_8064; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_8083 = _T_262 ? marchid : _GEN_8065; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_8084 = _T_262 ? mimpid : _GEN_8066; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_8085 = _T_262 ? mhartid : _GEN_8067; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_8086 = _T_261 ? _satp_T_3 : satp; // @[decode.scala 469:28 652:39 658:38]
  wire [63:0] _GEN_8087 = _T_261 ? _mstatus_T_1 : _GEN_8068; // @[decode.scala 489:11 652:39]
  wire [126:0] _GEN_8088 = _T_261 ? 127'h8000000000101101 : _GEN_8069; // @[decode.scala 652:39 490:8]
  wire [63:0] _GEN_8089 = _T_261 ? medeleg : _GEN_8070; // @[decode.scala 472:28 652:39]
  wire [63:0] _GEN_8090 = _T_261 ? mideleg : _GEN_8071; // @[decode.scala 473:28 652:39]
  wire [63:0] _GEN_8091 = _T_261 ? mie : _GEN_8072; // @[decode.scala 474:28 652:39]
  wire [63:0] _GEN_8092 = _T_261 ? mtvec : _GEN_8073; // @[decode.scala 475:28 652:39]
  wire [63:0] _GEN_8093 = _T_261 ? mcounteren : _GEN_8074; // @[decode.scala 476:28 652:39]
  wire [63:0] _GEN_8094 = _T_261 ? mscratch : _GEN_8075; // @[decode.scala 477:28 652:39]
  wire [63:0] _GEN_8095 = _T_261 ? mepc : _GEN_8076; // @[decode.scala 478:28 652:39]
  wire [63:0] _GEN_8096 = _T_261 ? mcause : _GEN_8077; // @[decode.scala 479:28 652:39]
  wire [63:0] _GEN_8097 = _T_261 ? mtval : _GEN_8078; // @[decode.scala 480:28 652:39]
  wire [63:0] _GEN_8098 = _T_261 ? mip : _GEN_8079; // @[decode.scala 481:28 652:39]
  wire [63:0] _GEN_8099 = _T_261 ? pmpcfg0 : _GEN_8080; // @[decode.scala 482:28 652:39]
  wire [63:0] _GEN_8100 = _T_261 ? pmpaddr0 : _GEN_8081; // @[decode.scala 483:28 652:39]
  wire [63:0] _GEN_8101 = _T_261 ? mvendorid : _GEN_8082; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_8102 = _T_261 ? marchid : _GEN_8083; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_8103 = _T_261 ? mimpid : _GEN_8084; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_8104 = _T_261 ? mhartid : _GEN_8085; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_8105 = _T_260 ? _scounteren_T_3 : scounteren; // @[decode.scala 468:28 652:39 657:38]
  wire [63:0] _GEN_8106 = _T_260 ? satp : _GEN_8086; // @[decode.scala 469:28 652:39]
  wire [63:0] _GEN_8107 = _T_260 ? _mstatus_T_1 : _GEN_8087; // @[decode.scala 489:11 652:39]
  wire [126:0] _GEN_8108 = _T_260 ? 127'h8000000000101101 : _GEN_8088; // @[decode.scala 652:39 490:8]
  wire [63:0] _GEN_8109 = _T_260 ? medeleg : _GEN_8089; // @[decode.scala 472:28 652:39]
  wire [63:0] _GEN_8110 = _T_260 ? mideleg : _GEN_8090; // @[decode.scala 473:28 652:39]
  wire [63:0] _GEN_8111 = _T_260 ? mie : _GEN_8091; // @[decode.scala 474:28 652:39]
  wire [63:0] _GEN_8112 = _T_260 ? mtvec : _GEN_8092; // @[decode.scala 475:28 652:39]
  wire [63:0] _GEN_8113 = _T_260 ? mcounteren : _GEN_8093; // @[decode.scala 476:28 652:39]
  wire [63:0] _GEN_8114 = _T_260 ? mscratch : _GEN_8094; // @[decode.scala 477:28 652:39]
  wire [63:0] _GEN_8115 = _T_260 ? mepc : _GEN_8095; // @[decode.scala 478:28 652:39]
  wire [63:0] _GEN_8116 = _T_260 ? mcause : _GEN_8096; // @[decode.scala 479:28 652:39]
  wire [63:0] _GEN_8117 = _T_260 ? mtval : _GEN_8097; // @[decode.scala 480:28 652:39]
  wire [63:0] _GEN_8118 = _T_260 ? mip : _GEN_8098; // @[decode.scala 481:28 652:39]
  wire [63:0] _GEN_8119 = _T_260 ? pmpcfg0 : _GEN_8099; // @[decode.scala 482:28 652:39]
  wire [63:0] _GEN_8120 = _T_260 ? pmpaddr0 : _GEN_8100; // @[decode.scala 483:28 652:39]
  wire [63:0] _GEN_8121 = _T_260 ? mvendorid : _GEN_8101; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_8122 = _T_260 ? marchid : _GEN_8102; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_8123 = _T_260 ? mimpid : _GEN_8103; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_8124 = _T_260 ? mhartid : _GEN_8104; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_8125 = _T_259 ? _ucause_T_3 : ucause; // @[decode.scala 467:28 652:39 656:38]
  wire [63:0] _GEN_8126 = _T_259 ? scounteren : _GEN_8105; // @[decode.scala 468:28 652:39]
  wire [63:0] _GEN_8127 = _T_259 ? satp : _GEN_8106; // @[decode.scala 469:28 652:39]
  wire [63:0] _GEN_8128 = _T_259 ? _mstatus_T_1 : _GEN_8107; // @[decode.scala 489:11 652:39]
  wire [126:0] _GEN_8129 = _T_259 ? 127'h8000000000101101 : _GEN_8108; // @[decode.scala 652:39 490:8]
  wire [63:0] _GEN_8130 = _T_259 ? medeleg : _GEN_8109; // @[decode.scala 472:28 652:39]
  wire [63:0] _GEN_8131 = _T_259 ? mideleg : _GEN_8110; // @[decode.scala 473:28 652:39]
  wire [63:0] _GEN_8132 = _T_259 ? mie : _GEN_8111; // @[decode.scala 474:28 652:39]
  wire [63:0] _GEN_8133 = _T_259 ? mtvec : _GEN_8112; // @[decode.scala 475:28 652:39]
  wire [63:0] _GEN_8134 = _T_259 ? mcounteren : _GEN_8113; // @[decode.scala 476:28 652:39]
  wire [63:0] _GEN_8135 = _T_259 ? mscratch : _GEN_8114; // @[decode.scala 477:28 652:39]
  wire [63:0] _GEN_8136 = _T_259 ? mepc : _GEN_8115; // @[decode.scala 478:28 652:39]
  wire [63:0] _GEN_8137 = _T_259 ? mcause : _GEN_8116; // @[decode.scala 479:28 652:39]
  wire [63:0] _GEN_8138 = _T_259 ? mtval : _GEN_8117; // @[decode.scala 480:28 652:39]
  wire [63:0] _GEN_8139 = _T_259 ? mip : _GEN_8118; // @[decode.scala 481:28 652:39]
  wire [63:0] _GEN_8140 = _T_259 ? pmpcfg0 : _GEN_8119; // @[decode.scala 482:28 652:39]
  wire [63:0] _GEN_8141 = _T_259 ? pmpaddr0 : _GEN_8120; // @[decode.scala 483:28 652:39]
  wire [63:0] _GEN_8142 = _T_259 ? mvendorid : _GEN_8121; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_8143 = _T_259 ? marchid : _GEN_8122; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_8144 = _T_259 ? mimpid : _GEN_8123; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_8145 = _T_259 ? mhartid : _GEN_8124; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_8146 = _T_258 ? _uepc_T_3 : uepc; // @[decode.scala 466:28 652:39 655:38]
  wire [63:0] _GEN_8147 = _T_258 ? ucause : _GEN_8125; // @[decode.scala 467:28 652:39]
  wire [63:0] _GEN_8148 = _T_258 ? scounteren : _GEN_8126; // @[decode.scala 468:28 652:39]
  wire [63:0] _GEN_8149 = _T_258 ? satp : _GEN_8127; // @[decode.scala 469:28 652:39]
  wire [63:0] _GEN_8150 = _T_258 ? _mstatus_T_1 : _GEN_8128; // @[decode.scala 489:11 652:39]
  wire [126:0] _GEN_8151 = _T_258 ? 127'h8000000000101101 : _GEN_8129; // @[decode.scala 652:39 490:8]
  wire [63:0] _GEN_8152 = _T_258 ? medeleg : _GEN_8130; // @[decode.scala 472:28 652:39]
  wire [63:0] _GEN_8153 = _T_258 ? mideleg : _GEN_8131; // @[decode.scala 473:28 652:39]
  wire [63:0] _GEN_8154 = _T_258 ? mie : _GEN_8132; // @[decode.scala 474:28 652:39]
  wire [63:0] _GEN_8155 = _T_258 ? mtvec : _GEN_8133; // @[decode.scala 475:28 652:39]
  wire [63:0] _GEN_8156 = _T_258 ? mcounteren : _GEN_8134; // @[decode.scala 476:28 652:39]
  wire [63:0] _GEN_8157 = _T_258 ? mscratch : _GEN_8135; // @[decode.scala 477:28 652:39]
  wire [63:0] _GEN_8158 = _T_258 ? mepc : _GEN_8136; // @[decode.scala 478:28 652:39]
  wire [63:0] _GEN_8159 = _T_258 ? mcause : _GEN_8137; // @[decode.scala 479:28 652:39]
  wire [63:0] _GEN_8160 = _T_258 ? mtval : _GEN_8138; // @[decode.scala 480:28 652:39]
  wire [63:0] _GEN_8161 = _T_258 ? mip : _GEN_8139; // @[decode.scala 481:28 652:39]
  wire [63:0] _GEN_8162 = _T_258 ? pmpcfg0 : _GEN_8140; // @[decode.scala 482:28 652:39]
  wire [63:0] _GEN_8163 = _T_258 ? pmpaddr0 : _GEN_8141; // @[decode.scala 483:28 652:39]
  wire [63:0] _GEN_8164 = _T_258 ? mvendorid : _GEN_8142; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_8165 = _T_258 ? marchid : _GEN_8143; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_8166 = _T_258 ? mimpid : _GEN_8144; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_8167 = _T_258 ? mhartid : _GEN_8145; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_8168 = _T_257 ? _utvec_T_3 : utvec; // @[decode.scala 465:28 652:39 654:38]
  wire [63:0] _GEN_8169 = _T_257 ? uepc : _GEN_8146; // @[decode.scala 466:28 652:39]
  wire [63:0] _GEN_8170 = _T_257 ? ucause : _GEN_8147; // @[decode.scala 467:28 652:39]
  wire [63:0] _GEN_8171 = _T_257 ? scounteren : _GEN_8148; // @[decode.scala 468:28 652:39]
  wire [63:0] _GEN_8172 = _T_257 ? satp : _GEN_8149; // @[decode.scala 469:28 652:39]
  wire [63:0] _GEN_8173 = _T_257 ? _mstatus_T_1 : _GEN_8150; // @[decode.scala 489:11 652:39]
  wire [126:0] _GEN_8174 = _T_257 ? 127'h8000000000101101 : _GEN_8151; // @[decode.scala 652:39 490:8]
  wire [63:0] _GEN_8175 = _T_257 ? medeleg : _GEN_8152; // @[decode.scala 472:28 652:39]
  wire [63:0] _GEN_8176 = _T_257 ? mideleg : _GEN_8153; // @[decode.scala 473:28 652:39]
  wire [63:0] _GEN_8177 = _T_257 ? mie : _GEN_8154; // @[decode.scala 474:28 652:39]
  wire [63:0] _GEN_8178 = _T_257 ? mtvec : _GEN_8155; // @[decode.scala 475:28 652:39]
  wire [63:0] _GEN_8179 = _T_257 ? mcounteren : _GEN_8156; // @[decode.scala 476:28 652:39]
  wire [63:0] _GEN_8180 = _T_257 ? mscratch : _GEN_8157; // @[decode.scala 477:28 652:39]
  wire [63:0] _GEN_8181 = _T_257 ? mepc : _GEN_8158; // @[decode.scala 478:28 652:39]
  wire [63:0] _GEN_8182 = _T_257 ? mcause : _GEN_8159; // @[decode.scala 479:28 652:39]
  wire [63:0] _GEN_8183 = _T_257 ? mtval : _GEN_8160; // @[decode.scala 480:28 652:39]
  wire [63:0] _GEN_8184 = _T_257 ? mip : _GEN_8161; // @[decode.scala 481:28 652:39]
  wire [63:0] _GEN_8185 = _T_257 ? pmpcfg0 : _GEN_8162; // @[decode.scala 482:28 652:39]
  wire [63:0] _GEN_8186 = _T_257 ? pmpaddr0 : _GEN_8163; // @[decode.scala 483:28 652:39]
  wire [63:0] _GEN_8187 = _T_257 ? mvendorid : _GEN_8164; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_8188 = _T_257 ? marchid : _GEN_8165; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_8189 = _T_257 ? mimpid : _GEN_8166; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_8190 = _T_257 ? mhartid : _GEN_8167; // @[decode.scala 487:28 652:39]
  wire [63:0] _GEN_8191 = _T_256 ? _ustatus_T_3 : ustatus; // @[decode.scala 464:28 652:39 653:38]
  wire [63:0] _GEN_8192 = _T_256 ? utvec : _GEN_8168; // @[decode.scala 465:28 652:39]
  wire [63:0] _GEN_8193 = _T_256 ? uepc : _GEN_8169; // @[decode.scala 466:28 652:39]
  wire [63:0] _GEN_8194 = _T_256 ? ucause : _GEN_8170; // @[decode.scala 467:28 652:39]
  wire [63:0] _GEN_8195 = _T_256 ? scounteren : _GEN_8171; // @[decode.scala 468:28 652:39]
  wire [63:0] _GEN_8196 = _T_256 ? satp : _GEN_8172; // @[decode.scala 469:28 652:39]
  wire [63:0] _GEN_8197 = _T_256 ? _mstatus_T_1 : _GEN_8173; // @[decode.scala 489:11 652:39]
  wire [126:0] _GEN_8198 = _T_256 ? 127'h8000000000101101 : _GEN_8174; // @[decode.scala 652:39 490:8]
  wire [63:0] _GEN_8199 = _T_256 ? medeleg : _GEN_8175; // @[decode.scala 472:28 652:39]
  wire [63:0] _GEN_8200 = _T_256 ? mideleg : _GEN_8176; // @[decode.scala 473:28 652:39]
  wire [63:0] _GEN_8201 = _T_256 ? mie : _GEN_8177; // @[decode.scala 474:28 652:39]
  wire [63:0] _GEN_8202 = _T_256 ? mtvec : _GEN_8178; // @[decode.scala 475:28 652:39]
  wire [63:0] _GEN_8203 = _T_256 ? mcounteren : _GEN_8179; // @[decode.scala 476:28 652:39]
  wire [63:0] _GEN_8204 = _T_256 ? mscratch : _GEN_8180; // @[decode.scala 477:28 652:39]
  wire [63:0] _GEN_8205 = _T_256 ? mepc : _GEN_8181; // @[decode.scala 478:28 652:39]
  wire [63:0] _GEN_8206 = _T_256 ? mcause : _GEN_8182; // @[decode.scala 479:28 652:39]
  wire [63:0] _GEN_8207 = _T_256 ? mtval : _GEN_8183; // @[decode.scala 480:28 652:39]
  wire [63:0] _GEN_8208 = _T_256 ? mip : _GEN_8184; // @[decode.scala 481:28 652:39]
  wire [63:0] _GEN_8209 = _T_256 ? pmpcfg0 : _GEN_8185; // @[decode.scala 482:28 652:39]
  wire [63:0] _GEN_8210 = _T_256 ? pmpaddr0 : _GEN_8186; // @[decode.scala 483:28 652:39]
  wire [63:0] _GEN_8211 = _T_256 ? mvendorid : _GEN_8187; // @[decode.scala 484:28 652:39]
  wire [63:0] _GEN_8212 = _T_256 ? marchid : _GEN_8188; // @[decode.scala 485:28 652:39]
  wire [63:0] _GEN_8213 = _T_256 ? mimpid : _GEN_8189; // @[decode.scala 486:28 652:39]
  wire [63:0] _GEN_8214 = _T_256 ? mhartid : _GEN_8190; // @[decode.scala 487:28 652:39]
  wire [63:0] _ustatus_T_4 = ~csrImmReg; // @[decode.scala 681:51]
  wire [63:0] _ustatus_T_5 = ustatus & _ustatus_T_4; // @[decode.scala 681:49]
  wire [63:0] _utvec_T_5 = utvec & _ustatus_T_4; // @[decode.scala 682:47]
  wire [63:0] _uepc_T_5 = uepc & _ustatus_T_4; // @[decode.scala 683:46]
  wire [63:0] _ucause_T_5 = ucause & _ustatus_T_4; // @[decode.scala 684:48]
  wire [63:0] _scounteren_T_5 = scounteren & _ustatus_T_4; // @[decode.scala 685:52]
  wire [63:0] _satp_T_5 = satp & _ustatus_T_4; // @[decode.scala 686:46]
  wire [63:0] _mstatus_T_7 = mstatus & _ustatus_T_4; // @[decode.scala 687:49]
  wire [63:0] _misa_T_7 = misa & _ustatus_T_4; // @[decode.scala 688:46]
  wire [63:0] _medeleg_T_5 = medeleg & _ustatus_T_4; // @[decode.scala 689:49]
  wire [63:0] _mideleg_T_5 = mideleg & _ustatus_T_4; // @[decode.scala 690:49]
  wire [63:0] _mie_T_5 = mie & _ustatus_T_4; // @[decode.scala 691:45]
  wire [63:0] _mtvec_T_5 = mtvec & _ustatus_T_4; // @[decode.scala 692:47]
  wire [63:0] _mcounteren_T_5 = mcounteren & _ustatus_T_4; // @[decode.scala 693:52]
  wire [63:0] _mscratch_T_5 = mscratch & _ustatus_T_4; // @[decode.scala 694:50]
  wire [63:0] _mepc_T_5 = mepc & _ustatus_T_4; // @[decode.scala 695:46]
  wire [63:0] _mcause_T_5 = mcause & _ustatus_T_4; // @[decode.scala 696:48]
  wire [63:0] _mtval_T_5 = mtval & _ustatus_T_4; // @[decode.scala 697:47]
  wire [63:0] _mip_T_5 = mip & _ustatus_T_4; // @[decode.scala 698:45]
  wire [63:0] _pmpcfg0_T_5 = pmpcfg0 & _ustatus_T_4; // @[decode.scala 699:49]
  wire [63:0] _pmpaddr0_T_5 = pmpaddr0 & _ustatus_T_4; // @[decode.scala 700:50]
  wire [63:0] _mvendorid_T_5 = mvendorid & _ustatus_T_4; // @[decode.scala 701:51]
  wire [63:0] _marchid_T_5 = marchid & _ustatus_T_4; // @[decode.scala 702:49]
  wire [63:0] _mimpid_T_5 = mimpid & _ustatus_T_4; // @[decode.scala 703:48]
  wire [63:0] _mhartid_T_5 = mhartid & _ustatus_T_4; // @[decode.scala 704:49]
  wire [63:0] _GEN_8215 = _T_279 ? _mhartid_T_5 : mhartid; // @[decode.scala 487:28 680:39 704:38]
  wire [63:0] _GEN_8216 = _T_278 ? _mimpid_T_5 : mimpid; // @[decode.scala 486:28 680:39 703:38]
  wire [63:0] _GEN_8217 = _T_278 ? mhartid : _GEN_8215; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8218 = _T_277 ? _marchid_T_5 : marchid; // @[decode.scala 485:28 680:39 702:38]
  wire [63:0] _GEN_8219 = _T_277 ? mimpid : _GEN_8216; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8220 = _T_277 ? mhartid : _GEN_8217; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8221 = _T_276 ? _mvendorid_T_5 : mvendorid; // @[decode.scala 484:28 680:39 701:38]
  wire [63:0] _GEN_8222 = _T_276 ? marchid : _GEN_8218; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8223 = _T_276 ? mimpid : _GEN_8219; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8224 = _T_276 ? mhartid : _GEN_8220; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8225 = _T_275 ? _pmpaddr0_T_5 : pmpaddr0; // @[decode.scala 483:28 680:39 700:38]
  wire [63:0] _GEN_8226 = _T_275 ? mvendorid : _GEN_8221; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8227 = _T_275 ? marchid : _GEN_8222; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8228 = _T_275 ? mimpid : _GEN_8223; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8229 = _T_275 ? mhartid : _GEN_8224; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8230 = _T_274 ? _pmpcfg0_T_5 : pmpcfg0; // @[decode.scala 482:28 680:39 699:38]
  wire [63:0] _GEN_8231 = _T_274 ? pmpaddr0 : _GEN_8225; // @[decode.scala 483:28 680:39]
  wire [63:0] _GEN_8232 = _T_274 ? mvendorid : _GEN_8226; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8233 = _T_274 ? marchid : _GEN_8227; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8234 = _T_274 ? mimpid : _GEN_8228; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8235 = _T_274 ? mhartid : _GEN_8229; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8236 = _T_273 ? _mip_T_5 : mip; // @[decode.scala 481:28 680:39 698:38]
  wire [63:0] _GEN_8237 = _T_273 ? pmpcfg0 : _GEN_8230; // @[decode.scala 482:28 680:39]
  wire [63:0] _GEN_8238 = _T_273 ? pmpaddr0 : _GEN_8231; // @[decode.scala 483:28 680:39]
  wire [63:0] _GEN_8239 = _T_273 ? mvendorid : _GEN_8232; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8240 = _T_273 ? marchid : _GEN_8233; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8241 = _T_273 ? mimpid : _GEN_8234; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8242 = _T_273 ? mhartid : _GEN_8235; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8243 = _T_272 ? _mtval_T_5 : mtval; // @[decode.scala 480:28 680:39 697:38]
  wire [63:0] _GEN_8244 = _T_272 ? mip : _GEN_8236; // @[decode.scala 481:28 680:39]
  wire [63:0] _GEN_8245 = _T_272 ? pmpcfg0 : _GEN_8237; // @[decode.scala 482:28 680:39]
  wire [63:0] _GEN_8246 = _T_272 ? pmpaddr0 : _GEN_8238; // @[decode.scala 483:28 680:39]
  wire [63:0] _GEN_8247 = _T_272 ? mvendorid : _GEN_8239; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8248 = _T_272 ? marchid : _GEN_8240; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8249 = _T_272 ? mimpid : _GEN_8241; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8250 = _T_272 ? mhartid : _GEN_8242; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8251 = _T_271 ? _mcause_T_5 : mcause; // @[decode.scala 479:28 680:39 696:38]
  wire [63:0] _GEN_8252 = _T_271 ? mtval : _GEN_8243; // @[decode.scala 480:28 680:39]
  wire [63:0] _GEN_8253 = _T_271 ? mip : _GEN_8244; // @[decode.scala 481:28 680:39]
  wire [63:0] _GEN_8254 = _T_271 ? pmpcfg0 : _GEN_8245; // @[decode.scala 482:28 680:39]
  wire [63:0] _GEN_8255 = _T_271 ? pmpaddr0 : _GEN_8246; // @[decode.scala 483:28 680:39]
  wire [63:0] _GEN_8256 = _T_271 ? mvendorid : _GEN_8247; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8257 = _T_271 ? marchid : _GEN_8248; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8258 = _T_271 ? mimpid : _GEN_8249; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8259 = _T_271 ? mhartid : _GEN_8250; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8260 = _T_270 ? _mepc_T_5 : mepc; // @[decode.scala 478:28 680:39 695:38]
  wire [63:0] _GEN_8261 = _T_270 ? mcause : _GEN_8251; // @[decode.scala 479:28 680:39]
  wire [63:0] _GEN_8262 = _T_270 ? mtval : _GEN_8252; // @[decode.scala 480:28 680:39]
  wire [63:0] _GEN_8263 = _T_270 ? mip : _GEN_8253; // @[decode.scala 481:28 680:39]
  wire [63:0] _GEN_8264 = _T_270 ? pmpcfg0 : _GEN_8254; // @[decode.scala 482:28 680:39]
  wire [63:0] _GEN_8265 = _T_270 ? pmpaddr0 : _GEN_8255; // @[decode.scala 483:28 680:39]
  wire [63:0] _GEN_8266 = _T_270 ? mvendorid : _GEN_8256; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8267 = _T_270 ? marchid : _GEN_8257; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8268 = _T_270 ? mimpid : _GEN_8258; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8269 = _T_270 ? mhartid : _GEN_8259; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8270 = _T_269 ? _mscratch_T_5 : mscratch; // @[decode.scala 477:28 680:39 694:38]
  wire [63:0] _GEN_8271 = _T_269 ? mepc : _GEN_8260; // @[decode.scala 478:28 680:39]
  wire [63:0] _GEN_8272 = _T_269 ? mcause : _GEN_8261; // @[decode.scala 479:28 680:39]
  wire [63:0] _GEN_8273 = _T_269 ? mtval : _GEN_8262; // @[decode.scala 480:28 680:39]
  wire [63:0] _GEN_8274 = _T_269 ? mip : _GEN_8263; // @[decode.scala 481:28 680:39]
  wire [63:0] _GEN_8275 = _T_269 ? pmpcfg0 : _GEN_8264; // @[decode.scala 482:28 680:39]
  wire [63:0] _GEN_8276 = _T_269 ? pmpaddr0 : _GEN_8265; // @[decode.scala 483:28 680:39]
  wire [63:0] _GEN_8277 = _T_269 ? mvendorid : _GEN_8266; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8278 = _T_269 ? marchid : _GEN_8267; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8279 = _T_269 ? mimpid : _GEN_8268; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8280 = _T_269 ? mhartid : _GEN_8269; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8281 = _T_268 ? _mcounteren_T_5 : mcounteren; // @[decode.scala 476:28 680:39 693:38]
  wire [63:0] _GEN_8282 = _T_268 ? mscratch : _GEN_8270; // @[decode.scala 477:28 680:39]
  wire [63:0] _GEN_8283 = _T_268 ? mepc : _GEN_8271; // @[decode.scala 478:28 680:39]
  wire [63:0] _GEN_8284 = _T_268 ? mcause : _GEN_8272; // @[decode.scala 479:28 680:39]
  wire [63:0] _GEN_8285 = _T_268 ? mtval : _GEN_8273; // @[decode.scala 480:28 680:39]
  wire [63:0] _GEN_8286 = _T_268 ? mip : _GEN_8274; // @[decode.scala 481:28 680:39]
  wire [63:0] _GEN_8287 = _T_268 ? pmpcfg0 : _GEN_8275; // @[decode.scala 482:28 680:39]
  wire [63:0] _GEN_8288 = _T_268 ? pmpaddr0 : _GEN_8276; // @[decode.scala 483:28 680:39]
  wire [63:0] _GEN_8289 = _T_268 ? mvendorid : _GEN_8277; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8290 = _T_268 ? marchid : _GEN_8278; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8291 = _T_268 ? mimpid : _GEN_8279; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8292 = _T_268 ? mhartid : _GEN_8280; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8293 = _T_267 ? _mtvec_T_5 : mtvec; // @[decode.scala 475:28 680:39 692:38]
  wire [63:0] _GEN_8294 = _T_267 ? mcounteren : _GEN_8281; // @[decode.scala 476:28 680:39]
  wire [63:0] _GEN_8295 = _T_267 ? mscratch : _GEN_8282; // @[decode.scala 477:28 680:39]
  wire [63:0] _GEN_8296 = _T_267 ? mepc : _GEN_8283; // @[decode.scala 478:28 680:39]
  wire [63:0] _GEN_8297 = _T_267 ? mcause : _GEN_8284; // @[decode.scala 479:28 680:39]
  wire [63:0] _GEN_8298 = _T_267 ? mtval : _GEN_8285; // @[decode.scala 480:28 680:39]
  wire [63:0] _GEN_8299 = _T_267 ? mip : _GEN_8286; // @[decode.scala 481:28 680:39]
  wire [63:0] _GEN_8300 = _T_267 ? pmpcfg0 : _GEN_8287; // @[decode.scala 482:28 680:39]
  wire [63:0] _GEN_8301 = _T_267 ? pmpaddr0 : _GEN_8288; // @[decode.scala 483:28 680:39]
  wire [63:0] _GEN_8302 = _T_267 ? mvendorid : _GEN_8289; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8303 = _T_267 ? marchid : _GEN_8290; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8304 = _T_267 ? mimpid : _GEN_8291; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8305 = _T_267 ? mhartid : _GEN_8292; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8306 = _T_266 ? _mie_T_5 : mie; // @[decode.scala 474:28 680:39 691:38]
  wire [63:0] _GEN_8307 = _T_266 ? mtvec : _GEN_8293; // @[decode.scala 475:28 680:39]
  wire [63:0] _GEN_8308 = _T_266 ? mcounteren : _GEN_8294; // @[decode.scala 476:28 680:39]
  wire [63:0] _GEN_8309 = _T_266 ? mscratch : _GEN_8295; // @[decode.scala 477:28 680:39]
  wire [63:0] _GEN_8310 = _T_266 ? mepc : _GEN_8296; // @[decode.scala 478:28 680:39]
  wire [63:0] _GEN_8311 = _T_266 ? mcause : _GEN_8297; // @[decode.scala 479:28 680:39]
  wire [63:0] _GEN_8312 = _T_266 ? mtval : _GEN_8298; // @[decode.scala 480:28 680:39]
  wire [63:0] _GEN_8313 = _T_266 ? mip : _GEN_8299; // @[decode.scala 481:28 680:39]
  wire [63:0] _GEN_8314 = _T_266 ? pmpcfg0 : _GEN_8300; // @[decode.scala 482:28 680:39]
  wire [63:0] _GEN_8315 = _T_266 ? pmpaddr0 : _GEN_8301; // @[decode.scala 483:28 680:39]
  wire [63:0] _GEN_8316 = _T_266 ? mvendorid : _GEN_8302; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8317 = _T_266 ? marchid : _GEN_8303; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8318 = _T_266 ? mimpid : _GEN_8304; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8319 = _T_266 ? mhartid : _GEN_8305; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8320 = _T_265 ? _mideleg_T_5 : mideleg; // @[decode.scala 473:28 680:39 690:38]
  wire [63:0] _GEN_8321 = _T_265 ? mie : _GEN_8306; // @[decode.scala 474:28 680:39]
  wire [63:0] _GEN_8322 = _T_265 ? mtvec : _GEN_8307; // @[decode.scala 475:28 680:39]
  wire [63:0] _GEN_8323 = _T_265 ? mcounteren : _GEN_8308; // @[decode.scala 476:28 680:39]
  wire [63:0] _GEN_8324 = _T_265 ? mscratch : _GEN_8309; // @[decode.scala 477:28 680:39]
  wire [63:0] _GEN_8325 = _T_265 ? mepc : _GEN_8310; // @[decode.scala 478:28 680:39]
  wire [63:0] _GEN_8326 = _T_265 ? mcause : _GEN_8311; // @[decode.scala 479:28 680:39]
  wire [63:0] _GEN_8327 = _T_265 ? mtval : _GEN_8312; // @[decode.scala 480:28 680:39]
  wire [63:0] _GEN_8328 = _T_265 ? mip : _GEN_8313; // @[decode.scala 481:28 680:39]
  wire [63:0] _GEN_8329 = _T_265 ? pmpcfg0 : _GEN_8314; // @[decode.scala 482:28 680:39]
  wire [63:0] _GEN_8330 = _T_265 ? pmpaddr0 : _GEN_8315; // @[decode.scala 483:28 680:39]
  wire [63:0] _GEN_8331 = _T_265 ? mvendorid : _GEN_8316; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8332 = _T_265 ? marchid : _GEN_8317; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8333 = _T_265 ? mimpid : _GEN_8318; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8334 = _T_265 ? mhartid : _GEN_8319; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8335 = _T_264 ? _medeleg_T_5 : medeleg; // @[decode.scala 472:28 680:39 689:38]
  wire [63:0] _GEN_8336 = _T_264 ? mideleg : _GEN_8320; // @[decode.scala 473:28 680:39]
  wire [63:0] _GEN_8337 = _T_264 ? mie : _GEN_8321; // @[decode.scala 474:28 680:39]
  wire [63:0] _GEN_8338 = _T_264 ? mtvec : _GEN_8322; // @[decode.scala 475:28 680:39]
  wire [63:0] _GEN_8339 = _T_264 ? mcounteren : _GEN_8323; // @[decode.scala 476:28 680:39]
  wire [63:0] _GEN_8340 = _T_264 ? mscratch : _GEN_8324; // @[decode.scala 477:28 680:39]
  wire [63:0] _GEN_8341 = _T_264 ? mepc : _GEN_8325; // @[decode.scala 478:28 680:39]
  wire [63:0] _GEN_8342 = _T_264 ? mcause : _GEN_8326; // @[decode.scala 479:28 680:39]
  wire [63:0] _GEN_8343 = _T_264 ? mtval : _GEN_8327; // @[decode.scala 480:28 680:39]
  wire [63:0] _GEN_8344 = _T_264 ? mip : _GEN_8328; // @[decode.scala 481:28 680:39]
  wire [63:0] _GEN_8345 = _T_264 ? pmpcfg0 : _GEN_8329; // @[decode.scala 482:28 680:39]
  wire [63:0] _GEN_8346 = _T_264 ? pmpaddr0 : _GEN_8330; // @[decode.scala 483:28 680:39]
  wire [63:0] _GEN_8347 = _T_264 ? mvendorid : _GEN_8331; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8348 = _T_264 ? marchid : _GEN_8332; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8349 = _T_264 ? mimpid : _GEN_8333; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8350 = _T_264 ? mhartid : _GEN_8334; // @[decode.scala 487:28 680:39]
  wire [126:0] _GEN_8351 = _T_263 ? {{63'd0}, _misa_T_7} : 127'h8000000000101101; // @[decode.scala 680:39 688:38 490:8]
  wire [63:0] _GEN_8352 = _T_263 ? medeleg : _GEN_8335; // @[decode.scala 472:28 680:39]
  wire [63:0] _GEN_8353 = _T_263 ? mideleg : _GEN_8336; // @[decode.scala 473:28 680:39]
  wire [63:0] _GEN_8354 = _T_263 ? mie : _GEN_8337; // @[decode.scala 474:28 680:39]
  wire [63:0] _GEN_8355 = _T_263 ? mtvec : _GEN_8338; // @[decode.scala 475:28 680:39]
  wire [63:0] _GEN_8356 = _T_263 ? mcounteren : _GEN_8339; // @[decode.scala 476:28 680:39]
  wire [63:0] _GEN_8357 = _T_263 ? mscratch : _GEN_8340; // @[decode.scala 477:28 680:39]
  wire [63:0] _GEN_8358 = _T_263 ? mepc : _GEN_8341; // @[decode.scala 478:28 680:39]
  wire [63:0] _GEN_8359 = _T_263 ? mcause : _GEN_8342; // @[decode.scala 479:28 680:39]
  wire [63:0] _GEN_8360 = _T_263 ? mtval : _GEN_8343; // @[decode.scala 480:28 680:39]
  wire [63:0] _GEN_8361 = _T_263 ? mip : _GEN_8344; // @[decode.scala 481:28 680:39]
  wire [63:0] _GEN_8362 = _T_263 ? pmpcfg0 : _GEN_8345; // @[decode.scala 482:28 680:39]
  wire [63:0] _GEN_8363 = _T_263 ? pmpaddr0 : _GEN_8346; // @[decode.scala 483:28 680:39]
  wire [63:0] _GEN_8364 = _T_263 ? mvendorid : _GEN_8347; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8365 = _T_263 ? marchid : _GEN_8348; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8366 = _T_263 ? mimpid : _GEN_8349; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8367 = _T_263 ? mhartid : _GEN_8350; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8368 = _T_262 ? _mstatus_T_7 : _mstatus_T_1; // @[decode.scala 489:11 680:39 687:38]
  wire [126:0] _GEN_8369 = _T_262 ? 127'h8000000000101101 : _GEN_8351; // @[decode.scala 680:39 490:8]
  wire [63:0] _GEN_8370 = _T_262 ? medeleg : _GEN_8352; // @[decode.scala 472:28 680:39]
  wire [63:0] _GEN_8371 = _T_262 ? mideleg : _GEN_8353; // @[decode.scala 473:28 680:39]
  wire [63:0] _GEN_8372 = _T_262 ? mie : _GEN_8354; // @[decode.scala 474:28 680:39]
  wire [63:0] _GEN_8373 = _T_262 ? mtvec : _GEN_8355; // @[decode.scala 475:28 680:39]
  wire [63:0] _GEN_8374 = _T_262 ? mcounteren : _GEN_8356; // @[decode.scala 476:28 680:39]
  wire [63:0] _GEN_8375 = _T_262 ? mscratch : _GEN_8357; // @[decode.scala 477:28 680:39]
  wire [63:0] _GEN_8376 = _T_262 ? mepc : _GEN_8358; // @[decode.scala 478:28 680:39]
  wire [63:0] _GEN_8377 = _T_262 ? mcause : _GEN_8359; // @[decode.scala 479:28 680:39]
  wire [63:0] _GEN_8378 = _T_262 ? mtval : _GEN_8360; // @[decode.scala 480:28 680:39]
  wire [63:0] _GEN_8379 = _T_262 ? mip : _GEN_8361; // @[decode.scala 481:28 680:39]
  wire [63:0] _GEN_8380 = _T_262 ? pmpcfg0 : _GEN_8362; // @[decode.scala 482:28 680:39]
  wire [63:0] _GEN_8381 = _T_262 ? pmpaddr0 : _GEN_8363; // @[decode.scala 483:28 680:39]
  wire [63:0] _GEN_8382 = _T_262 ? mvendorid : _GEN_8364; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8383 = _T_262 ? marchid : _GEN_8365; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8384 = _T_262 ? mimpid : _GEN_8366; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8385 = _T_262 ? mhartid : _GEN_8367; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8386 = _T_261 ? _satp_T_5 : satp; // @[decode.scala 469:28 680:39 686:38]
  wire [63:0] _GEN_8387 = _T_261 ? _mstatus_T_1 : _GEN_8368; // @[decode.scala 489:11 680:39]
  wire [126:0] _GEN_8388 = _T_261 ? 127'h8000000000101101 : _GEN_8369; // @[decode.scala 680:39 490:8]
  wire [63:0] _GEN_8389 = _T_261 ? medeleg : _GEN_8370; // @[decode.scala 472:28 680:39]
  wire [63:0] _GEN_8390 = _T_261 ? mideleg : _GEN_8371; // @[decode.scala 473:28 680:39]
  wire [63:0] _GEN_8391 = _T_261 ? mie : _GEN_8372; // @[decode.scala 474:28 680:39]
  wire [63:0] _GEN_8392 = _T_261 ? mtvec : _GEN_8373; // @[decode.scala 475:28 680:39]
  wire [63:0] _GEN_8393 = _T_261 ? mcounteren : _GEN_8374; // @[decode.scala 476:28 680:39]
  wire [63:0] _GEN_8394 = _T_261 ? mscratch : _GEN_8375; // @[decode.scala 477:28 680:39]
  wire [63:0] _GEN_8395 = _T_261 ? mepc : _GEN_8376; // @[decode.scala 478:28 680:39]
  wire [63:0] _GEN_8396 = _T_261 ? mcause : _GEN_8377; // @[decode.scala 479:28 680:39]
  wire [63:0] _GEN_8397 = _T_261 ? mtval : _GEN_8378; // @[decode.scala 480:28 680:39]
  wire [63:0] _GEN_8398 = _T_261 ? mip : _GEN_8379; // @[decode.scala 481:28 680:39]
  wire [63:0] _GEN_8399 = _T_261 ? pmpcfg0 : _GEN_8380; // @[decode.scala 482:28 680:39]
  wire [63:0] _GEN_8400 = _T_261 ? pmpaddr0 : _GEN_8381; // @[decode.scala 483:28 680:39]
  wire [63:0] _GEN_8401 = _T_261 ? mvendorid : _GEN_8382; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8402 = _T_261 ? marchid : _GEN_8383; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8403 = _T_261 ? mimpid : _GEN_8384; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8404 = _T_261 ? mhartid : _GEN_8385; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8405 = _T_260 ? _scounteren_T_5 : scounteren; // @[decode.scala 468:28 680:39 685:38]
  wire [63:0] _GEN_8406 = _T_260 ? satp : _GEN_8386; // @[decode.scala 469:28 680:39]
  wire [63:0] _GEN_8407 = _T_260 ? _mstatus_T_1 : _GEN_8387; // @[decode.scala 489:11 680:39]
  wire [126:0] _GEN_8408 = _T_260 ? 127'h8000000000101101 : _GEN_8388; // @[decode.scala 680:39 490:8]
  wire [63:0] _GEN_8409 = _T_260 ? medeleg : _GEN_8389; // @[decode.scala 472:28 680:39]
  wire [63:0] _GEN_8410 = _T_260 ? mideleg : _GEN_8390; // @[decode.scala 473:28 680:39]
  wire [63:0] _GEN_8411 = _T_260 ? mie : _GEN_8391; // @[decode.scala 474:28 680:39]
  wire [63:0] _GEN_8412 = _T_260 ? mtvec : _GEN_8392; // @[decode.scala 475:28 680:39]
  wire [63:0] _GEN_8413 = _T_260 ? mcounteren : _GEN_8393; // @[decode.scala 476:28 680:39]
  wire [63:0] _GEN_8414 = _T_260 ? mscratch : _GEN_8394; // @[decode.scala 477:28 680:39]
  wire [63:0] _GEN_8415 = _T_260 ? mepc : _GEN_8395; // @[decode.scala 478:28 680:39]
  wire [63:0] _GEN_8416 = _T_260 ? mcause : _GEN_8396; // @[decode.scala 479:28 680:39]
  wire [63:0] _GEN_8417 = _T_260 ? mtval : _GEN_8397; // @[decode.scala 480:28 680:39]
  wire [63:0] _GEN_8418 = _T_260 ? mip : _GEN_8398; // @[decode.scala 481:28 680:39]
  wire [63:0] _GEN_8419 = _T_260 ? pmpcfg0 : _GEN_8399; // @[decode.scala 482:28 680:39]
  wire [63:0] _GEN_8420 = _T_260 ? pmpaddr0 : _GEN_8400; // @[decode.scala 483:28 680:39]
  wire [63:0] _GEN_8421 = _T_260 ? mvendorid : _GEN_8401; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8422 = _T_260 ? marchid : _GEN_8402; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8423 = _T_260 ? mimpid : _GEN_8403; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8424 = _T_260 ? mhartid : _GEN_8404; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8425 = _T_259 ? _ucause_T_5 : ucause; // @[decode.scala 467:28 680:39 684:38]
  wire [63:0] _GEN_8426 = _T_259 ? scounteren : _GEN_8405; // @[decode.scala 468:28 680:39]
  wire [63:0] _GEN_8427 = _T_259 ? satp : _GEN_8406; // @[decode.scala 469:28 680:39]
  wire [63:0] _GEN_8428 = _T_259 ? _mstatus_T_1 : _GEN_8407; // @[decode.scala 489:11 680:39]
  wire [126:0] _GEN_8429 = _T_259 ? 127'h8000000000101101 : _GEN_8408; // @[decode.scala 680:39 490:8]
  wire [63:0] _GEN_8430 = _T_259 ? medeleg : _GEN_8409; // @[decode.scala 472:28 680:39]
  wire [63:0] _GEN_8431 = _T_259 ? mideleg : _GEN_8410; // @[decode.scala 473:28 680:39]
  wire [63:0] _GEN_8432 = _T_259 ? mie : _GEN_8411; // @[decode.scala 474:28 680:39]
  wire [63:0] _GEN_8433 = _T_259 ? mtvec : _GEN_8412; // @[decode.scala 475:28 680:39]
  wire [63:0] _GEN_8434 = _T_259 ? mcounteren : _GEN_8413; // @[decode.scala 476:28 680:39]
  wire [63:0] _GEN_8435 = _T_259 ? mscratch : _GEN_8414; // @[decode.scala 477:28 680:39]
  wire [63:0] _GEN_8436 = _T_259 ? mepc : _GEN_8415; // @[decode.scala 478:28 680:39]
  wire [63:0] _GEN_8437 = _T_259 ? mcause : _GEN_8416; // @[decode.scala 479:28 680:39]
  wire [63:0] _GEN_8438 = _T_259 ? mtval : _GEN_8417; // @[decode.scala 480:28 680:39]
  wire [63:0] _GEN_8439 = _T_259 ? mip : _GEN_8418; // @[decode.scala 481:28 680:39]
  wire [63:0] _GEN_8440 = _T_259 ? pmpcfg0 : _GEN_8419; // @[decode.scala 482:28 680:39]
  wire [63:0] _GEN_8441 = _T_259 ? pmpaddr0 : _GEN_8420; // @[decode.scala 483:28 680:39]
  wire [63:0] _GEN_8442 = _T_259 ? mvendorid : _GEN_8421; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8443 = _T_259 ? marchid : _GEN_8422; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8444 = _T_259 ? mimpid : _GEN_8423; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8445 = _T_259 ? mhartid : _GEN_8424; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8446 = _T_258 ? _uepc_T_5 : uepc; // @[decode.scala 466:28 680:39 683:38]
  wire [63:0] _GEN_8447 = _T_258 ? ucause : _GEN_8425; // @[decode.scala 467:28 680:39]
  wire [63:0] _GEN_8448 = _T_258 ? scounteren : _GEN_8426; // @[decode.scala 468:28 680:39]
  wire [63:0] _GEN_8449 = _T_258 ? satp : _GEN_8427; // @[decode.scala 469:28 680:39]
  wire [63:0] _GEN_8450 = _T_258 ? _mstatus_T_1 : _GEN_8428; // @[decode.scala 489:11 680:39]
  wire [126:0] _GEN_8451 = _T_258 ? 127'h8000000000101101 : _GEN_8429; // @[decode.scala 680:39 490:8]
  wire [63:0] _GEN_8452 = _T_258 ? medeleg : _GEN_8430; // @[decode.scala 472:28 680:39]
  wire [63:0] _GEN_8453 = _T_258 ? mideleg : _GEN_8431; // @[decode.scala 473:28 680:39]
  wire [63:0] _GEN_8454 = _T_258 ? mie : _GEN_8432; // @[decode.scala 474:28 680:39]
  wire [63:0] _GEN_8455 = _T_258 ? mtvec : _GEN_8433; // @[decode.scala 475:28 680:39]
  wire [63:0] _GEN_8456 = _T_258 ? mcounteren : _GEN_8434; // @[decode.scala 476:28 680:39]
  wire [63:0] _GEN_8457 = _T_258 ? mscratch : _GEN_8435; // @[decode.scala 477:28 680:39]
  wire [63:0] _GEN_8458 = _T_258 ? mepc : _GEN_8436; // @[decode.scala 478:28 680:39]
  wire [63:0] _GEN_8459 = _T_258 ? mcause : _GEN_8437; // @[decode.scala 479:28 680:39]
  wire [63:0] _GEN_8460 = _T_258 ? mtval : _GEN_8438; // @[decode.scala 480:28 680:39]
  wire [63:0] _GEN_8461 = _T_258 ? mip : _GEN_8439; // @[decode.scala 481:28 680:39]
  wire [63:0] _GEN_8462 = _T_258 ? pmpcfg0 : _GEN_8440; // @[decode.scala 482:28 680:39]
  wire [63:0] _GEN_8463 = _T_258 ? pmpaddr0 : _GEN_8441; // @[decode.scala 483:28 680:39]
  wire [63:0] _GEN_8464 = _T_258 ? mvendorid : _GEN_8442; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8465 = _T_258 ? marchid : _GEN_8443; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8466 = _T_258 ? mimpid : _GEN_8444; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8467 = _T_258 ? mhartid : _GEN_8445; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8468 = _T_257 ? _utvec_T_5 : utvec; // @[decode.scala 465:28 680:39 682:38]
  wire [63:0] _GEN_8469 = _T_257 ? uepc : _GEN_8446; // @[decode.scala 466:28 680:39]
  wire [63:0] _GEN_8470 = _T_257 ? ucause : _GEN_8447; // @[decode.scala 467:28 680:39]
  wire [63:0] _GEN_8471 = _T_257 ? scounteren : _GEN_8448; // @[decode.scala 468:28 680:39]
  wire [63:0] _GEN_8472 = _T_257 ? satp : _GEN_8449; // @[decode.scala 469:28 680:39]
  wire [63:0] _GEN_8473 = _T_257 ? _mstatus_T_1 : _GEN_8450; // @[decode.scala 489:11 680:39]
  wire [126:0] _GEN_8474 = _T_257 ? 127'h8000000000101101 : _GEN_8451; // @[decode.scala 680:39 490:8]
  wire [63:0] _GEN_8475 = _T_257 ? medeleg : _GEN_8452; // @[decode.scala 472:28 680:39]
  wire [63:0] _GEN_8476 = _T_257 ? mideleg : _GEN_8453; // @[decode.scala 473:28 680:39]
  wire [63:0] _GEN_8477 = _T_257 ? mie : _GEN_8454; // @[decode.scala 474:28 680:39]
  wire [63:0] _GEN_8478 = _T_257 ? mtvec : _GEN_8455; // @[decode.scala 475:28 680:39]
  wire [63:0] _GEN_8479 = _T_257 ? mcounteren : _GEN_8456; // @[decode.scala 476:28 680:39]
  wire [63:0] _GEN_8480 = _T_257 ? mscratch : _GEN_8457; // @[decode.scala 477:28 680:39]
  wire [63:0] _GEN_8481 = _T_257 ? mepc : _GEN_8458; // @[decode.scala 478:28 680:39]
  wire [63:0] _GEN_8482 = _T_257 ? mcause : _GEN_8459; // @[decode.scala 479:28 680:39]
  wire [63:0] _GEN_8483 = _T_257 ? mtval : _GEN_8460; // @[decode.scala 480:28 680:39]
  wire [63:0] _GEN_8484 = _T_257 ? mip : _GEN_8461; // @[decode.scala 481:28 680:39]
  wire [63:0] _GEN_8485 = _T_257 ? pmpcfg0 : _GEN_8462; // @[decode.scala 482:28 680:39]
  wire [63:0] _GEN_8486 = _T_257 ? pmpaddr0 : _GEN_8463; // @[decode.scala 483:28 680:39]
  wire [63:0] _GEN_8487 = _T_257 ? mvendorid : _GEN_8464; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8488 = _T_257 ? marchid : _GEN_8465; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8489 = _T_257 ? mimpid : _GEN_8466; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8490 = _T_257 ? mhartid : _GEN_8467; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8491 = _T_256 ? _ustatus_T_5 : ustatus; // @[decode.scala 464:28 680:39 681:38]
  wire [63:0] _GEN_8492 = _T_256 ? utvec : _GEN_8468; // @[decode.scala 465:28 680:39]
  wire [63:0] _GEN_8493 = _T_256 ? uepc : _GEN_8469; // @[decode.scala 466:28 680:39]
  wire [63:0] _GEN_8494 = _T_256 ? ucause : _GEN_8470; // @[decode.scala 467:28 680:39]
  wire [63:0] _GEN_8495 = _T_256 ? scounteren : _GEN_8471; // @[decode.scala 468:28 680:39]
  wire [63:0] _GEN_8496 = _T_256 ? satp : _GEN_8472; // @[decode.scala 469:28 680:39]
  wire [63:0] _GEN_8497 = _T_256 ? _mstatus_T_1 : _GEN_8473; // @[decode.scala 489:11 680:39]
  wire [126:0] _GEN_8498 = _T_256 ? 127'h8000000000101101 : _GEN_8474; // @[decode.scala 680:39 490:8]
  wire [63:0] _GEN_8499 = _T_256 ? medeleg : _GEN_8475; // @[decode.scala 472:28 680:39]
  wire [63:0] _GEN_8500 = _T_256 ? mideleg : _GEN_8476; // @[decode.scala 473:28 680:39]
  wire [63:0] _GEN_8501 = _T_256 ? mie : _GEN_8477; // @[decode.scala 474:28 680:39]
  wire [63:0] _GEN_8502 = _T_256 ? mtvec : _GEN_8478; // @[decode.scala 475:28 680:39]
  wire [63:0] _GEN_8503 = _T_256 ? mcounteren : _GEN_8479; // @[decode.scala 476:28 680:39]
  wire [63:0] _GEN_8504 = _T_256 ? mscratch : _GEN_8480; // @[decode.scala 477:28 680:39]
  wire [63:0] _GEN_8505 = _T_256 ? mepc : _GEN_8481; // @[decode.scala 478:28 680:39]
  wire [63:0] _GEN_8506 = _T_256 ? mcause : _GEN_8482; // @[decode.scala 479:28 680:39]
  wire [63:0] _GEN_8507 = _T_256 ? mtval : _GEN_8483; // @[decode.scala 480:28 680:39]
  wire [63:0] _GEN_8508 = _T_256 ? mip : _GEN_8484; // @[decode.scala 481:28 680:39]
  wire [63:0] _GEN_8509 = _T_256 ? pmpcfg0 : _GEN_8485; // @[decode.scala 482:28 680:39]
  wire [63:0] _GEN_8510 = _T_256 ? pmpaddr0 : _GEN_8486; // @[decode.scala 483:28 680:39]
  wire [63:0] _GEN_8511 = _T_256 ? mvendorid : _GEN_8487; // @[decode.scala 484:28 680:39]
  wire [63:0] _GEN_8512 = _T_256 ? marchid : _GEN_8488; // @[decode.scala 485:28 680:39]
  wire [63:0] _GEN_8513 = _T_256 ? mimpid : _GEN_8489; // @[decode.scala 486:28 680:39]
  wire [63:0] _GEN_8514 = _T_256 ? mhartid : _GEN_8490; // @[decode.scala 487:28 680:39]
  wire [63:0] _GEN_8515 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8491 : ustatus; // @[decode.scala 464:28 538:48]
  wire [63:0] _GEN_8516 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8492 : utvec; // @[decode.scala 465:28 538:48]
  wire [63:0] _GEN_8517 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8493 : uepc; // @[decode.scala 466:28 538:48]
  wire [63:0] _GEN_8518 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8494 : ucause; // @[decode.scala 467:28 538:48]
  wire [63:0] _GEN_8519 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8495 : scounteren; // @[decode.scala 468:28 538:48]
  wire [63:0] _GEN_8520 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8496 : satp; // @[decode.scala 469:28 538:48]
  wire [63:0] _GEN_8521 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8497 : _mstatus_T_1; // @[decode.scala 489:11 538:48]
  wire [126:0] _GEN_8522 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8498 : 127'h8000000000101101; // @[decode.scala 538:48 490:8]
  wire [63:0] _GEN_8523 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8499 : medeleg; // @[decode.scala 472:28 538:48]
  wire [63:0] _GEN_8524 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8500 : mideleg; // @[decode.scala 473:28 538:48]
  wire [63:0] _GEN_8525 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8501 : mie; // @[decode.scala 474:28 538:48]
  wire [63:0] _GEN_8526 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8502 : mtvec; // @[decode.scala 475:28 538:48]
  wire [63:0] _GEN_8527 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8503 : mcounteren; // @[decode.scala 476:28 538:48]
  wire [63:0] _GEN_8528 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8504 : mscratch; // @[decode.scala 477:28 538:48]
  wire [63:0] _GEN_8529 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8505 : mepc; // @[decode.scala 478:28 538:48]
  wire [63:0] _GEN_8530 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8506 : mcause; // @[decode.scala 479:28 538:48]
  wire [63:0] _GEN_8531 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8507 : mtval; // @[decode.scala 480:28 538:48]
  wire [63:0] _GEN_8532 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8508 : mip; // @[decode.scala 481:28 538:48]
  wire [63:0] _GEN_8533 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8509 : pmpcfg0; // @[decode.scala 482:28 538:48]
  wire [63:0] _GEN_8534 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8510 : pmpaddr0; // @[decode.scala 483:28 538:48]
  wire [63:0] _GEN_8535 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8511 : mvendorid; // @[decode.scala 484:28 538:48]
  wire [63:0] _GEN_8536 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8512 : marchid; // @[decode.scala 485:28 538:48]
  wire [63:0] _GEN_8537 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8513 : mimpid; // @[decode.scala 486:28 538:48]
  wire [63:0] _GEN_8538 = 3'h7 == writeBackResult_instruction[14:12] ? _GEN_8514 : mhartid; // @[decode.scala 487:28 538:48]
  wire [63:0] _GEN_8539 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8191 : _GEN_8515; // @[decode.scala 538:48]
  wire [63:0] _GEN_8540 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8192 : _GEN_8516; // @[decode.scala 538:48]
  wire [63:0] _GEN_8541 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8193 : _GEN_8517; // @[decode.scala 538:48]
  wire [63:0] _GEN_8542 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8194 : _GEN_8518; // @[decode.scala 538:48]
  wire [63:0] _GEN_8543 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8195 : _GEN_8519; // @[decode.scala 538:48]
  wire [63:0] _GEN_8544 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8196 : _GEN_8520; // @[decode.scala 538:48]
  wire [63:0] _GEN_8545 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8197 : _GEN_8521; // @[decode.scala 538:48]
  wire [126:0] _GEN_8546 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8198 : _GEN_8522; // @[decode.scala 538:48]
  wire [63:0] _GEN_8547 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8199 : _GEN_8523; // @[decode.scala 538:48]
  wire [63:0] _GEN_8548 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8200 : _GEN_8524; // @[decode.scala 538:48]
  wire [63:0] _GEN_8549 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8201 : _GEN_8525; // @[decode.scala 538:48]
  wire [63:0] _GEN_8550 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8202 : _GEN_8526; // @[decode.scala 538:48]
  wire [63:0] _GEN_8551 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8203 : _GEN_8527; // @[decode.scala 538:48]
  wire [63:0] _GEN_8552 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8204 : _GEN_8528; // @[decode.scala 538:48]
  wire [63:0] _GEN_8553 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8205 : _GEN_8529; // @[decode.scala 538:48]
  wire [63:0] _GEN_8554 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8206 : _GEN_8530; // @[decode.scala 538:48]
  wire [63:0] _GEN_8555 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8207 : _GEN_8531; // @[decode.scala 538:48]
  wire [63:0] _GEN_8556 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8208 : _GEN_8532; // @[decode.scala 538:48]
  wire [63:0] _GEN_8557 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8209 : _GEN_8533; // @[decode.scala 538:48]
  wire [63:0] _GEN_8558 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8210 : _GEN_8534; // @[decode.scala 538:48]
  wire [63:0] _GEN_8559 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8211 : _GEN_8535; // @[decode.scala 538:48]
  wire [63:0] _GEN_8560 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8212 : _GEN_8536; // @[decode.scala 538:48]
  wire [63:0] _GEN_8561 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8213 : _GEN_8537; // @[decode.scala 538:48]
  wire [63:0] _GEN_8562 = 3'h6 == writeBackResult_instruction[14:12] ? _GEN_8214 : _GEN_8538; // @[decode.scala 538:48]
  wire [63:0] _GEN_8563 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7891 : _GEN_8539; // @[decode.scala 538:48]
  wire [63:0] _GEN_8564 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7892 : _GEN_8540; // @[decode.scala 538:48]
  wire [63:0] _GEN_8565 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7893 : _GEN_8541; // @[decode.scala 538:48]
  wire [63:0] _GEN_8566 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7894 : _GEN_8542; // @[decode.scala 538:48]
  wire [63:0] _GEN_8567 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7895 : _GEN_8543; // @[decode.scala 538:48]
  wire [63:0] _GEN_8568 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7896 : _GEN_8544; // @[decode.scala 538:48]
  wire [63:0] _GEN_8569 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7897 : _GEN_8545; // @[decode.scala 538:48]
  wire [126:0] _GEN_8570 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7898 : _GEN_8546; // @[decode.scala 538:48]
  wire [63:0] _GEN_8571 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7899 : _GEN_8547; // @[decode.scala 538:48]
  wire [63:0] _GEN_8572 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7900 : _GEN_8548; // @[decode.scala 538:48]
  wire [63:0] _GEN_8573 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7901 : _GEN_8549; // @[decode.scala 538:48]
  wire [63:0] _GEN_8574 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7902 : _GEN_8550; // @[decode.scala 538:48]
  wire [63:0] _GEN_8575 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7903 : _GEN_8551; // @[decode.scala 538:48]
  wire [63:0] _GEN_8576 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7904 : _GEN_8552; // @[decode.scala 538:48]
  wire [63:0] _GEN_8577 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7905 : _GEN_8553; // @[decode.scala 538:48]
  wire [63:0] _GEN_8578 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7906 : _GEN_8554; // @[decode.scala 538:48]
  wire [63:0] _GEN_8579 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7907 : _GEN_8555; // @[decode.scala 538:48]
  wire [63:0] _GEN_8580 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7908 : _GEN_8556; // @[decode.scala 538:48]
  wire [63:0] _GEN_8581 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7909 : _GEN_8557; // @[decode.scala 538:48]
  wire [63:0] _GEN_8582 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7910 : _GEN_8558; // @[decode.scala 538:48]
  wire [63:0] _GEN_8583 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7911 : _GEN_8559; // @[decode.scala 538:48]
  wire [63:0] _GEN_8584 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7912 : _GEN_8560; // @[decode.scala 538:48]
  wire [63:0] _GEN_8585 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7913 : _GEN_8561; // @[decode.scala 538:48]
  wire [63:0] _GEN_8586 = 3'h5 == writeBackResult_instruction[14:12] ? _GEN_7914 : _GEN_8562; // @[decode.scala 538:48]
  wire [63:0] _GEN_8587 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7591 : _GEN_8563; // @[decode.scala 538:48]
  wire [63:0] _GEN_8588 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7592 : _GEN_8564; // @[decode.scala 538:48]
  wire [63:0] _GEN_8589 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7593 : _GEN_8565; // @[decode.scala 538:48]
  wire [63:0] _GEN_8590 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7594 : _GEN_8566; // @[decode.scala 538:48]
  wire [63:0] _GEN_8591 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7595 : _GEN_8567; // @[decode.scala 538:48]
  wire [63:0] _GEN_8592 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7596 : _GEN_8568; // @[decode.scala 538:48]
  wire [63:0] _GEN_8593 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7597 : _GEN_8569; // @[decode.scala 538:48]
  wire [126:0] _GEN_8594 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7598 : _GEN_8570; // @[decode.scala 538:48]
  wire [63:0] _GEN_8595 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7599 : _GEN_8571; // @[decode.scala 538:48]
  wire [63:0] _GEN_8596 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7600 : _GEN_8572; // @[decode.scala 538:48]
  wire [63:0] _GEN_8597 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7601 : _GEN_8573; // @[decode.scala 538:48]
  wire [63:0] _GEN_8598 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7602 : _GEN_8574; // @[decode.scala 538:48]
  wire [63:0] _GEN_8599 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7603 : _GEN_8575; // @[decode.scala 538:48]
  wire [63:0] _GEN_8600 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7604 : _GEN_8576; // @[decode.scala 538:48]
  wire [63:0] _GEN_8601 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7605 : _GEN_8577; // @[decode.scala 538:48]
  wire [63:0] _GEN_8602 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7606 : _GEN_8578; // @[decode.scala 538:48]
  wire [63:0] _GEN_8603 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7607 : _GEN_8579; // @[decode.scala 538:48]
  wire [63:0] _GEN_8604 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7608 : _GEN_8580; // @[decode.scala 538:48]
  wire [63:0] _GEN_8605 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7609 : _GEN_8581; // @[decode.scala 538:48]
  wire [63:0] _GEN_8606 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7610 : _GEN_8582; // @[decode.scala 538:48]
  wire [63:0] _GEN_8607 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7611 : _GEN_8583; // @[decode.scala 538:48]
  wire [63:0] _GEN_8608 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7612 : _GEN_8584; // @[decode.scala 538:48]
  wire [63:0] _GEN_8609 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7613 : _GEN_8585; // @[decode.scala 538:48]
  wire [63:0] _GEN_8610 = 3'h3 == writeBackResult_instruction[14:12] ? _GEN_7614 : _GEN_8586; // @[decode.scala 538:48]
  wire [63:0] _GEN_8617 = 3'h2 == writeBackResult_instruction[14:12] ? _GEN_7297 : _GEN_8593; // @[decode.scala 538:48]
  wire [126:0] _GEN_8618 = 3'h2 == writeBackResult_instruction[14:12] ? _GEN_7298 : _GEN_8594; // @[decode.scala 538:48]
  wire [63:0] _GEN_8625 = 3'h2 == writeBackResult_instruction[14:12] ? _GEN_7305 : _GEN_8601; // @[decode.scala 538:48]
  wire [63:0] _GEN_8626 = 3'h2 == writeBackResult_instruction[14:12] ? _GEN_7306 : _GEN_8602; // @[decode.scala 538:48]
  wire [63:0] _GEN_8641 = 3'h1 == writeBackResult_instruction[14:12] ? _GEN_6997 : _GEN_8617; // @[decode.scala 538:48]
  wire [126:0] _GEN_8642 = 3'h1 == writeBackResult_instruction[14:12] ? _GEN_6998 : _GEN_8618; // @[decode.scala 538:48]
  wire [63:0] _GEN_8649 = 3'h1 == writeBackResult_instruction[14:12] ? _GEN_7005 : _GEN_8625; // @[decode.scala 538:48]
  wire [63:0] _GEN_8650 = 3'h1 == writeBackResult_instruction[14:12] ? _GEN_7006 : _GEN_8626; // @[decode.scala 538:48]
  wire [63:0] _GEN_8666 = _T_246 & writeBackResult_instruction[14:12] != 3'h0 ? _GEN_8641 : _mstatus_T_1; // @[decode.scala 489:11 535:126]
  wire [126:0] _GEN_8667 = _T_246 & writeBackResult_instruction[14:12] != 3'h0 ? _GEN_8642 : 127'h8000000000101101; // @[decode.scala 535:126 490:8]
  wire [63:0] _GEN_8674 = _T_246 & writeBackResult_instruction[14:12] != 3'h0 ? _GEN_8649 : mepc; // @[decode.scala 535:126 478:28]
  wire [63:0] _GEN_8675 = _T_246 & writeBackResult_instruction[14:12] != 3'h0 ? _GEN_8650 : mcause; // @[decode.scala 535:126 479:28]
  reg [63:0] currentPrivilege; // @[decode.scala 710:33]
  wire [37:0] _GEN_8685 = mstatus[12] ? 38'h2200000000 : 38'h2200001800; // @[decode.scala 714:{24,24}]
  wire [63:0] _mstatus_T_9 = {60'ha0000008,mstatus[7:4]}; // @[Cat.scala 33:92]
  wire  _T_421 = currentPrivilege == 64'h2200000000; // @[decode.scala 720:29]
  wire [3:0] _GEN_8686 = currentPrivilege == 64'h2200000000 ? 4'hb : 4'h8; // @[decode.scala 720:{42,51} 721:27]
  wire [4:0] _mstatus_T_11 = _T_421 ? 5'h18 : 5'h0; // @[decode.scala 724:66]
  wire [63:0] _mstatus_T_13 = {51'h0,_mstatus_T_11,mstatus[3:0],4'h0}; // @[Cat.scala 33:92]
  wire [63:0] _mstatus_T_14 = 64'ha00000000 | _mstatus_T_13; // @[decode.scala 724:46]
  wire [63:0] _GEN_9883 = {{32'd0}, writeBackResult_instruction}; // @[decode.scala 725:44]
  wire [63:0] _mepc_T_6 = stallReg ? ecallPC : interruptedPC; // @[decode.scala 728:18]
  wire [63:0] _GEN_8687 = _GEN_9883 == 64'h80000073 ? _mepc_T_6 : _GEN_8674; // @[decode.scala 725:69 728:12]
  wire [63:0] _GEN_8688 = _GEN_9883 == 64'h80000073 ? 64'h8000000000000007 : _GEN_8675; // @[decode.scala 725:69 729:14]
  wire [63:0] _GEN_8689 = _GEN_9883 == 64'h80000073 ? 64'h2200000000 : currentPrivilege; // @[decode.scala 725:69 730:24 710:33]
  wire [63:0] _GEN_8690 = _GEN_9883 == 64'h80000073 ? mtvec : _GEN_6681; // @[decode.scala 725:69 731:18]
  wire [63:0] _GEN_8691 = _GEN_9883 == 64'h80000073 ? _mstatus_T_14 : _GEN_8666; // @[decode.scala 725:69 732:15]
  wire  _GEN_8771 = writeAddrPRF_exec1Valid ? 6'h0 == writeAddrPRF_exec1Addr | _GEN_1952 : _GEN_1952; // @[decode.scala 751:33]
  wire  _GEN_8772 = writeAddrPRF_exec1Valid ? 6'h1 == writeAddrPRF_exec1Addr | _GEN_1953 : _GEN_1953; // @[decode.scala 751:33]
  wire  _GEN_8773 = writeAddrPRF_exec1Valid ? 6'h2 == writeAddrPRF_exec1Addr | _GEN_1954 : _GEN_1954; // @[decode.scala 751:33]
  wire  _GEN_8774 = writeAddrPRF_exec1Valid ? 6'h3 == writeAddrPRF_exec1Addr | _GEN_1955 : _GEN_1955; // @[decode.scala 751:33]
  wire  _GEN_8775 = writeAddrPRF_exec1Valid ? 6'h4 == writeAddrPRF_exec1Addr | _GEN_1956 : _GEN_1956; // @[decode.scala 751:33]
  wire  _GEN_8776 = writeAddrPRF_exec1Valid ? 6'h5 == writeAddrPRF_exec1Addr | _GEN_1957 : _GEN_1957; // @[decode.scala 751:33]
  wire  _GEN_8777 = writeAddrPRF_exec1Valid ? 6'h6 == writeAddrPRF_exec1Addr | _GEN_1958 : _GEN_1958; // @[decode.scala 751:33]
  wire  _GEN_8778 = writeAddrPRF_exec1Valid ? 6'h7 == writeAddrPRF_exec1Addr | _GEN_1959 : _GEN_1959; // @[decode.scala 751:33]
  wire  _GEN_8779 = writeAddrPRF_exec1Valid ? 6'h8 == writeAddrPRF_exec1Addr | _GEN_1960 : _GEN_1960; // @[decode.scala 751:33]
  wire  _GEN_8780 = writeAddrPRF_exec1Valid ? 6'h9 == writeAddrPRF_exec1Addr | _GEN_1961 : _GEN_1961; // @[decode.scala 751:33]
  wire  _GEN_8781 = writeAddrPRF_exec1Valid ? 6'ha == writeAddrPRF_exec1Addr | _GEN_1962 : _GEN_1962; // @[decode.scala 751:33]
  wire  _GEN_8782 = writeAddrPRF_exec1Valid ? 6'hb == writeAddrPRF_exec1Addr | _GEN_1963 : _GEN_1963; // @[decode.scala 751:33]
  wire  _GEN_8783 = writeAddrPRF_exec1Valid ? 6'hc == writeAddrPRF_exec1Addr | _GEN_1964 : _GEN_1964; // @[decode.scala 751:33]
  wire  _GEN_8784 = writeAddrPRF_exec1Valid ? 6'hd == writeAddrPRF_exec1Addr | _GEN_1965 : _GEN_1965; // @[decode.scala 751:33]
  wire  _GEN_8785 = writeAddrPRF_exec1Valid ? 6'he == writeAddrPRF_exec1Addr | _GEN_1966 : _GEN_1966; // @[decode.scala 751:33]
  wire  _GEN_8786 = writeAddrPRF_exec1Valid ? 6'hf == writeAddrPRF_exec1Addr | _GEN_1967 : _GEN_1967; // @[decode.scala 751:33]
  wire  _GEN_8787 = writeAddrPRF_exec1Valid ? 6'h10 == writeAddrPRF_exec1Addr | _GEN_1968 : _GEN_1968; // @[decode.scala 751:33]
  wire  _GEN_8788 = writeAddrPRF_exec1Valid ? 6'h11 == writeAddrPRF_exec1Addr | _GEN_1969 : _GEN_1969; // @[decode.scala 751:33]
  wire  _GEN_8789 = writeAddrPRF_exec1Valid ? 6'h12 == writeAddrPRF_exec1Addr | _GEN_1970 : _GEN_1970; // @[decode.scala 751:33]
  wire  _GEN_8790 = writeAddrPRF_exec1Valid ? 6'h13 == writeAddrPRF_exec1Addr | _GEN_1971 : _GEN_1971; // @[decode.scala 751:33]
  wire  _GEN_8791 = writeAddrPRF_exec1Valid ? 6'h14 == writeAddrPRF_exec1Addr | _GEN_1972 : _GEN_1972; // @[decode.scala 751:33]
  wire  _GEN_8792 = writeAddrPRF_exec1Valid ? 6'h15 == writeAddrPRF_exec1Addr | _GEN_1973 : _GEN_1973; // @[decode.scala 751:33]
  wire  _GEN_8793 = writeAddrPRF_exec1Valid ? 6'h16 == writeAddrPRF_exec1Addr | _GEN_1974 : _GEN_1974; // @[decode.scala 751:33]
  wire  _GEN_8794 = writeAddrPRF_exec1Valid ? 6'h17 == writeAddrPRF_exec1Addr | _GEN_1975 : _GEN_1975; // @[decode.scala 751:33]
  wire  _GEN_8795 = writeAddrPRF_exec1Valid ? 6'h18 == writeAddrPRF_exec1Addr | _GEN_1976 : _GEN_1976; // @[decode.scala 751:33]
  wire  _GEN_8796 = writeAddrPRF_exec1Valid ? 6'h19 == writeAddrPRF_exec1Addr | _GEN_1977 : _GEN_1977; // @[decode.scala 751:33]
  wire  _GEN_8797 = writeAddrPRF_exec1Valid ? 6'h1a == writeAddrPRF_exec1Addr | _GEN_1978 : _GEN_1978; // @[decode.scala 751:33]
  wire  _GEN_8798 = writeAddrPRF_exec1Valid ? 6'h1b == writeAddrPRF_exec1Addr | _GEN_1979 : _GEN_1979; // @[decode.scala 751:33]
  wire  _GEN_8799 = writeAddrPRF_exec1Valid ? 6'h1c == writeAddrPRF_exec1Addr | _GEN_1980 : _GEN_1980; // @[decode.scala 751:33]
  wire  _GEN_8800 = writeAddrPRF_exec1Valid ? 6'h1d == writeAddrPRF_exec1Addr | _GEN_1981 : _GEN_1981; // @[decode.scala 751:33]
  wire  _GEN_8801 = writeAddrPRF_exec1Valid ? 6'h1e == writeAddrPRF_exec1Addr | _GEN_1982 : _GEN_1982; // @[decode.scala 751:33]
  wire  _GEN_8802 = writeAddrPRF_exec1Valid ? 6'h1f == writeAddrPRF_exec1Addr | _GEN_1983 : _GEN_1983; // @[decode.scala 751:33]
  wire  _GEN_8803 = writeAddrPRF_exec1Valid ? 6'h20 == writeAddrPRF_exec1Addr | _GEN_1984 : _GEN_1984; // @[decode.scala 751:33]
  wire  _GEN_8804 = writeAddrPRF_exec1Valid ? 6'h21 == writeAddrPRF_exec1Addr | _GEN_1985 : _GEN_1985; // @[decode.scala 751:33]
  wire  _GEN_8805 = writeAddrPRF_exec1Valid ? 6'h22 == writeAddrPRF_exec1Addr | _GEN_1986 : _GEN_1986; // @[decode.scala 751:33]
  wire  _GEN_8806 = writeAddrPRF_exec1Valid ? 6'h23 == writeAddrPRF_exec1Addr | _GEN_1987 : _GEN_1987; // @[decode.scala 751:33]
  wire  _GEN_8807 = writeAddrPRF_exec1Valid ? 6'h24 == writeAddrPRF_exec1Addr | _GEN_1988 : _GEN_1988; // @[decode.scala 751:33]
  wire  _GEN_8808 = writeAddrPRF_exec1Valid ? 6'h25 == writeAddrPRF_exec1Addr | _GEN_1989 : _GEN_1989; // @[decode.scala 751:33]
  wire  _GEN_8809 = writeAddrPRF_exec1Valid ? 6'h26 == writeAddrPRF_exec1Addr | _GEN_1990 : _GEN_1990; // @[decode.scala 751:33]
  wire  _GEN_8810 = writeAddrPRF_exec1Valid ? 6'h27 == writeAddrPRF_exec1Addr | _GEN_1991 : _GEN_1991; // @[decode.scala 751:33]
  wire  _GEN_8811 = writeAddrPRF_exec1Valid ? 6'h28 == writeAddrPRF_exec1Addr | _GEN_1992 : _GEN_1992; // @[decode.scala 751:33]
  wire  _GEN_8812 = writeAddrPRF_exec1Valid ? 6'h29 == writeAddrPRF_exec1Addr | _GEN_1993 : _GEN_1993; // @[decode.scala 751:33]
  wire  _GEN_8813 = writeAddrPRF_exec1Valid ? 6'h2a == writeAddrPRF_exec1Addr | _GEN_1994 : _GEN_1994; // @[decode.scala 751:33]
  wire  _GEN_8814 = writeAddrPRF_exec1Valid ? 6'h2b == writeAddrPRF_exec1Addr | _GEN_1995 : _GEN_1995; // @[decode.scala 751:33]
  wire  _GEN_8815 = writeAddrPRF_exec1Valid ? 6'h2c == writeAddrPRF_exec1Addr | _GEN_1996 : _GEN_1996; // @[decode.scala 751:33]
  wire  _GEN_8816 = writeAddrPRF_exec1Valid ? 6'h2d == writeAddrPRF_exec1Addr | _GEN_1997 : _GEN_1997; // @[decode.scala 751:33]
  wire  _GEN_8817 = writeAddrPRF_exec1Valid ? 6'h2e == writeAddrPRF_exec1Addr | _GEN_1998 : _GEN_1998; // @[decode.scala 751:33]
  wire  _GEN_8818 = writeAddrPRF_exec1Valid ? 6'h2f == writeAddrPRF_exec1Addr | _GEN_1999 : _GEN_1999; // @[decode.scala 751:33]
  wire  _GEN_8819 = writeAddrPRF_exec1Valid ? 6'h30 == writeAddrPRF_exec1Addr | _GEN_2000 : _GEN_2000; // @[decode.scala 751:33]
  wire  _GEN_8820 = writeAddrPRF_exec1Valid ? 6'h31 == writeAddrPRF_exec1Addr | _GEN_2001 : _GEN_2001; // @[decode.scala 751:33]
  wire  _GEN_8821 = writeAddrPRF_exec1Valid ? 6'h32 == writeAddrPRF_exec1Addr | _GEN_2002 : _GEN_2002; // @[decode.scala 751:33]
  wire  _GEN_8822 = writeAddrPRF_exec1Valid ? 6'h33 == writeAddrPRF_exec1Addr | _GEN_2003 : _GEN_2003; // @[decode.scala 751:33]
  wire  _GEN_8823 = writeAddrPRF_exec1Valid ? 6'h34 == writeAddrPRF_exec1Addr | _GEN_2004 : _GEN_2004; // @[decode.scala 751:33]
  wire  _GEN_8824 = writeAddrPRF_exec1Valid ? 6'h35 == writeAddrPRF_exec1Addr | _GEN_2005 : _GEN_2005; // @[decode.scala 751:33]
  wire  _GEN_8825 = writeAddrPRF_exec1Valid ? 6'h36 == writeAddrPRF_exec1Addr | _GEN_2006 : _GEN_2006; // @[decode.scala 751:33]
  wire  _GEN_8826 = writeAddrPRF_exec1Valid ? 6'h37 == writeAddrPRF_exec1Addr | _GEN_2007 : _GEN_2007; // @[decode.scala 751:33]
  wire  _GEN_8827 = writeAddrPRF_exec1Valid ? 6'h38 == writeAddrPRF_exec1Addr | _GEN_2008 : _GEN_2008; // @[decode.scala 751:33]
  wire  _GEN_8828 = writeAddrPRF_exec1Valid ? 6'h39 == writeAddrPRF_exec1Addr | _GEN_2009 : _GEN_2009; // @[decode.scala 751:33]
  wire  _GEN_8829 = writeAddrPRF_exec1Valid ? 6'h3a == writeAddrPRF_exec1Addr | _GEN_2010 : _GEN_2010; // @[decode.scala 751:33]
  wire  _GEN_8830 = writeAddrPRF_exec1Valid ? 6'h3b == writeAddrPRF_exec1Addr | _GEN_2011 : _GEN_2011; // @[decode.scala 751:33]
  wire  _GEN_8831 = writeAddrPRF_exec1Valid ? 6'h3c == writeAddrPRF_exec1Addr | _GEN_2012 : _GEN_2012; // @[decode.scala 751:33]
  wire  _GEN_8832 = writeAddrPRF_exec1Valid ? 6'h3d == writeAddrPRF_exec1Addr | _GEN_2013 : _GEN_2013; // @[decode.scala 751:33]
  wire  _GEN_8833 = writeAddrPRF_exec1Valid ? 6'h3e == writeAddrPRF_exec1Addr | _GEN_2014 : _GEN_2014; // @[decode.scala 751:33]
  wire  _GEN_8834 = writeAddrPRF_exec1Valid ? 6'h3f == writeAddrPRF_exec1Addr | _GEN_2015 : _GEN_2015; // @[decode.scala 751:33]
  wire  _GEN_8899 = writeAddrPRF_exec2Valid ? 6'h0 == writeAddrPRF_exec2Addr | _GEN_8771 : _GEN_8771; // @[decode.scala 752:33]
  wire  _GEN_8900 = writeAddrPRF_exec2Valid ? 6'h1 == writeAddrPRF_exec2Addr | _GEN_8772 : _GEN_8772; // @[decode.scala 752:33]
  wire  _GEN_8901 = writeAddrPRF_exec2Valid ? 6'h2 == writeAddrPRF_exec2Addr | _GEN_8773 : _GEN_8773; // @[decode.scala 752:33]
  wire  _GEN_8902 = writeAddrPRF_exec2Valid ? 6'h3 == writeAddrPRF_exec2Addr | _GEN_8774 : _GEN_8774; // @[decode.scala 752:33]
  wire  _GEN_8903 = writeAddrPRF_exec2Valid ? 6'h4 == writeAddrPRF_exec2Addr | _GEN_8775 : _GEN_8775; // @[decode.scala 752:33]
  wire  _GEN_8904 = writeAddrPRF_exec2Valid ? 6'h5 == writeAddrPRF_exec2Addr | _GEN_8776 : _GEN_8776; // @[decode.scala 752:33]
  wire  _GEN_8905 = writeAddrPRF_exec2Valid ? 6'h6 == writeAddrPRF_exec2Addr | _GEN_8777 : _GEN_8777; // @[decode.scala 752:33]
  wire  _GEN_8906 = writeAddrPRF_exec2Valid ? 6'h7 == writeAddrPRF_exec2Addr | _GEN_8778 : _GEN_8778; // @[decode.scala 752:33]
  wire  _GEN_8907 = writeAddrPRF_exec2Valid ? 6'h8 == writeAddrPRF_exec2Addr | _GEN_8779 : _GEN_8779; // @[decode.scala 752:33]
  wire  _GEN_8908 = writeAddrPRF_exec2Valid ? 6'h9 == writeAddrPRF_exec2Addr | _GEN_8780 : _GEN_8780; // @[decode.scala 752:33]
  wire  _GEN_8909 = writeAddrPRF_exec2Valid ? 6'ha == writeAddrPRF_exec2Addr | _GEN_8781 : _GEN_8781; // @[decode.scala 752:33]
  wire  _GEN_8910 = writeAddrPRF_exec2Valid ? 6'hb == writeAddrPRF_exec2Addr | _GEN_8782 : _GEN_8782; // @[decode.scala 752:33]
  wire  _GEN_8911 = writeAddrPRF_exec2Valid ? 6'hc == writeAddrPRF_exec2Addr | _GEN_8783 : _GEN_8783; // @[decode.scala 752:33]
  wire  _GEN_8912 = writeAddrPRF_exec2Valid ? 6'hd == writeAddrPRF_exec2Addr | _GEN_8784 : _GEN_8784; // @[decode.scala 752:33]
  wire  _GEN_8913 = writeAddrPRF_exec2Valid ? 6'he == writeAddrPRF_exec2Addr | _GEN_8785 : _GEN_8785; // @[decode.scala 752:33]
  wire  _GEN_8914 = writeAddrPRF_exec2Valid ? 6'hf == writeAddrPRF_exec2Addr | _GEN_8786 : _GEN_8786; // @[decode.scala 752:33]
  wire  _GEN_8915 = writeAddrPRF_exec2Valid ? 6'h10 == writeAddrPRF_exec2Addr | _GEN_8787 : _GEN_8787; // @[decode.scala 752:33]
  wire  _GEN_8916 = writeAddrPRF_exec2Valid ? 6'h11 == writeAddrPRF_exec2Addr | _GEN_8788 : _GEN_8788; // @[decode.scala 752:33]
  wire  _GEN_8917 = writeAddrPRF_exec2Valid ? 6'h12 == writeAddrPRF_exec2Addr | _GEN_8789 : _GEN_8789; // @[decode.scala 752:33]
  wire  _GEN_8918 = writeAddrPRF_exec2Valid ? 6'h13 == writeAddrPRF_exec2Addr | _GEN_8790 : _GEN_8790; // @[decode.scala 752:33]
  wire  _GEN_8919 = writeAddrPRF_exec2Valid ? 6'h14 == writeAddrPRF_exec2Addr | _GEN_8791 : _GEN_8791; // @[decode.scala 752:33]
  wire  _GEN_8920 = writeAddrPRF_exec2Valid ? 6'h15 == writeAddrPRF_exec2Addr | _GEN_8792 : _GEN_8792; // @[decode.scala 752:33]
  wire  _GEN_8921 = writeAddrPRF_exec2Valid ? 6'h16 == writeAddrPRF_exec2Addr | _GEN_8793 : _GEN_8793; // @[decode.scala 752:33]
  wire  _GEN_8922 = writeAddrPRF_exec2Valid ? 6'h17 == writeAddrPRF_exec2Addr | _GEN_8794 : _GEN_8794; // @[decode.scala 752:33]
  wire  _GEN_8923 = writeAddrPRF_exec2Valid ? 6'h18 == writeAddrPRF_exec2Addr | _GEN_8795 : _GEN_8795; // @[decode.scala 752:33]
  wire  _GEN_8924 = writeAddrPRF_exec2Valid ? 6'h19 == writeAddrPRF_exec2Addr | _GEN_8796 : _GEN_8796; // @[decode.scala 752:33]
  wire  _GEN_8925 = writeAddrPRF_exec2Valid ? 6'h1a == writeAddrPRF_exec2Addr | _GEN_8797 : _GEN_8797; // @[decode.scala 752:33]
  wire  _GEN_8926 = writeAddrPRF_exec2Valid ? 6'h1b == writeAddrPRF_exec2Addr | _GEN_8798 : _GEN_8798; // @[decode.scala 752:33]
  wire  _GEN_8927 = writeAddrPRF_exec2Valid ? 6'h1c == writeAddrPRF_exec2Addr | _GEN_8799 : _GEN_8799; // @[decode.scala 752:33]
  wire  _GEN_8928 = writeAddrPRF_exec2Valid ? 6'h1d == writeAddrPRF_exec2Addr | _GEN_8800 : _GEN_8800; // @[decode.scala 752:33]
  wire  _GEN_8929 = writeAddrPRF_exec2Valid ? 6'h1e == writeAddrPRF_exec2Addr | _GEN_8801 : _GEN_8801; // @[decode.scala 752:33]
  wire  _GEN_8930 = writeAddrPRF_exec2Valid ? 6'h1f == writeAddrPRF_exec2Addr | _GEN_8802 : _GEN_8802; // @[decode.scala 752:33]
  wire  _GEN_8931 = writeAddrPRF_exec2Valid ? 6'h20 == writeAddrPRF_exec2Addr | _GEN_8803 : _GEN_8803; // @[decode.scala 752:33]
  wire  _GEN_8932 = writeAddrPRF_exec2Valid ? 6'h21 == writeAddrPRF_exec2Addr | _GEN_8804 : _GEN_8804; // @[decode.scala 752:33]
  wire  _GEN_8933 = writeAddrPRF_exec2Valid ? 6'h22 == writeAddrPRF_exec2Addr | _GEN_8805 : _GEN_8805; // @[decode.scala 752:33]
  wire  _GEN_8934 = writeAddrPRF_exec2Valid ? 6'h23 == writeAddrPRF_exec2Addr | _GEN_8806 : _GEN_8806; // @[decode.scala 752:33]
  wire  _GEN_8935 = writeAddrPRF_exec2Valid ? 6'h24 == writeAddrPRF_exec2Addr | _GEN_8807 : _GEN_8807; // @[decode.scala 752:33]
  wire  _GEN_8936 = writeAddrPRF_exec2Valid ? 6'h25 == writeAddrPRF_exec2Addr | _GEN_8808 : _GEN_8808; // @[decode.scala 752:33]
  wire  _GEN_8937 = writeAddrPRF_exec2Valid ? 6'h26 == writeAddrPRF_exec2Addr | _GEN_8809 : _GEN_8809; // @[decode.scala 752:33]
  wire  _GEN_8938 = writeAddrPRF_exec2Valid ? 6'h27 == writeAddrPRF_exec2Addr | _GEN_8810 : _GEN_8810; // @[decode.scala 752:33]
  wire  _GEN_8939 = writeAddrPRF_exec2Valid ? 6'h28 == writeAddrPRF_exec2Addr | _GEN_8811 : _GEN_8811; // @[decode.scala 752:33]
  wire  _GEN_8940 = writeAddrPRF_exec2Valid ? 6'h29 == writeAddrPRF_exec2Addr | _GEN_8812 : _GEN_8812; // @[decode.scala 752:33]
  wire  _GEN_8941 = writeAddrPRF_exec2Valid ? 6'h2a == writeAddrPRF_exec2Addr | _GEN_8813 : _GEN_8813; // @[decode.scala 752:33]
  wire  _GEN_8942 = writeAddrPRF_exec2Valid ? 6'h2b == writeAddrPRF_exec2Addr | _GEN_8814 : _GEN_8814; // @[decode.scala 752:33]
  wire  _GEN_8943 = writeAddrPRF_exec2Valid ? 6'h2c == writeAddrPRF_exec2Addr | _GEN_8815 : _GEN_8815; // @[decode.scala 752:33]
  wire  _GEN_8944 = writeAddrPRF_exec2Valid ? 6'h2d == writeAddrPRF_exec2Addr | _GEN_8816 : _GEN_8816; // @[decode.scala 752:33]
  wire  _GEN_8945 = writeAddrPRF_exec2Valid ? 6'h2e == writeAddrPRF_exec2Addr | _GEN_8817 : _GEN_8817; // @[decode.scala 752:33]
  wire  _GEN_8946 = writeAddrPRF_exec2Valid ? 6'h2f == writeAddrPRF_exec2Addr | _GEN_8818 : _GEN_8818; // @[decode.scala 752:33]
  wire  _GEN_8947 = writeAddrPRF_exec2Valid ? 6'h30 == writeAddrPRF_exec2Addr | _GEN_8819 : _GEN_8819; // @[decode.scala 752:33]
  wire  _GEN_8948 = writeAddrPRF_exec2Valid ? 6'h31 == writeAddrPRF_exec2Addr | _GEN_8820 : _GEN_8820; // @[decode.scala 752:33]
  wire  _GEN_8949 = writeAddrPRF_exec2Valid ? 6'h32 == writeAddrPRF_exec2Addr | _GEN_8821 : _GEN_8821; // @[decode.scala 752:33]
  wire  _GEN_8950 = writeAddrPRF_exec2Valid ? 6'h33 == writeAddrPRF_exec2Addr | _GEN_8822 : _GEN_8822; // @[decode.scala 752:33]
  wire  _GEN_8951 = writeAddrPRF_exec2Valid ? 6'h34 == writeAddrPRF_exec2Addr | _GEN_8823 : _GEN_8823; // @[decode.scala 752:33]
  wire  _GEN_8952 = writeAddrPRF_exec2Valid ? 6'h35 == writeAddrPRF_exec2Addr | _GEN_8824 : _GEN_8824; // @[decode.scala 752:33]
  wire  _GEN_8953 = writeAddrPRF_exec2Valid ? 6'h36 == writeAddrPRF_exec2Addr | _GEN_8825 : _GEN_8825; // @[decode.scala 752:33]
  wire  _GEN_8954 = writeAddrPRF_exec2Valid ? 6'h37 == writeAddrPRF_exec2Addr | _GEN_8826 : _GEN_8826; // @[decode.scala 752:33]
  wire  _GEN_8955 = writeAddrPRF_exec2Valid ? 6'h38 == writeAddrPRF_exec2Addr | _GEN_8827 : _GEN_8827; // @[decode.scala 752:33]
  wire  _GEN_8956 = writeAddrPRF_exec2Valid ? 6'h39 == writeAddrPRF_exec2Addr | _GEN_8828 : _GEN_8828; // @[decode.scala 752:33]
  wire  _GEN_8957 = writeAddrPRF_exec2Valid ? 6'h3a == writeAddrPRF_exec2Addr | _GEN_8829 : _GEN_8829; // @[decode.scala 752:33]
  wire  _GEN_8958 = writeAddrPRF_exec2Valid ? 6'h3b == writeAddrPRF_exec2Addr | _GEN_8830 : _GEN_8830; // @[decode.scala 752:33]
  wire  _GEN_8959 = writeAddrPRF_exec2Valid ? 6'h3c == writeAddrPRF_exec2Addr | _GEN_8831 : _GEN_8831; // @[decode.scala 752:33]
  wire  _GEN_8960 = writeAddrPRF_exec2Valid ? 6'h3d == writeAddrPRF_exec2Addr | _GEN_8832 : _GEN_8832; // @[decode.scala 752:33]
  wire  _GEN_8961 = writeAddrPRF_exec2Valid ? 6'h3e == writeAddrPRF_exec2Addr | _GEN_8833 : _GEN_8833; // @[decode.scala 752:33]
  wire  _GEN_8962 = writeAddrPRF_exec2Valid ? 6'h3f == writeAddrPRF_exec2Addr | _GEN_8834 : _GEN_8834; // @[decode.scala 752:33]
  wire  _GEN_9027 = writeAddrPRF_exec3Valid ? 6'h0 == writeAddrPRF_exec3Addr | _GEN_8899 : _GEN_8899; // @[decode.scala 753:33]
  wire  _GEN_9028 = writeAddrPRF_exec3Valid ? 6'h1 == writeAddrPRF_exec3Addr | _GEN_8900 : _GEN_8900; // @[decode.scala 753:33]
  wire  _GEN_9029 = writeAddrPRF_exec3Valid ? 6'h2 == writeAddrPRF_exec3Addr | _GEN_8901 : _GEN_8901; // @[decode.scala 753:33]
  wire  _GEN_9030 = writeAddrPRF_exec3Valid ? 6'h3 == writeAddrPRF_exec3Addr | _GEN_8902 : _GEN_8902; // @[decode.scala 753:33]
  wire  _GEN_9031 = writeAddrPRF_exec3Valid ? 6'h4 == writeAddrPRF_exec3Addr | _GEN_8903 : _GEN_8903; // @[decode.scala 753:33]
  wire  _GEN_9032 = writeAddrPRF_exec3Valid ? 6'h5 == writeAddrPRF_exec3Addr | _GEN_8904 : _GEN_8904; // @[decode.scala 753:33]
  wire  _GEN_9033 = writeAddrPRF_exec3Valid ? 6'h6 == writeAddrPRF_exec3Addr | _GEN_8905 : _GEN_8905; // @[decode.scala 753:33]
  wire  _GEN_9034 = writeAddrPRF_exec3Valid ? 6'h7 == writeAddrPRF_exec3Addr | _GEN_8906 : _GEN_8906; // @[decode.scala 753:33]
  wire  _GEN_9035 = writeAddrPRF_exec3Valid ? 6'h8 == writeAddrPRF_exec3Addr | _GEN_8907 : _GEN_8907; // @[decode.scala 753:33]
  wire  _GEN_9036 = writeAddrPRF_exec3Valid ? 6'h9 == writeAddrPRF_exec3Addr | _GEN_8908 : _GEN_8908; // @[decode.scala 753:33]
  wire  _GEN_9037 = writeAddrPRF_exec3Valid ? 6'ha == writeAddrPRF_exec3Addr | _GEN_8909 : _GEN_8909; // @[decode.scala 753:33]
  wire  _GEN_9038 = writeAddrPRF_exec3Valid ? 6'hb == writeAddrPRF_exec3Addr | _GEN_8910 : _GEN_8910; // @[decode.scala 753:33]
  wire  _GEN_9039 = writeAddrPRF_exec3Valid ? 6'hc == writeAddrPRF_exec3Addr | _GEN_8911 : _GEN_8911; // @[decode.scala 753:33]
  wire  _GEN_9040 = writeAddrPRF_exec3Valid ? 6'hd == writeAddrPRF_exec3Addr | _GEN_8912 : _GEN_8912; // @[decode.scala 753:33]
  wire  _GEN_9041 = writeAddrPRF_exec3Valid ? 6'he == writeAddrPRF_exec3Addr | _GEN_8913 : _GEN_8913; // @[decode.scala 753:33]
  wire  _GEN_9042 = writeAddrPRF_exec3Valid ? 6'hf == writeAddrPRF_exec3Addr | _GEN_8914 : _GEN_8914; // @[decode.scala 753:33]
  wire  _GEN_9043 = writeAddrPRF_exec3Valid ? 6'h10 == writeAddrPRF_exec3Addr | _GEN_8915 : _GEN_8915; // @[decode.scala 753:33]
  wire  _GEN_9044 = writeAddrPRF_exec3Valid ? 6'h11 == writeAddrPRF_exec3Addr | _GEN_8916 : _GEN_8916; // @[decode.scala 753:33]
  wire  _GEN_9045 = writeAddrPRF_exec3Valid ? 6'h12 == writeAddrPRF_exec3Addr | _GEN_8917 : _GEN_8917; // @[decode.scala 753:33]
  wire  _GEN_9046 = writeAddrPRF_exec3Valid ? 6'h13 == writeAddrPRF_exec3Addr | _GEN_8918 : _GEN_8918; // @[decode.scala 753:33]
  wire  _GEN_9047 = writeAddrPRF_exec3Valid ? 6'h14 == writeAddrPRF_exec3Addr | _GEN_8919 : _GEN_8919; // @[decode.scala 753:33]
  wire  _GEN_9048 = writeAddrPRF_exec3Valid ? 6'h15 == writeAddrPRF_exec3Addr | _GEN_8920 : _GEN_8920; // @[decode.scala 753:33]
  wire  _GEN_9049 = writeAddrPRF_exec3Valid ? 6'h16 == writeAddrPRF_exec3Addr | _GEN_8921 : _GEN_8921; // @[decode.scala 753:33]
  wire  _GEN_9050 = writeAddrPRF_exec3Valid ? 6'h17 == writeAddrPRF_exec3Addr | _GEN_8922 : _GEN_8922; // @[decode.scala 753:33]
  wire  _GEN_9051 = writeAddrPRF_exec3Valid ? 6'h18 == writeAddrPRF_exec3Addr | _GEN_8923 : _GEN_8923; // @[decode.scala 753:33]
  wire  _GEN_9052 = writeAddrPRF_exec3Valid ? 6'h19 == writeAddrPRF_exec3Addr | _GEN_8924 : _GEN_8924; // @[decode.scala 753:33]
  wire  _GEN_9053 = writeAddrPRF_exec3Valid ? 6'h1a == writeAddrPRF_exec3Addr | _GEN_8925 : _GEN_8925; // @[decode.scala 753:33]
  wire  _GEN_9054 = writeAddrPRF_exec3Valid ? 6'h1b == writeAddrPRF_exec3Addr | _GEN_8926 : _GEN_8926; // @[decode.scala 753:33]
  wire  _GEN_9055 = writeAddrPRF_exec3Valid ? 6'h1c == writeAddrPRF_exec3Addr | _GEN_8927 : _GEN_8927; // @[decode.scala 753:33]
  wire  _GEN_9056 = writeAddrPRF_exec3Valid ? 6'h1d == writeAddrPRF_exec3Addr | _GEN_8928 : _GEN_8928; // @[decode.scala 753:33]
  wire  _GEN_9057 = writeAddrPRF_exec3Valid ? 6'h1e == writeAddrPRF_exec3Addr | _GEN_8929 : _GEN_8929; // @[decode.scala 753:33]
  wire  _GEN_9058 = writeAddrPRF_exec3Valid ? 6'h1f == writeAddrPRF_exec3Addr | _GEN_8930 : _GEN_8930; // @[decode.scala 753:33]
  wire  _GEN_9091 = _T_212 | stateRegInputBuf; // @[decode.scala 771:58 772:32 187:34]
  wire  _GEN_9092 = fromFetch_expected_valid ? _GEN_9091 : 1'h1; // @[decode.scala 770:42 775:30]
  wire  _GEN_9097 = branchEvalIn_fired & ~branchEvalIn_passFail ? 1'h0 : _GEN_6714; // @[decode.scala 761:58 765:18]
  wire  _GEN_9099 = ~fromFetch_fired | _T_214 & fun3 == 3'h0 & immediate_immediate == 64'h302 ? 1'h0 : stateRegInputBuf; // @[decode.scala 794:100 795:32 187:34]
  wire  _GEN_9101 = readyOutputBuf ? _GEN_9099 : stateRegInputBuf; // @[decode.scala 792:32 187:34]
  wire  _GEN_9104 = ~stall & ~(branchEvalIn_fired & (opcode == 7'h63 | opcode == 7'h6f | opcode == 7'h67)) ? _GEN_9101
     : stateRegInputBuf; // @[decode.scala 790:114 187:34]
  wire  _GEN_9118 = validInputBuf | stateRegOutputBuf; // @[decode.scala 822:29 823:29 188:34]
  wire  _GEN_9122 = ~validInputBuf ? 1'h0 : stateRegOutputBuf; // @[decode.scala 836:32 837:31 188:34]
  wire  _GEN_9124 = toExec_fired ? _GEN_9122 : stateRegOutputBuf; // @[decode.scala 834:28 188:34]
  wire  _T_456 = writeBackResult_instruction[6:0] != 7'h63; // @[decode.scala 852:38]
  wire  _T_457 = writeBackResult_fired & writeBackResult_rdAddr != 5'h0 & _T_456; // @[decode.scala 851:61]
  wire  _T_459 = writeBackResult_instruction[6:0] != 7'h23; // @[decode.scala 853:38]
  wire  _T_460 = _T_457 & _T_459; // @[decode.scala 852:50]
  wire [5:0] _GEN_9135 = 5'h1 == writeBackResult_rdAddr ? architecturalRegMap_1 : architecturalRegMap_0; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9136 = 5'h2 == writeBackResult_rdAddr ? architecturalRegMap_2 : _GEN_9135; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9137 = 5'h3 == writeBackResult_rdAddr ? architecturalRegMap_3 : _GEN_9136; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9138 = 5'h4 == writeBackResult_rdAddr ? architecturalRegMap_4 : _GEN_9137; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9139 = 5'h5 == writeBackResult_rdAddr ? architecturalRegMap_5 : _GEN_9138; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9140 = 5'h6 == writeBackResult_rdAddr ? architecturalRegMap_6 : _GEN_9139; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9141 = 5'h7 == writeBackResult_rdAddr ? architecturalRegMap_7 : _GEN_9140; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9142 = 5'h8 == writeBackResult_rdAddr ? architecturalRegMap_8 : _GEN_9141; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9143 = 5'h9 == writeBackResult_rdAddr ? architecturalRegMap_9 : _GEN_9142; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9144 = 5'ha == writeBackResult_rdAddr ? architecturalRegMap_10 : _GEN_9143; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9145 = 5'hb == writeBackResult_rdAddr ? architecturalRegMap_11 : _GEN_9144; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9146 = 5'hc == writeBackResult_rdAddr ? architecturalRegMap_12 : _GEN_9145; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9147 = 5'hd == writeBackResult_rdAddr ? architecturalRegMap_13 : _GEN_9146; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9148 = 5'he == writeBackResult_rdAddr ? architecturalRegMap_14 : _GEN_9147; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9149 = 5'hf == writeBackResult_rdAddr ? architecturalRegMap_15 : _GEN_9148; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9150 = 5'h10 == writeBackResult_rdAddr ? architecturalRegMap_16 : _GEN_9149; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9151 = 5'h11 == writeBackResult_rdAddr ? architecturalRegMap_17 : _GEN_9150; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9152 = 5'h12 == writeBackResult_rdAddr ? architecturalRegMap_18 : _GEN_9151; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9153 = 5'h13 == writeBackResult_rdAddr ? architecturalRegMap_19 : _GEN_9152; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9154 = 5'h14 == writeBackResult_rdAddr ? architecturalRegMap_20 : _GEN_9153; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9155 = 5'h15 == writeBackResult_rdAddr ? architecturalRegMap_21 : _GEN_9154; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9156 = 5'h16 == writeBackResult_rdAddr ? architecturalRegMap_22 : _GEN_9155; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9157 = 5'h17 == writeBackResult_rdAddr ? architecturalRegMap_23 : _GEN_9156; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9158 = 5'h18 == writeBackResult_rdAddr ? architecturalRegMap_24 : _GEN_9157; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9159 = 5'h19 == writeBackResult_rdAddr ? architecturalRegMap_25 : _GEN_9158; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9160 = 5'h1a == writeBackResult_rdAddr ? architecturalRegMap_26 : _GEN_9159; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9161 = 5'h1b == writeBackResult_rdAddr ? architecturalRegMap_27 : _GEN_9160; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9162 = 5'h1c == writeBackResult_rdAddr ? architecturalRegMap_28 : _GEN_9161; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9163 = 5'h1d == writeBackResult_rdAddr ? architecturalRegMap_29 : _GEN_9162; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9164 = 5'h1e == writeBackResult_rdAddr ? architecturalRegMap_30 : _GEN_9163; // @[decode.scala 854:{49,49}]
  wire [5:0] _GEN_9165 = 5'h1f == writeBackResult_rdAddr ? architecturalRegMap_31 : _GEN_9164; // @[decode.scala 854:{49,49}]
  wire  _T_461 = _GEN_9165 != writeBackResult_PRFDest; // @[decode.scala 854:49]
  wire  _T_462 = _T_460 & _T_461; // @[decode.scala 853:50]
  wire  _T_463 = writeBackResult_instruction != 32'h80000073; // @[decode.scala 855:33]
  wire  _T_464 = _T_462 & _T_463; // @[decode.scala 854:77]
  wire  _GEN_10076 = 6'h0 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9198 = 6'h0 == _GEN_9165 | _GEN_1888; // @[decode.scala 858:{62,62}]
  wire  _GEN_10077 = 6'h1 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9199 = 6'h1 == _GEN_9165 | _GEN_1889; // @[decode.scala 858:{62,62}]
  wire  _GEN_10078 = 6'h2 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9200 = 6'h2 == _GEN_9165 | _GEN_1890; // @[decode.scala 858:{62,62}]
  wire  _GEN_10079 = 6'h3 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9201 = 6'h3 == _GEN_9165 | _GEN_1891; // @[decode.scala 858:{62,62}]
  wire  _GEN_10080 = 6'h4 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9202 = 6'h4 == _GEN_9165 | _GEN_1892; // @[decode.scala 858:{62,62}]
  wire  _GEN_10081 = 6'h5 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9203 = 6'h5 == _GEN_9165 | _GEN_1893; // @[decode.scala 858:{62,62}]
  wire  _GEN_10082 = 6'h6 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9204 = 6'h6 == _GEN_9165 | _GEN_1894; // @[decode.scala 858:{62,62}]
  wire  _GEN_10083 = 6'h7 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9205 = 6'h7 == _GEN_9165 | _GEN_1895; // @[decode.scala 858:{62,62}]
  wire  _GEN_10084 = 6'h8 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9206 = 6'h8 == _GEN_9165 | _GEN_1896; // @[decode.scala 858:{62,62}]
  wire  _GEN_10085 = 6'h9 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9207 = 6'h9 == _GEN_9165 | _GEN_1897; // @[decode.scala 858:{62,62}]
  wire  _GEN_10086 = 6'ha == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9208 = 6'ha == _GEN_9165 | _GEN_1898; // @[decode.scala 858:{62,62}]
  wire  _GEN_10087 = 6'hb == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9209 = 6'hb == _GEN_9165 | _GEN_1899; // @[decode.scala 858:{62,62}]
  wire  _GEN_10088 = 6'hc == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9210 = 6'hc == _GEN_9165 | _GEN_1900; // @[decode.scala 858:{62,62}]
  wire  _GEN_10089 = 6'hd == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9211 = 6'hd == _GEN_9165 | _GEN_1901; // @[decode.scala 858:{62,62}]
  wire  _GEN_10090 = 6'he == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9212 = 6'he == _GEN_9165 | _GEN_1902; // @[decode.scala 858:{62,62}]
  wire  _GEN_10091 = 6'hf == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9213 = 6'hf == _GEN_9165 | _GEN_1903; // @[decode.scala 858:{62,62}]
  wire  _GEN_10092 = 6'h10 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9214 = 6'h10 == _GEN_9165 | _GEN_1904; // @[decode.scala 858:{62,62}]
  wire  _GEN_10093 = 6'h11 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9215 = 6'h11 == _GEN_9165 | _GEN_1905; // @[decode.scala 858:{62,62}]
  wire  _GEN_10094 = 6'h12 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9216 = 6'h12 == _GEN_9165 | _GEN_1906; // @[decode.scala 858:{62,62}]
  wire  _GEN_10095 = 6'h13 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9217 = 6'h13 == _GEN_9165 | _GEN_1907; // @[decode.scala 858:{62,62}]
  wire  _GEN_10096 = 6'h14 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9218 = 6'h14 == _GEN_9165 | _GEN_1908; // @[decode.scala 858:{62,62}]
  wire  _GEN_10097 = 6'h15 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9219 = 6'h15 == _GEN_9165 | _GEN_1909; // @[decode.scala 858:{62,62}]
  wire  _GEN_10098 = 6'h16 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9220 = 6'h16 == _GEN_9165 | _GEN_1910; // @[decode.scala 858:{62,62}]
  wire  _GEN_10099 = 6'h17 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9221 = 6'h17 == _GEN_9165 | _GEN_1911; // @[decode.scala 858:{62,62}]
  wire  _GEN_10100 = 6'h18 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9222 = 6'h18 == _GEN_9165 | _GEN_1912; // @[decode.scala 858:{62,62}]
  wire  _GEN_10101 = 6'h19 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9223 = 6'h19 == _GEN_9165 | _GEN_1913; // @[decode.scala 858:{62,62}]
  wire  _GEN_10102 = 6'h1a == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9224 = 6'h1a == _GEN_9165 | _GEN_1914; // @[decode.scala 858:{62,62}]
  wire  _GEN_10103 = 6'h1b == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9225 = 6'h1b == _GEN_9165 | _GEN_1915; // @[decode.scala 858:{62,62}]
  wire  _GEN_10104 = 6'h1c == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9226 = 6'h1c == _GEN_9165 | _GEN_1916; // @[decode.scala 858:{62,62}]
  wire  _GEN_10105 = 6'h1d == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9227 = 6'h1d == _GEN_9165 | _GEN_1917; // @[decode.scala 858:{62,62}]
  wire  _GEN_10106 = 6'h1e == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9228 = 6'h1e == _GEN_9165 | _GEN_1918; // @[decode.scala 858:{62,62}]
  wire  _GEN_10107 = 6'h1f == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9229 = 6'h1f == _GEN_9165 | _GEN_1919; // @[decode.scala 858:{62,62}]
  wire  _GEN_10108 = 6'h20 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9230 = 6'h20 == _GEN_9165 | _GEN_1920; // @[decode.scala 858:{62,62}]
  wire  _GEN_10109 = 6'h21 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9231 = 6'h21 == _GEN_9165 | _GEN_1921; // @[decode.scala 858:{62,62}]
  wire  _GEN_10110 = 6'h22 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9232 = 6'h22 == _GEN_9165 | _GEN_1922; // @[decode.scala 858:{62,62}]
  wire  _GEN_10111 = 6'h23 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9233 = 6'h23 == _GEN_9165 | _GEN_1923; // @[decode.scala 858:{62,62}]
  wire  _GEN_10112 = 6'h24 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9234 = 6'h24 == _GEN_9165 | _GEN_1924; // @[decode.scala 858:{62,62}]
  wire  _GEN_10113 = 6'h25 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9235 = 6'h25 == _GEN_9165 | _GEN_1925; // @[decode.scala 858:{62,62}]
  wire  _GEN_10114 = 6'h26 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9236 = 6'h26 == _GEN_9165 | _GEN_1926; // @[decode.scala 858:{62,62}]
  wire  _GEN_10115 = 6'h27 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9237 = 6'h27 == _GEN_9165 | _GEN_1927; // @[decode.scala 858:{62,62}]
  wire  _GEN_10116 = 6'h28 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9238 = 6'h28 == _GEN_9165 | _GEN_1928; // @[decode.scala 858:{62,62}]
  wire  _GEN_10117 = 6'h29 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9239 = 6'h29 == _GEN_9165 | _GEN_1929; // @[decode.scala 858:{62,62}]
  wire  _GEN_10118 = 6'h2a == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9240 = 6'h2a == _GEN_9165 | _GEN_1930; // @[decode.scala 858:{62,62}]
  wire  _GEN_10119 = 6'h2b == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9241 = 6'h2b == _GEN_9165 | _GEN_1931; // @[decode.scala 858:{62,62}]
  wire  _GEN_10120 = 6'h2c == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9242 = 6'h2c == _GEN_9165 | _GEN_1932; // @[decode.scala 858:{62,62}]
  wire  _GEN_10121 = 6'h2d == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9243 = 6'h2d == _GEN_9165 | _GEN_1933; // @[decode.scala 858:{62,62}]
  wire  _GEN_10122 = 6'h2e == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9244 = 6'h2e == _GEN_9165 | _GEN_1934; // @[decode.scala 858:{62,62}]
  wire  _GEN_10123 = 6'h2f == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9245 = 6'h2f == _GEN_9165 | _GEN_1935; // @[decode.scala 858:{62,62}]
  wire  _GEN_10124 = 6'h30 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9246 = 6'h30 == _GEN_9165 | _GEN_1936; // @[decode.scala 858:{62,62}]
  wire  _GEN_10125 = 6'h31 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9247 = 6'h31 == _GEN_9165 | _GEN_1937; // @[decode.scala 858:{62,62}]
  wire  _GEN_10126 = 6'h32 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9248 = 6'h32 == _GEN_9165 | _GEN_1938; // @[decode.scala 858:{62,62}]
  wire  _GEN_10127 = 6'h33 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9249 = 6'h33 == _GEN_9165 | _GEN_1939; // @[decode.scala 858:{62,62}]
  wire  _GEN_10128 = 6'h34 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9250 = 6'h34 == _GEN_9165 | _GEN_1940; // @[decode.scala 858:{62,62}]
  wire  _GEN_10129 = 6'h35 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9251 = 6'h35 == _GEN_9165 | _GEN_1941; // @[decode.scala 858:{62,62}]
  wire  _GEN_10130 = 6'h36 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9252 = 6'h36 == _GEN_9165 | _GEN_1942; // @[decode.scala 858:{62,62}]
  wire  _GEN_10131 = 6'h37 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9253 = 6'h37 == _GEN_9165 | _GEN_1943; // @[decode.scala 858:{62,62}]
  wire  _GEN_10132 = 6'h38 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9254 = 6'h38 == _GEN_9165 | _GEN_1944; // @[decode.scala 858:{62,62}]
  wire  _GEN_10133 = 6'h39 == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9255 = 6'h39 == _GEN_9165 | _GEN_1945; // @[decode.scala 858:{62,62}]
  wire  _GEN_10134 = 6'h3a == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9256 = 6'h3a == _GEN_9165 | _GEN_1946; // @[decode.scala 858:{62,62}]
  wire  _GEN_10135 = 6'h3b == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9257 = 6'h3b == _GEN_9165 | _GEN_1947; // @[decode.scala 858:{62,62}]
  wire  _GEN_10136 = 6'h3c == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9258 = 6'h3c == _GEN_9165 | _GEN_1948; // @[decode.scala 858:{62,62}]
  wire  _GEN_10137 = 6'h3d == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9259 = 6'h3d == _GEN_9165 | _GEN_1949; // @[decode.scala 858:{62,62}]
  wire  _GEN_10138 = 6'h3e == _GEN_9165; // @[decode.scala 858:{62,62}]
  wire  _GEN_9260 = 6'h3e == _GEN_9165 | _GEN_1950; // @[decode.scala 858:{62,62}]
  wire  _GEN_9262 = _GEN_10076 | _GEN_6071; // @[decode.scala 859:{68,68}]
  wire  _GEN_9263 = _GEN_10077 | _GEN_6072; // @[decode.scala 859:{68,68}]
  wire  _GEN_9264 = _GEN_10078 | _GEN_6073; // @[decode.scala 859:{68,68}]
  wire  _GEN_9265 = _GEN_10079 | _GEN_6074; // @[decode.scala 859:{68,68}]
  wire  _GEN_9266 = _GEN_10080 | _GEN_6075; // @[decode.scala 859:{68,68}]
  wire  _GEN_9267 = _GEN_10081 | _GEN_6076; // @[decode.scala 859:{68,68}]
  wire  _GEN_9268 = _GEN_10082 | _GEN_6077; // @[decode.scala 859:{68,68}]
  wire  _GEN_9269 = _GEN_10083 | _GEN_6078; // @[decode.scala 859:{68,68}]
  wire  _GEN_9270 = _GEN_10084 | _GEN_6079; // @[decode.scala 859:{68,68}]
  wire  _GEN_9271 = _GEN_10085 | _GEN_6080; // @[decode.scala 859:{68,68}]
  wire  _GEN_9272 = _GEN_10086 | _GEN_6081; // @[decode.scala 859:{68,68}]
  wire  _GEN_9273 = _GEN_10087 | _GEN_6082; // @[decode.scala 859:{68,68}]
  wire  _GEN_9274 = _GEN_10088 | _GEN_6083; // @[decode.scala 859:{68,68}]
  wire  _GEN_9275 = _GEN_10089 | _GEN_6084; // @[decode.scala 859:{68,68}]
  wire  _GEN_9276 = _GEN_10090 | _GEN_6085; // @[decode.scala 859:{68,68}]
  wire  _GEN_9277 = _GEN_10091 | _GEN_6086; // @[decode.scala 859:{68,68}]
  wire  _GEN_9278 = _GEN_10092 | _GEN_6087; // @[decode.scala 859:{68,68}]
  wire  _GEN_9279 = _GEN_10093 | _GEN_6088; // @[decode.scala 859:{68,68}]
  wire  _GEN_9280 = _GEN_10094 | _GEN_6089; // @[decode.scala 859:{68,68}]
  wire  _GEN_9281 = _GEN_10095 | _GEN_6090; // @[decode.scala 859:{68,68}]
  wire  _GEN_9282 = _GEN_10096 | _GEN_6091; // @[decode.scala 859:{68,68}]
  wire  _GEN_9283 = _GEN_10097 | _GEN_6092; // @[decode.scala 859:{68,68}]
  wire  _GEN_9284 = _GEN_10098 | _GEN_6093; // @[decode.scala 859:{68,68}]
  wire  _GEN_9285 = _GEN_10099 | _GEN_6094; // @[decode.scala 859:{68,68}]
  wire  _GEN_9286 = _GEN_10100 | _GEN_6095; // @[decode.scala 859:{68,68}]
  wire  _GEN_9287 = _GEN_10101 | _GEN_6096; // @[decode.scala 859:{68,68}]
  wire  _GEN_9288 = _GEN_10102 | _GEN_6097; // @[decode.scala 859:{68,68}]
  wire  _GEN_9289 = _GEN_10103 | _GEN_6098; // @[decode.scala 859:{68,68}]
  wire  _GEN_9290 = _GEN_10104 | _GEN_6099; // @[decode.scala 859:{68,68}]
  wire  _GEN_9291 = _GEN_10105 | _GEN_6100; // @[decode.scala 859:{68,68}]
  wire  _GEN_9292 = _GEN_10106 | _GEN_6101; // @[decode.scala 859:{68,68}]
  wire  _GEN_9293 = _GEN_10107 | _GEN_6102; // @[decode.scala 859:{68,68}]
  wire  _GEN_9294 = _GEN_10108 | _GEN_6103; // @[decode.scala 859:{68,68}]
  wire  _GEN_9295 = _GEN_10109 | _GEN_6104; // @[decode.scala 859:{68,68}]
  wire  _GEN_9296 = _GEN_10110 | _GEN_6105; // @[decode.scala 859:{68,68}]
  wire  _GEN_9297 = _GEN_10111 | _GEN_6106; // @[decode.scala 859:{68,68}]
  wire  _GEN_9298 = _GEN_10112 | _GEN_6107; // @[decode.scala 859:{68,68}]
  wire  _GEN_9299 = _GEN_10113 | _GEN_6108; // @[decode.scala 859:{68,68}]
  wire  _GEN_9300 = _GEN_10114 | _GEN_6109; // @[decode.scala 859:{68,68}]
  wire  _GEN_9301 = _GEN_10115 | _GEN_6110; // @[decode.scala 859:{68,68}]
  wire  _GEN_9302 = _GEN_10116 | _GEN_6111; // @[decode.scala 859:{68,68}]
  wire  _GEN_9303 = _GEN_10117 | _GEN_6112; // @[decode.scala 859:{68,68}]
  wire  _GEN_9304 = _GEN_10118 | _GEN_6113; // @[decode.scala 859:{68,68}]
  wire  _GEN_9305 = _GEN_10119 | _GEN_6114; // @[decode.scala 859:{68,68}]
  wire  _GEN_9306 = _GEN_10120 | _GEN_6115; // @[decode.scala 859:{68,68}]
  wire  _GEN_9307 = _GEN_10121 | _GEN_6116; // @[decode.scala 859:{68,68}]
  wire  _GEN_9308 = _GEN_10122 | _GEN_6117; // @[decode.scala 859:{68,68}]
  wire  _GEN_9309 = _GEN_10123 | _GEN_6118; // @[decode.scala 859:{68,68}]
  wire  _GEN_9310 = _GEN_10124 | _GEN_6119; // @[decode.scala 859:{68,68}]
  wire  _GEN_9311 = _GEN_10125 | _GEN_6120; // @[decode.scala 859:{68,68}]
  wire  _GEN_9312 = _GEN_10126 | _GEN_6121; // @[decode.scala 859:{68,68}]
  wire  _GEN_9313 = _GEN_10127 | _GEN_6122; // @[decode.scala 859:{68,68}]
  wire  _GEN_9314 = _GEN_10128 | _GEN_6123; // @[decode.scala 859:{68,68}]
  wire  _GEN_9315 = _GEN_10129 | _GEN_6124; // @[decode.scala 859:{68,68}]
  wire  _GEN_9316 = _GEN_10130 | _GEN_6125; // @[decode.scala 859:{68,68}]
  wire  _GEN_9317 = _GEN_10131 | _GEN_6126; // @[decode.scala 859:{68,68}]
  wire  _GEN_9318 = _GEN_10132 | _GEN_6127; // @[decode.scala 859:{68,68}]
  wire  _GEN_9319 = _GEN_10133 | _GEN_6128; // @[decode.scala 859:{68,68}]
  wire  _GEN_9320 = _GEN_10134 | _GEN_6129; // @[decode.scala 859:{68,68}]
  wire  _GEN_9321 = _GEN_10135 | _GEN_6130; // @[decode.scala 859:{68,68}]
  wire  _GEN_9322 = _GEN_10136 | _GEN_6131; // @[decode.scala 859:{68,68}]
  wire  _GEN_9323 = _GEN_10137 | _GEN_6132; // @[decode.scala 859:{68,68}]
  wire  _GEN_9324 = _GEN_10138 | _GEN_6133; // @[decode.scala 859:{68,68}]
  wire  _GEN_9326 = _GEN_10076 | _GEN_6231; // @[decode.scala 860:{68,68}]
  wire  _GEN_9327 = _GEN_10077 | _GEN_6232; // @[decode.scala 860:{68,68}]
  wire  _GEN_9328 = _GEN_10078 | _GEN_6233; // @[decode.scala 860:{68,68}]
  wire  _GEN_9329 = _GEN_10079 | _GEN_6234; // @[decode.scala 860:{68,68}]
  wire  _GEN_9330 = _GEN_10080 | _GEN_6235; // @[decode.scala 860:{68,68}]
  wire  _GEN_9331 = _GEN_10081 | _GEN_6236; // @[decode.scala 860:{68,68}]
  wire  _GEN_9332 = _GEN_10082 | _GEN_6237; // @[decode.scala 860:{68,68}]
  wire  _GEN_9333 = _GEN_10083 | _GEN_6238; // @[decode.scala 860:{68,68}]
  wire  _GEN_9334 = _GEN_10084 | _GEN_6239; // @[decode.scala 860:{68,68}]
  wire  _GEN_9335 = _GEN_10085 | _GEN_6240; // @[decode.scala 860:{68,68}]
  wire  _GEN_9336 = _GEN_10086 | _GEN_6241; // @[decode.scala 860:{68,68}]
  wire  _GEN_9337 = _GEN_10087 | _GEN_6242; // @[decode.scala 860:{68,68}]
  wire  _GEN_9338 = _GEN_10088 | _GEN_6243; // @[decode.scala 860:{68,68}]
  wire  _GEN_9339 = _GEN_10089 | _GEN_6244; // @[decode.scala 860:{68,68}]
  wire  _GEN_9340 = _GEN_10090 | _GEN_6245; // @[decode.scala 860:{68,68}]
  wire  _GEN_9341 = _GEN_10091 | _GEN_6246; // @[decode.scala 860:{68,68}]
  wire  _GEN_9342 = _GEN_10092 | _GEN_6247; // @[decode.scala 860:{68,68}]
  wire  _GEN_9343 = _GEN_10093 | _GEN_6248; // @[decode.scala 860:{68,68}]
  wire  _GEN_9344 = _GEN_10094 | _GEN_6249; // @[decode.scala 860:{68,68}]
  wire  _GEN_9345 = _GEN_10095 | _GEN_6250; // @[decode.scala 860:{68,68}]
  wire  _GEN_9346 = _GEN_10096 | _GEN_6251; // @[decode.scala 860:{68,68}]
  wire  _GEN_9347 = _GEN_10097 | _GEN_6252; // @[decode.scala 860:{68,68}]
  wire  _GEN_9348 = _GEN_10098 | _GEN_6253; // @[decode.scala 860:{68,68}]
  wire  _GEN_9349 = _GEN_10099 | _GEN_6254; // @[decode.scala 860:{68,68}]
  wire  _GEN_9350 = _GEN_10100 | _GEN_6255; // @[decode.scala 860:{68,68}]
  wire  _GEN_9351 = _GEN_10101 | _GEN_6256; // @[decode.scala 860:{68,68}]
  wire  _GEN_9352 = _GEN_10102 | _GEN_6257; // @[decode.scala 860:{68,68}]
  wire  _GEN_9353 = _GEN_10103 | _GEN_6258; // @[decode.scala 860:{68,68}]
  wire  _GEN_9354 = _GEN_10104 | _GEN_6259; // @[decode.scala 860:{68,68}]
  wire  _GEN_9355 = _GEN_10105 | _GEN_6260; // @[decode.scala 860:{68,68}]
  wire  _GEN_9356 = _GEN_10106 | _GEN_6261; // @[decode.scala 860:{68,68}]
  wire  _GEN_9357 = _GEN_10107 | _GEN_6262; // @[decode.scala 860:{68,68}]
  wire  _GEN_9358 = _GEN_10108 | _GEN_6263; // @[decode.scala 860:{68,68}]
  wire  _GEN_9359 = _GEN_10109 | _GEN_6264; // @[decode.scala 860:{68,68}]
  wire  _GEN_9360 = _GEN_10110 | _GEN_6265; // @[decode.scala 860:{68,68}]
  wire  _GEN_9361 = _GEN_10111 | _GEN_6266; // @[decode.scala 860:{68,68}]
  wire  _GEN_9362 = _GEN_10112 | _GEN_6267; // @[decode.scala 860:{68,68}]
  wire  _GEN_9363 = _GEN_10113 | _GEN_6268; // @[decode.scala 860:{68,68}]
  wire  _GEN_9364 = _GEN_10114 | _GEN_6269; // @[decode.scala 860:{68,68}]
  wire  _GEN_9365 = _GEN_10115 | _GEN_6270; // @[decode.scala 860:{68,68}]
  wire  _GEN_9366 = _GEN_10116 | _GEN_6271; // @[decode.scala 860:{68,68}]
  wire  _GEN_9367 = _GEN_10117 | _GEN_6272; // @[decode.scala 860:{68,68}]
  wire  _GEN_9368 = _GEN_10118 | _GEN_6273; // @[decode.scala 860:{68,68}]
  wire  _GEN_9369 = _GEN_10119 | _GEN_6274; // @[decode.scala 860:{68,68}]
  wire  _GEN_9370 = _GEN_10120 | _GEN_6275; // @[decode.scala 860:{68,68}]
  wire  _GEN_9371 = _GEN_10121 | _GEN_6276; // @[decode.scala 860:{68,68}]
  wire  _GEN_9372 = _GEN_10122 | _GEN_6277; // @[decode.scala 860:{68,68}]
  wire  _GEN_9373 = _GEN_10123 | _GEN_6278; // @[decode.scala 860:{68,68}]
  wire  _GEN_9374 = _GEN_10124 | _GEN_6279; // @[decode.scala 860:{68,68}]
  wire  _GEN_9375 = _GEN_10125 | _GEN_6280; // @[decode.scala 860:{68,68}]
  wire  _GEN_9376 = _GEN_10126 | _GEN_6281; // @[decode.scala 860:{68,68}]
  wire  _GEN_9377 = _GEN_10127 | _GEN_6282; // @[decode.scala 860:{68,68}]
  wire  _GEN_9378 = _GEN_10128 | _GEN_6283; // @[decode.scala 860:{68,68}]
  wire  _GEN_9379 = _GEN_10129 | _GEN_6284; // @[decode.scala 860:{68,68}]
  wire  _GEN_9380 = _GEN_10130 | _GEN_6285; // @[decode.scala 860:{68,68}]
  wire  _GEN_9381 = _GEN_10131 | _GEN_6286; // @[decode.scala 860:{68,68}]
  wire  _GEN_9382 = _GEN_10132 | _GEN_6287; // @[decode.scala 860:{68,68}]
  wire  _GEN_9383 = _GEN_10133 | _GEN_6288; // @[decode.scala 860:{68,68}]
  wire  _GEN_9384 = _GEN_10134 | _GEN_6289; // @[decode.scala 860:{68,68}]
  wire  _GEN_9385 = _GEN_10135 | _GEN_6290; // @[decode.scala 860:{68,68}]
  wire  _GEN_9386 = _GEN_10136 | _GEN_6291; // @[decode.scala 860:{68,68}]
  wire  _GEN_9387 = _GEN_10137 | _GEN_6292; // @[decode.scala 860:{68,68}]
  wire  _GEN_9388 = _GEN_10138 | _GEN_6293; // @[decode.scala 860:{68,68}]
  wire  _GEN_9390 = _GEN_10076 | _GEN_6391; // @[decode.scala 861:{68,68}]
  wire  _GEN_9391 = _GEN_10077 | _GEN_6392; // @[decode.scala 861:{68,68}]
  wire  _GEN_9392 = _GEN_10078 | _GEN_6393; // @[decode.scala 861:{68,68}]
  wire  _GEN_9393 = _GEN_10079 | _GEN_6394; // @[decode.scala 861:{68,68}]
  wire  _GEN_9394 = _GEN_10080 | _GEN_6395; // @[decode.scala 861:{68,68}]
  wire  _GEN_9395 = _GEN_10081 | _GEN_6396; // @[decode.scala 861:{68,68}]
  wire  _GEN_9396 = _GEN_10082 | _GEN_6397; // @[decode.scala 861:{68,68}]
  wire  _GEN_9397 = _GEN_10083 | _GEN_6398; // @[decode.scala 861:{68,68}]
  wire  _GEN_9398 = _GEN_10084 | _GEN_6399; // @[decode.scala 861:{68,68}]
  wire  _GEN_9399 = _GEN_10085 | _GEN_6400; // @[decode.scala 861:{68,68}]
  wire  _GEN_9400 = _GEN_10086 | _GEN_6401; // @[decode.scala 861:{68,68}]
  wire  _GEN_9401 = _GEN_10087 | _GEN_6402; // @[decode.scala 861:{68,68}]
  wire  _GEN_9402 = _GEN_10088 | _GEN_6403; // @[decode.scala 861:{68,68}]
  wire  _GEN_9403 = _GEN_10089 | _GEN_6404; // @[decode.scala 861:{68,68}]
  wire  _GEN_9404 = _GEN_10090 | _GEN_6405; // @[decode.scala 861:{68,68}]
  wire  _GEN_9405 = _GEN_10091 | _GEN_6406; // @[decode.scala 861:{68,68}]
  wire  _GEN_9406 = _GEN_10092 | _GEN_6407; // @[decode.scala 861:{68,68}]
  wire  _GEN_9407 = _GEN_10093 | _GEN_6408; // @[decode.scala 861:{68,68}]
  wire  _GEN_9408 = _GEN_10094 | _GEN_6409; // @[decode.scala 861:{68,68}]
  wire  _GEN_9409 = _GEN_10095 | _GEN_6410; // @[decode.scala 861:{68,68}]
  wire  _GEN_9410 = _GEN_10096 | _GEN_6411; // @[decode.scala 861:{68,68}]
  wire  _GEN_9411 = _GEN_10097 | _GEN_6412; // @[decode.scala 861:{68,68}]
  wire  _GEN_9412 = _GEN_10098 | _GEN_6413; // @[decode.scala 861:{68,68}]
  wire  _GEN_9413 = _GEN_10099 | _GEN_6414; // @[decode.scala 861:{68,68}]
  wire  _GEN_9414 = _GEN_10100 | _GEN_6415; // @[decode.scala 861:{68,68}]
  wire  _GEN_9415 = _GEN_10101 | _GEN_6416; // @[decode.scala 861:{68,68}]
  wire  _GEN_9416 = _GEN_10102 | _GEN_6417; // @[decode.scala 861:{68,68}]
  wire  _GEN_9417 = _GEN_10103 | _GEN_6418; // @[decode.scala 861:{68,68}]
  wire  _GEN_9418 = _GEN_10104 | _GEN_6419; // @[decode.scala 861:{68,68}]
  wire  _GEN_9419 = _GEN_10105 | _GEN_6420; // @[decode.scala 861:{68,68}]
  wire  _GEN_9420 = _GEN_10106 | _GEN_6421; // @[decode.scala 861:{68,68}]
  wire  _GEN_9421 = _GEN_10107 | _GEN_6422; // @[decode.scala 861:{68,68}]
  wire  _GEN_9422 = _GEN_10108 | _GEN_6423; // @[decode.scala 861:{68,68}]
  wire  _GEN_9423 = _GEN_10109 | _GEN_6424; // @[decode.scala 861:{68,68}]
  wire  _GEN_9424 = _GEN_10110 | _GEN_6425; // @[decode.scala 861:{68,68}]
  wire  _GEN_9425 = _GEN_10111 | _GEN_6426; // @[decode.scala 861:{68,68}]
  wire  _GEN_9426 = _GEN_10112 | _GEN_6427; // @[decode.scala 861:{68,68}]
  wire  _GEN_9427 = _GEN_10113 | _GEN_6428; // @[decode.scala 861:{68,68}]
  wire  _GEN_9428 = _GEN_10114 | _GEN_6429; // @[decode.scala 861:{68,68}]
  wire  _GEN_9429 = _GEN_10115 | _GEN_6430; // @[decode.scala 861:{68,68}]
  wire  _GEN_9430 = _GEN_10116 | _GEN_6431; // @[decode.scala 861:{68,68}]
  wire  _GEN_9431 = _GEN_10117 | _GEN_6432; // @[decode.scala 861:{68,68}]
  wire  _GEN_9432 = _GEN_10118 | _GEN_6433; // @[decode.scala 861:{68,68}]
  wire  _GEN_9433 = _GEN_10119 | _GEN_6434; // @[decode.scala 861:{68,68}]
  wire  _GEN_9434 = _GEN_10120 | _GEN_6435; // @[decode.scala 861:{68,68}]
  wire  _GEN_9435 = _GEN_10121 | _GEN_6436; // @[decode.scala 861:{68,68}]
  wire  _GEN_9436 = _GEN_10122 | _GEN_6437; // @[decode.scala 861:{68,68}]
  wire  _GEN_9437 = _GEN_10123 | _GEN_6438; // @[decode.scala 861:{68,68}]
  wire  _GEN_9438 = _GEN_10124 | _GEN_6439; // @[decode.scala 861:{68,68}]
  wire  _GEN_9439 = _GEN_10125 | _GEN_6440; // @[decode.scala 861:{68,68}]
  wire  _GEN_9440 = _GEN_10126 | _GEN_6441; // @[decode.scala 861:{68,68}]
  wire  _GEN_9441 = _GEN_10127 | _GEN_6442; // @[decode.scala 861:{68,68}]
  wire  _GEN_9442 = _GEN_10128 | _GEN_6443; // @[decode.scala 861:{68,68}]
  wire  _GEN_9443 = _GEN_10129 | _GEN_6444; // @[decode.scala 861:{68,68}]
  wire  _GEN_9444 = _GEN_10130 | _GEN_6445; // @[decode.scala 861:{68,68}]
  wire  _GEN_9445 = _GEN_10131 | _GEN_6446; // @[decode.scala 861:{68,68}]
  wire  _GEN_9446 = _GEN_10132 | _GEN_6447; // @[decode.scala 861:{68,68}]
  wire  _GEN_9447 = _GEN_10133 | _GEN_6448; // @[decode.scala 861:{68,68}]
  wire  _GEN_9448 = _GEN_10134 | _GEN_6449; // @[decode.scala 861:{68,68}]
  wire  _GEN_9449 = _GEN_10135 | _GEN_6450; // @[decode.scala 861:{68,68}]
  wire  _GEN_9450 = _GEN_10136 | _GEN_6451; // @[decode.scala 861:{68,68}]
  wire  _GEN_9451 = _GEN_10137 | _GEN_6452; // @[decode.scala 861:{68,68}]
  wire  _GEN_9452 = _GEN_10138 | _GEN_6453; // @[decode.scala 861:{68,68}]
  wire  _GEN_9454 = _GEN_10076 | _GEN_6551; // @[decode.scala 862:{68,68}]
  wire  _GEN_9455 = _GEN_10077 | _GEN_6552; // @[decode.scala 862:{68,68}]
  wire  _GEN_9456 = _GEN_10078 | _GEN_6553; // @[decode.scala 862:{68,68}]
  wire  _GEN_9457 = _GEN_10079 | _GEN_6554; // @[decode.scala 862:{68,68}]
  wire  _GEN_9458 = _GEN_10080 | _GEN_6555; // @[decode.scala 862:{68,68}]
  wire  _GEN_9459 = _GEN_10081 | _GEN_6556; // @[decode.scala 862:{68,68}]
  wire  _GEN_9460 = _GEN_10082 | _GEN_6557; // @[decode.scala 862:{68,68}]
  wire  _GEN_9461 = _GEN_10083 | _GEN_6558; // @[decode.scala 862:{68,68}]
  wire  _GEN_9462 = _GEN_10084 | _GEN_6559; // @[decode.scala 862:{68,68}]
  wire  _GEN_9463 = _GEN_10085 | _GEN_6560; // @[decode.scala 862:{68,68}]
  wire  _GEN_9464 = _GEN_10086 | _GEN_6561; // @[decode.scala 862:{68,68}]
  wire  _GEN_9465 = _GEN_10087 | _GEN_6562; // @[decode.scala 862:{68,68}]
  wire  _GEN_9466 = _GEN_10088 | _GEN_6563; // @[decode.scala 862:{68,68}]
  wire  _GEN_9467 = _GEN_10089 | _GEN_6564; // @[decode.scala 862:{68,68}]
  wire  _GEN_9468 = _GEN_10090 | _GEN_6565; // @[decode.scala 862:{68,68}]
  wire  _GEN_9469 = _GEN_10091 | _GEN_6566; // @[decode.scala 862:{68,68}]
  wire  _GEN_9470 = _GEN_10092 | _GEN_6567; // @[decode.scala 862:{68,68}]
  wire  _GEN_9471 = _GEN_10093 | _GEN_6568; // @[decode.scala 862:{68,68}]
  wire  _GEN_9472 = _GEN_10094 | _GEN_6569; // @[decode.scala 862:{68,68}]
  wire  _GEN_9473 = _GEN_10095 | _GEN_6570; // @[decode.scala 862:{68,68}]
  wire  _GEN_9474 = _GEN_10096 | _GEN_6571; // @[decode.scala 862:{68,68}]
  wire  _GEN_9475 = _GEN_10097 | _GEN_6572; // @[decode.scala 862:{68,68}]
  wire  _GEN_9476 = _GEN_10098 | _GEN_6573; // @[decode.scala 862:{68,68}]
  wire  _GEN_9477 = _GEN_10099 | _GEN_6574; // @[decode.scala 862:{68,68}]
  wire  _GEN_9478 = _GEN_10100 | _GEN_6575; // @[decode.scala 862:{68,68}]
  wire  _GEN_9479 = _GEN_10101 | _GEN_6576; // @[decode.scala 862:{68,68}]
  wire  _GEN_9480 = _GEN_10102 | _GEN_6577; // @[decode.scala 862:{68,68}]
  wire  _GEN_9481 = _GEN_10103 | _GEN_6578; // @[decode.scala 862:{68,68}]
  wire  _GEN_9482 = _GEN_10104 | _GEN_6579; // @[decode.scala 862:{68,68}]
  wire  _GEN_9483 = _GEN_10105 | _GEN_6580; // @[decode.scala 862:{68,68}]
  wire  _GEN_9484 = _GEN_10106 | _GEN_6581; // @[decode.scala 862:{68,68}]
  wire  _GEN_9485 = _GEN_10107 | _GEN_6582; // @[decode.scala 862:{68,68}]
  wire  _GEN_9486 = _GEN_10108 | _GEN_6583; // @[decode.scala 862:{68,68}]
  wire  _GEN_9487 = _GEN_10109 | _GEN_6584; // @[decode.scala 862:{68,68}]
  wire  _GEN_9488 = _GEN_10110 | _GEN_6585; // @[decode.scala 862:{68,68}]
  wire  _GEN_9489 = _GEN_10111 | _GEN_6586; // @[decode.scala 862:{68,68}]
  wire  _GEN_9490 = _GEN_10112 | _GEN_6587; // @[decode.scala 862:{68,68}]
  wire  _GEN_9491 = _GEN_10113 | _GEN_6588; // @[decode.scala 862:{68,68}]
  wire  _GEN_9492 = _GEN_10114 | _GEN_6589; // @[decode.scala 862:{68,68}]
  wire  _GEN_9493 = _GEN_10115 | _GEN_6590; // @[decode.scala 862:{68,68}]
  wire  _GEN_9494 = _GEN_10116 | _GEN_6591; // @[decode.scala 862:{68,68}]
  wire  _GEN_9495 = _GEN_10117 | _GEN_6592; // @[decode.scala 862:{68,68}]
  wire  _GEN_9496 = _GEN_10118 | _GEN_6593; // @[decode.scala 862:{68,68}]
  wire  _GEN_9497 = _GEN_10119 | _GEN_6594; // @[decode.scala 862:{68,68}]
  wire  _GEN_9498 = _GEN_10120 | _GEN_6595; // @[decode.scala 862:{68,68}]
  wire  _GEN_9499 = _GEN_10121 | _GEN_6596; // @[decode.scala 862:{68,68}]
  wire  _GEN_9500 = _GEN_10122 | _GEN_6597; // @[decode.scala 862:{68,68}]
  wire  _GEN_9501 = _GEN_10123 | _GEN_6598; // @[decode.scala 862:{68,68}]
  wire  _GEN_9502 = _GEN_10124 | _GEN_6599; // @[decode.scala 862:{68,68}]
  wire  _GEN_9503 = _GEN_10125 | _GEN_6600; // @[decode.scala 862:{68,68}]
  wire  _GEN_9504 = _GEN_10126 | _GEN_6601; // @[decode.scala 862:{68,68}]
  wire  _GEN_9505 = _GEN_10127 | _GEN_6602; // @[decode.scala 862:{68,68}]
  wire  _GEN_9506 = _GEN_10128 | _GEN_6603; // @[decode.scala 862:{68,68}]
  wire  _GEN_9507 = _GEN_10129 | _GEN_6604; // @[decode.scala 862:{68,68}]
  wire  _GEN_9508 = _GEN_10130 | _GEN_6605; // @[decode.scala 862:{68,68}]
  wire  _GEN_9509 = _GEN_10131 | _GEN_6606; // @[decode.scala 862:{68,68}]
  wire  _GEN_9510 = _GEN_10132 | _GEN_6607; // @[decode.scala 862:{68,68}]
  wire  _GEN_9511 = _GEN_10133 | _GEN_6608; // @[decode.scala 862:{68,68}]
  wire  _GEN_9512 = _GEN_10134 | _GEN_6609; // @[decode.scala 862:{68,68}]
  wire  _GEN_9513 = _GEN_10135 | _GEN_6610; // @[decode.scala 862:{68,68}]
  wire  _GEN_9514 = _GEN_10136 | _GEN_6611; // @[decode.scala 862:{68,68}]
  wire  _GEN_9515 = _GEN_10137 | _GEN_6612; // @[decode.scala 862:{68,68}]
  wire  _GEN_9516 = _GEN_10138 | _GEN_6613; // @[decode.scala 862:{68,68}]
  wire  _GEN_9582 = _T_464 ? _GEN_9230 : _GEN_1920; // @[decode.scala 856:5]
  wire  _GEN_9583 = _T_464 ? _GEN_9231 : _GEN_1921; // @[decode.scala 856:5]
  wire  _GEN_9584 = _T_464 ? _GEN_9232 : _GEN_1922; // @[decode.scala 856:5]
  wire  _GEN_9585 = _T_464 ? _GEN_9233 : _GEN_1923; // @[decode.scala 856:5]
  wire  _GEN_9586 = _T_464 ? _GEN_9234 : _GEN_1924; // @[decode.scala 856:5]
  wire  _GEN_9587 = _T_464 ? _GEN_9235 : _GEN_1925; // @[decode.scala 856:5]
  wire  _GEN_9588 = _T_464 ? _GEN_9236 : _GEN_1926; // @[decode.scala 856:5]
  wire  _GEN_9589 = _T_464 ? _GEN_9237 : _GEN_1927; // @[decode.scala 856:5]
  wire  _GEN_9590 = _T_464 ? _GEN_9238 : _GEN_1928; // @[decode.scala 856:5]
  wire  _GEN_9591 = _T_464 ? _GEN_9239 : _GEN_1929; // @[decode.scala 856:5]
  wire  _GEN_9592 = _T_464 ? _GEN_9240 : _GEN_1930; // @[decode.scala 856:5]
  wire  _GEN_9593 = _T_464 ? _GEN_9241 : _GEN_1931; // @[decode.scala 856:5]
  wire  _GEN_9594 = _T_464 ? _GEN_9242 : _GEN_1932; // @[decode.scala 856:5]
  wire  _GEN_9595 = _T_464 ? _GEN_9243 : _GEN_1933; // @[decode.scala 856:5]
  wire  _GEN_9596 = _T_464 ? _GEN_9244 : _GEN_1934; // @[decode.scala 856:5]
  wire  _GEN_9597 = _T_464 ? _GEN_9245 : _GEN_1935; // @[decode.scala 856:5]
  wire  _GEN_9598 = _T_464 ? _GEN_9246 : _GEN_1936; // @[decode.scala 856:5]
  wire  _GEN_9599 = _T_464 ? _GEN_9247 : _GEN_1937; // @[decode.scala 856:5]
  wire  _GEN_9600 = _T_464 ? _GEN_9248 : _GEN_1938; // @[decode.scala 856:5]
  wire  _GEN_9601 = _T_464 ? _GEN_9249 : _GEN_1939; // @[decode.scala 856:5]
  wire  _GEN_9602 = _T_464 ? _GEN_9250 : _GEN_1940; // @[decode.scala 856:5]
  wire  _GEN_9603 = _T_464 ? _GEN_9251 : _GEN_1941; // @[decode.scala 856:5]
  wire  _GEN_9604 = _T_464 ? _GEN_9252 : _GEN_1942; // @[decode.scala 856:5]
  wire  _GEN_9605 = _T_464 ? _GEN_9253 : _GEN_1943; // @[decode.scala 856:5]
  wire  _GEN_9606 = _T_464 ? _GEN_9254 : _GEN_1944; // @[decode.scala 856:5]
  wire  _GEN_9607 = _T_464 ? _GEN_9255 : _GEN_1945; // @[decode.scala 856:5]
  wire  _GEN_9608 = _T_464 ? _GEN_9256 : _GEN_1946; // @[decode.scala 856:5]
  wire  _GEN_9609 = _T_464 ? _GEN_9257 : _GEN_1947; // @[decode.scala 856:5]
  wire  _GEN_9610 = _T_464 ? _GEN_9258 : _GEN_1948; // @[decode.scala 856:5]
  wire  _GEN_9611 = _T_464 ? _GEN_9259 : _GEN_1949; // @[decode.scala 856:5]
  wire  _GEN_9612 = _T_464 ? _GEN_9260 : _GEN_1950; // @[decode.scala 856:5]
  wire  _GEN_9870 = currentPrivilege == 64'h2200001800 ? mie[7] : mstatus[3] & mie[7]; // @[decode.scala 870:44 872:22 875:22]
  wire [63:0] _GEN_10391 = reset ? 64'h0 : _GEN_6686; // @[decode.scala 236:{27,27}]
  wire [126:0] _GEN_10392 = reset ? 127'h0 : _GEN_8667; // @[decode.scala 471:{28,28}]
  assign fromFetch_ready = ~stateRegInputBuf ? _GEN_9098 : stateRegInputBuf & _GEN_9109; // @[decode.scala 759:28]
  assign fromFetch_expected_valid = expectedPC != 64'h0; // @[decode.scala 255:42]
  assign fromFetch_expected_pc = expectedPC; // @[decode.scala 256:28]
  assign toExec_ready = ~stateRegOutputBuf ? 1'h0 : stateRegOutputBuf & _GEN_9096; // @[decode.scala 813:29]
  assign toExec_instruction = outputBuffer_instruction; // @[decode.scala 244:22]
  assign toExec_pc = outputBuffer_pc; // @[decode.scala 245:22]
  assign toExec_PRFDest = outputBuffer_PRFDest; // @[decode.scala 246:22]
  assign toExec_rs1Addr = outputBuffer_rs1Addr; // @[decode.scala 247:22]
  assign toExec_rs1Ready = 6'h3f == outputBuffer_rs1Addr ? PRFValidList_63 : _GEN_74; // @[decode.scala 248:{22,22}]
  assign toExec_rs2Addr = outputBuffer_rs2Addr; // @[decode.scala 249:22]
  assign toExec_rs2Ready = _GEN_181 | (3'h1 == toExec_rs2Ready_insType | 3'h4 == toExec_rs2Ready_insType | 3'h5 ==
    toExec_rs2Ready_insType); // @[decode.scala 250:60]
  assign toExec_branchMask = {toExec_branchMask_hi,toExec_branchMask_lo}; // @[decode.scala 252:49]
  assign jumpAddrWrite_ready = validOutputBuf & (unconditionalJumps | csrIns); // @[decode.scala 258:44]
  assign jumpAddrWrite_PRFDest = outputBuffer_PRFDest; // @[decode.scala 259:26]
  assign jumpAddrWrite_linkAddr = unconditionalJumps ? _GEN_185 : csrReadDataReg; // @[decode.scala 260:28 261:28 267:28]
  assign branchPCs_branchPCReady = branchBuffer_branchPCReady; // @[decode.scala 272:30]
  assign branchPCs_branchPC = branchBuffer_branchPC; // @[decode.scala 274:30]
  assign branchPCs_predictedPCReady = branchBuffer_predictedPCReady; // @[decode.scala 273:30]
  assign branchPCs_predictedPC = branchBuffer_predictedPC; // @[decode.scala 275:30]
  assign branchPCs_branchMask = branchPCMask; // @[decode.scala 276:30]
  assign canTakeInterrupt = stallReg ? 1'h0 : _GEN_9870; // @[decode.scala 866:18 869:22]
  always @(posedge clock) begin
    if (reset) begin // @[decode.scala 107:28]
      inputBuffer_pc <= 64'hffffffc; // @[decode.scala 107:28]
    end else if (fromFetch_fired & readyInputBuf) begin // @[decode.scala 196:42]
      inputBuffer_pc <= fromFetch_pc; // @[decode.scala 198:29]
    end
    if (reset) begin // @[decode.scala 107:28]
      inputBuffer_instruction <= 32'h0; // @[decode.scala 107:28]
    end else if (fromFetch_fired & readyInputBuf) begin // @[decode.scala 196:42]
      inputBuffer_instruction <= fromFetch_instruction; // @[decode.scala 197:29]
    end
    if (reset) begin // @[decode.scala 116:29]
      outputBuffer_instruction <= 32'h0; // @[decode.scala 116:29]
    end else if (validInputBuf & readyOutputBuf) begin // @[decode.scala 206:41]
      outputBuffer_instruction <= inputBuffer_instruction; // @[decode.scala 207:30]
    end
    if (reset) begin // @[decode.scala 116:29]
      outputBuffer_pc <= 64'h0; // @[decode.scala 116:29]
    end else if (validInputBuf & readyOutputBuf) begin // @[decode.scala 206:41]
      outputBuffer_pc <= inputBuffer_pc; // @[decode.scala 208:30]
    end
    if (reset) begin // @[decode.scala 116:29]
      outputBuffer_PRFDest <= 6'h0; // @[decode.scala 116:29]
    end else if (validInputBuf & readyOutputBuf) begin // @[decode.scala 206:41]
      if (PRFFreeList_0) begin // @[Mux.scala 47:70]
        outputBuffer_PRFDest <= 6'h0;
      end else if (PRFFreeList_1) begin // @[Mux.scala 47:70]
        outputBuffer_PRFDest <= 6'h1;
      end else begin
        outputBuffer_PRFDest <= _freeRegAddr_T_60;
      end
    end
    if (reset) begin // @[decode.scala 116:29]
      outputBuffer_rs1Addr <= 6'h0; // @[decode.scala 116:29]
    end else if (validInputBuf & readyOutputBuf) begin // @[decode.scala 206:41]
      if (5'h1f == rs1) begin // @[decode.scala 325:12]
        outputBuffer_rs1Addr <= frontEndRegMap_31; // @[decode.scala 325:12]
      end else if (5'h1e == rs1) begin // @[decode.scala 325:12]
        outputBuffer_rs1Addr <= frontEndRegMap_30; // @[decode.scala 325:12]
      end else begin
        outputBuffer_rs1Addr <= _GEN_237;
      end
    end
    if (reset) begin // @[decode.scala 116:29]
      outputBuffer_rs2Addr <= 6'h0; // @[decode.scala 116:29]
    end else if (validInputBuf & readyOutputBuf) begin // @[decode.scala 206:41]
      if (5'h1f == rs2) begin // @[decode.scala 326:12]
        outputBuffer_rs2Addr <= frontEndRegMap_31; // @[decode.scala 326:12]
      end else if (5'h1e == rs2) begin // @[decode.scala 326:12]
        outputBuffer_rs2Addr <= frontEndRegMap_30; // @[decode.scala 326:12]
      end else begin
        outputBuffer_rs2Addr <= _GEN_269;
      end
    end
    if (reset) begin // @[decode.scala 116:29]
      outputBuffer_immediate <= 64'h0; // @[decode.scala 116:29]
    end else if (validInputBuf & readyOutputBuf) begin // @[decode.scala 206:41]
      outputBuffer_immediate <= immediate_immediate; // @[decode.scala 212:30]
    end
    if (reset) begin // @[decode.scala 138:29]
      branchBuffer_branchPCReady <= 1'h0; // @[decode.scala 138:29]
    end else begin
      branchBuffer_branchPCReady <= _T_435 & validInputBuf & readyOutputBuf; // @[decode.scala 452:30]
    end
    if (reset) begin // @[decode.scala 138:29]
      branchBuffer_predictedPCReady <= 1'h0; // @[decode.scala 138:29]
    end else begin
      branchBuffer_predictedPCReady <= branchReg & validInputBuf & readyOutputBuf; // @[decode.scala 453:33]
    end
    if (reset) begin // @[decode.scala 138:29]
      branchBuffer_branchPC <= 64'h0; // @[decode.scala 138:29]
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        branchBuffer_branchPC <= inputBuffer_pc; // @[decode.scala 391:29]
      end
    end
    if (reset) begin // @[decode.scala 138:29]
      branchBuffer_predictedPC <= 64'h0; // @[decode.scala 138:29]
    end else if (_toExec_branchMask_T != 4'h0 & validInputBuf & readyOutputBuf) begin // @[decode.scala 448:83]
      branchBuffer_predictedPC <= inputBuffer_pc; // @[decode.scala 449:30]
    end
    if (reset) begin // @[decode.scala 138:29]
      branchBuffer_branchMask_0 <= 1'h0; // @[decode.scala 138:29]
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        branchBuffer_branchMask_0 <= _GEN_2496;
      end else begin
        branchBuffer_branchMask_0 <= _GEN_1850;
      end
    end else begin
      branchBuffer_branchMask_0 <= _GEN_1850;
    end
    if (reset) begin // @[decode.scala 138:29]
      branchBuffer_branchMask_1 <= 1'h0; // @[decode.scala 138:29]
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        branchBuffer_branchMask_1 <= _GEN_2497;
      end else begin
        branchBuffer_branchMask_1 <= _GEN_1851;
      end
    end else begin
      branchBuffer_branchMask_1 <= _GEN_1851;
    end
    if (reset) begin // @[decode.scala 138:29]
      branchBuffer_branchMask_2 <= 1'h0; // @[decode.scala 138:29]
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        branchBuffer_branchMask_2 <= _GEN_2498;
      end else begin
        branchBuffer_branchMask_2 <= _GEN_1852;
      end
    end else begin
      branchBuffer_branchMask_2 <= _GEN_1852;
    end
    if (reset) begin // @[decode.scala 138:29]
      branchBuffer_branchMask_3 <= 1'h0; // @[decode.scala 138:29]
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        branchBuffer_branchMask_3 <= _GEN_2499;
      end else begin
        branchBuffer_branchMask_3 <= _GEN_1853;
      end
    end else begin
      branchBuffer_branchMask_3 <= _GEN_1853;
    end
    if (reset) begin // @[decode.scala 173:30]
      branchTracker <= 3'h0; // @[decode.scala 173:30]
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        branchTracker <= _branchTracker_T_3; // @[decode.scala 442:21]
      end else begin
        branchTracker <= _GEN_1849;
      end
    end else begin
      branchTracker <= _GEN_1849;
    end
    if (reset) begin // @[decode.scala 183:27]
      expectedPC <= 64'h10000000; // @[decode.scala 183:27]
    end else if (_T_246 & writeBackResult_instruction[14:12] == 3'h0) begin // @[decode.scala 711:126]
      if (writeBackResult_instruction[31:20] == 12'h302) begin // @[decode.scala 712:60]
        expectedPC <= mepc; // @[decode.scala 715:18]
      end else if (~(|writeBackResult_instruction[31:20])) begin // @[decode.scala 717:58]
        expectedPC <= mtvec; // @[decode.scala 723:18]
      end else begin
        expectedPC <= _GEN_8690;
      end
    end else if (_fromFetch_expected_valid_T & fromFetch_fired & fromFetch_expected_pc == fromFetch_pc) begin // @[decode.scala 455:89]
      expectedPC <= 64'h0; // @[decode.scala 456:16]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      expectedPC <= _GEN_1207;
    end
    if (reset) begin // @[decode.scala 187:34]
      stateRegInputBuf <= 1'h0; // @[decode.scala 187:34]
    end else if (~stateRegInputBuf) begin // @[decode.scala 759:28]
      if (branchEvalIn_fired & ~branchEvalIn_passFail) begin // @[decode.scala 761:58]
        stateRegInputBuf <= 1'h0; // @[decode.scala 762:26]
      end else if (fromFetch_fired) begin // @[decode.scala 769:31]
        stateRegInputBuf <= _GEN_9092;
      end
    end else if (stateRegInputBuf) begin // @[decode.scala 759:28]
      if (_T_425) begin // @[decode.scala 784:58]
        stateRegInputBuf <= 1'h0; // @[decode.scala 785:26]
      end else begin
        stateRegInputBuf <= _GEN_9104;
      end
    end
    if (reset) begin // @[decode.scala 188:34]
      stateRegOutputBuf <= 1'h0; // @[decode.scala 188:34]
    end else if (~stateRegOutputBuf) begin // @[decode.scala 813:29]
      if (_T_425) begin // @[decode.scala 815:58]
        stateRegOutputBuf <= 1'h0; // @[decode.scala 816:27]
      end else begin
        stateRegOutputBuf <= _GEN_9118;
      end
    end else if (stateRegOutputBuf) begin // @[decode.scala 813:29]
      if (_T_425) begin // @[decode.scala 828:58]
        stateRegOutputBuf <= 1'h0; // @[decode.scala 829:27]
      end else begin
        stateRegOutputBuf <= _GEN_9124;
      end
    end
    if (reset) begin // @[decode.scala 190:25]
      stallReg <= 1'h0; // @[decode.scala 190:25]
    end else if (~stateRegInputBuf) begin // @[decode.scala 759:28]
      stallReg <= _GEN_9097;
    end else if (stateRegInputBuf) begin // @[decode.scala 759:28]
      stallReg <= _GEN_9097;
    end else begin
      stallReg <= _GEN_6714;
    end
    if (fromFetch_fired & readyInputBuf) begin // @[decode.scala 196:42]
      if (fromFetch_instruction[6:0] == 7'h73) begin // @[decode.scala 199:97]
        ecallPC <= fromFetch_pc; // @[decode.scala 201:15]
      end
    end
    PRFValidList_0 <= reset | _GEN_9027; // @[decode.scala 193:{29,29}]
    PRFValidList_1 <= reset | _GEN_9028; // @[decode.scala 193:{29,29}]
    PRFValidList_2 <= reset | _GEN_9029; // @[decode.scala 193:{29,29}]
    PRFValidList_3 <= reset | _GEN_9030; // @[decode.scala 193:{29,29}]
    PRFValidList_4 <= reset | _GEN_9031; // @[decode.scala 193:{29,29}]
    PRFValidList_5 <= reset | _GEN_9032; // @[decode.scala 193:{29,29}]
    PRFValidList_6 <= reset | _GEN_9033; // @[decode.scala 193:{29,29}]
    PRFValidList_7 <= reset | _GEN_9034; // @[decode.scala 193:{29,29}]
    PRFValidList_8 <= reset | _GEN_9035; // @[decode.scala 193:{29,29}]
    PRFValidList_9 <= reset | _GEN_9036; // @[decode.scala 193:{29,29}]
    PRFValidList_10 <= reset | _GEN_9037; // @[decode.scala 193:{29,29}]
    PRFValidList_11 <= reset | _GEN_9038; // @[decode.scala 193:{29,29}]
    PRFValidList_12 <= reset | _GEN_9039; // @[decode.scala 193:{29,29}]
    PRFValidList_13 <= reset | _GEN_9040; // @[decode.scala 193:{29,29}]
    PRFValidList_14 <= reset | _GEN_9041; // @[decode.scala 193:{29,29}]
    PRFValidList_15 <= reset | _GEN_9042; // @[decode.scala 193:{29,29}]
    PRFValidList_16 <= reset | _GEN_9043; // @[decode.scala 193:{29,29}]
    PRFValidList_17 <= reset | _GEN_9044; // @[decode.scala 193:{29,29}]
    PRFValidList_18 <= reset | _GEN_9045; // @[decode.scala 193:{29,29}]
    PRFValidList_19 <= reset | _GEN_9046; // @[decode.scala 193:{29,29}]
    PRFValidList_20 <= reset | _GEN_9047; // @[decode.scala 193:{29,29}]
    PRFValidList_21 <= reset | _GEN_9048; // @[decode.scala 193:{29,29}]
    PRFValidList_22 <= reset | _GEN_9049; // @[decode.scala 193:{29,29}]
    PRFValidList_23 <= reset | _GEN_9050; // @[decode.scala 193:{29,29}]
    PRFValidList_24 <= reset | _GEN_9051; // @[decode.scala 193:{29,29}]
    PRFValidList_25 <= reset | _GEN_9052; // @[decode.scala 193:{29,29}]
    PRFValidList_26 <= reset | _GEN_9053; // @[decode.scala 193:{29,29}]
    PRFValidList_27 <= reset | _GEN_9054; // @[decode.scala 193:{29,29}]
    PRFValidList_28 <= reset | _GEN_9055; // @[decode.scala 193:{29,29}]
    PRFValidList_29 <= reset | _GEN_9056; // @[decode.scala 193:{29,29}]
    PRFValidList_30 <= reset | _GEN_9057; // @[decode.scala 193:{29,29}]
    PRFValidList_31 <= reset | _GEN_9058; // @[decode.scala 193:{29,29}]
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_32 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_32 <= 6'h20 == writeAddrPRF_exec3Addr | _GEN_8931;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_32 <= 6'h20 == writeAddrPRF_exec2Addr | _GEN_8803;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_32 <= 6'h20 == writeAddrPRF_exec1Addr | _GEN_1984;
    end else begin
      PRFValidList_32 <= _GEN_1984;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_33 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_33 <= 6'h21 == writeAddrPRF_exec3Addr | _GEN_8932;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_33 <= 6'h21 == writeAddrPRF_exec2Addr | _GEN_8804;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_33 <= 6'h21 == writeAddrPRF_exec1Addr | _GEN_1985;
    end else begin
      PRFValidList_33 <= _GEN_1985;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_34 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_34 <= 6'h22 == writeAddrPRF_exec3Addr | _GEN_8933;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_34 <= 6'h22 == writeAddrPRF_exec2Addr | _GEN_8805;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_34 <= 6'h22 == writeAddrPRF_exec1Addr | _GEN_1986;
    end else begin
      PRFValidList_34 <= _GEN_1986;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_35 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_35 <= 6'h23 == writeAddrPRF_exec3Addr | _GEN_8934;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_35 <= 6'h23 == writeAddrPRF_exec2Addr | _GEN_8806;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_35 <= 6'h23 == writeAddrPRF_exec1Addr | _GEN_1987;
    end else begin
      PRFValidList_35 <= _GEN_1987;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_36 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_36 <= 6'h24 == writeAddrPRF_exec3Addr | _GEN_8935;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_36 <= 6'h24 == writeAddrPRF_exec2Addr | _GEN_8807;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_36 <= 6'h24 == writeAddrPRF_exec1Addr | _GEN_1988;
    end else begin
      PRFValidList_36 <= _GEN_1988;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_37 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_37 <= 6'h25 == writeAddrPRF_exec3Addr | _GEN_8936;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_37 <= 6'h25 == writeAddrPRF_exec2Addr | _GEN_8808;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_37 <= 6'h25 == writeAddrPRF_exec1Addr | _GEN_1989;
    end else begin
      PRFValidList_37 <= _GEN_1989;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_38 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_38 <= 6'h26 == writeAddrPRF_exec3Addr | _GEN_8937;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_38 <= 6'h26 == writeAddrPRF_exec2Addr | _GEN_8809;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_38 <= 6'h26 == writeAddrPRF_exec1Addr | _GEN_1990;
    end else begin
      PRFValidList_38 <= _GEN_1990;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_39 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_39 <= 6'h27 == writeAddrPRF_exec3Addr | _GEN_8938;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_39 <= 6'h27 == writeAddrPRF_exec2Addr | _GEN_8810;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_39 <= 6'h27 == writeAddrPRF_exec1Addr | _GEN_1991;
    end else begin
      PRFValidList_39 <= _GEN_1991;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_40 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_40 <= 6'h28 == writeAddrPRF_exec3Addr | _GEN_8939;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_40 <= 6'h28 == writeAddrPRF_exec2Addr | _GEN_8811;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_40 <= 6'h28 == writeAddrPRF_exec1Addr | _GEN_1992;
    end else begin
      PRFValidList_40 <= _GEN_1992;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_41 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_41 <= 6'h29 == writeAddrPRF_exec3Addr | _GEN_8940;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_41 <= 6'h29 == writeAddrPRF_exec2Addr | _GEN_8812;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_41 <= 6'h29 == writeAddrPRF_exec1Addr | _GEN_1993;
    end else begin
      PRFValidList_41 <= _GEN_1993;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_42 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_42 <= 6'h2a == writeAddrPRF_exec3Addr | _GEN_8941;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_42 <= 6'h2a == writeAddrPRF_exec2Addr | _GEN_8813;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_42 <= 6'h2a == writeAddrPRF_exec1Addr | _GEN_1994;
    end else begin
      PRFValidList_42 <= _GEN_1994;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_43 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_43 <= 6'h2b == writeAddrPRF_exec3Addr | _GEN_8942;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_43 <= 6'h2b == writeAddrPRF_exec2Addr | _GEN_8814;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_43 <= 6'h2b == writeAddrPRF_exec1Addr | _GEN_1995;
    end else begin
      PRFValidList_43 <= _GEN_1995;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_44 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_44 <= 6'h2c == writeAddrPRF_exec3Addr | _GEN_8943;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_44 <= 6'h2c == writeAddrPRF_exec2Addr | _GEN_8815;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_44 <= 6'h2c == writeAddrPRF_exec1Addr | _GEN_1996;
    end else begin
      PRFValidList_44 <= _GEN_1996;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_45 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_45 <= 6'h2d == writeAddrPRF_exec3Addr | _GEN_8944;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_45 <= 6'h2d == writeAddrPRF_exec2Addr | _GEN_8816;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_45 <= 6'h2d == writeAddrPRF_exec1Addr | _GEN_1997;
    end else begin
      PRFValidList_45 <= _GEN_1997;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_46 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_46 <= 6'h2e == writeAddrPRF_exec3Addr | _GEN_8945;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_46 <= 6'h2e == writeAddrPRF_exec2Addr | _GEN_8817;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_46 <= 6'h2e == writeAddrPRF_exec1Addr | _GEN_1998;
    end else begin
      PRFValidList_46 <= _GEN_1998;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_47 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_47 <= 6'h2f == writeAddrPRF_exec3Addr | _GEN_8946;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_47 <= 6'h2f == writeAddrPRF_exec2Addr | _GEN_8818;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_47 <= 6'h2f == writeAddrPRF_exec1Addr | _GEN_1999;
    end else begin
      PRFValidList_47 <= _GEN_1999;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_48 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_48 <= 6'h30 == writeAddrPRF_exec3Addr | _GEN_8947;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_48 <= 6'h30 == writeAddrPRF_exec2Addr | _GEN_8819;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_48 <= 6'h30 == writeAddrPRF_exec1Addr | _GEN_2000;
    end else begin
      PRFValidList_48 <= _GEN_2000;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_49 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_49 <= 6'h31 == writeAddrPRF_exec3Addr | _GEN_8948;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_49 <= 6'h31 == writeAddrPRF_exec2Addr | _GEN_8820;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_49 <= 6'h31 == writeAddrPRF_exec1Addr | _GEN_2001;
    end else begin
      PRFValidList_49 <= _GEN_2001;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_50 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_50 <= 6'h32 == writeAddrPRF_exec3Addr | _GEN_8949;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_50 <= 6'h32 == writeAddrPRF_exec2Addr | _GEN_8821;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_50 <= 6'h32 == writeAddrPRF_exec1Addr | _GEN_2002;
    end else begin
      PRFValidList_50 <= _GEN_2002;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_51 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_51 <= 6'h33 == writeAddrPRF_exec3Addr | _GEN_8950;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_51 <= 6'h33 == writeAddrPRF_exec2Addr | _GEN_8822;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_51 <= 6'h33 == writeAddrPRF_exec1Addr | _GEN_2003;
    end else begin
      PRFValidList_51 <= _GEN_2003;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_52 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_52 <= 6'h34 == writeAddrPRF_exec3Addr | _GEN_8951;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_52 <= 6'h34 == writeAddrPRF_exec2Addr | _GEN_8823;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_52 <= 6'h34 == writeAddrPRF_exec1Addr | _GEN_2004;
    end else begin
      PRFValidList_52 <= _GEN_2004;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_53 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_53 <= 6'h35 == writeAddrPRF_exec3Addr | _GEN_8952;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_53 <= 6'h35 == writeAddrPRF_exec2Addr | _GEN_8824;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_53 <= 6'h35 == writeAddrPRF_exec1Addr | _GEN_2005;
    end else begin
      PRFValidList_53 <= _GEN_2005;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_54 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_54 <= 6'h36 == writeAddrPRF_exec3Addr | _GEN_8953;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_54 <= 6'h36 == writeAddrPRF_exec2Addr | _GEN_8825;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_54 <= 6'h36 == writeAddrPRF_exec1Addr | _GEN_2006;
    end else begin
      PRFValidList_54 <= _GEN_2006;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_55 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_55 <= 6'h37 == writeAddrPRF_exec3Addr | _GEN_8954;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_55 <= 6'h37 == writeAddrPRF_exec2Addr | _GEN_8826;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_55 <= 6'h37 == writeAddrPRF_exec1Addr | _GEN_2007;
    end else begin
      PRFValidList_55 <= _GEN_2007;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_56 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_56 <= 6'h38 == writeAddrPRF_exec3Addr | _GEN_8955;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_56 <= 6'h38 == writeAddrPRF_exec2Addr | _GEN_8827;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_56 <= 6'h38 == writeAddrPRF_exec1Addr | _GEN_2008;
    end else begin
      PRFValidList_56 <= _GEN_2008;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_57 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_57 <= 6'h39 == writeAddrPRF_exec3Addr | _GEN_8956;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_57 <= 6'h39 == writeAddrPRF_exec2Addr | _GEN_8828;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_57 <= 6'h39 == writeAddrPRF_exec1Addr | _GEN_2009;
    end else begin
      PRFValidList_57 <= _GEN_2009;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_58 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_58 <= 6'h3a == writeAddrPRF_exec3Addr | _GEN_8957;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_58 <= 6'h3a == writeAddrPRF_exec2Addr | _GEN_8829;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_58 <= 6'h3a == writeAddrPRF_exec1Addr | _GEN_2010;
    end else begin
      PRFValidList_58 <= _GEN_2010;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_59 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_59 <= 6'h3b == writeAddrPRF_exec3Addr | _GEN_8958;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_59 <= 6'h3b == writeAddrPRF_exec2Addr | _GEN_8830;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_59 <= 6'h3b == writeAddrPRF_exec1Addr | _GEN_2011;
    end else begin
      PRFValidList_59 <= _GEN_2011;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_60 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_60 <= 6'h3c == writeAddrPRF_exec3Addr | _GEN_8959;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_60 <= 6'h3c == writeAddrPRF_exec2Addr | _GEN_8831;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_60 <= 6'h3c == writeAddrPRF_exec1Addr | _GEN_2012;
    end else begin
      PRFValidList_60 <= _GEN_2012;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_61 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_61 <= 6'h3d == writeAddrPRF_exec3Addr | _GEN_8960;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_61 <= 6'h3d == writeAddrPRF_exec2Addr | _GEN_8832;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_61 <= 6'h3d == writeAddrPRF_exec1Addr | _GEN_2013;
    end else begin
      PRFValidList_61 <= _GEN_2013;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_62 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_62 <= 6'h3e == writeAddrPRF_exec3Addr | _GEN_8961;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_62 <= 6'h3e == writeAddrPRF_exec2Addr | _GEN_8833;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_62 <= 6'h3e == writeAddrPRF_exec1Addr | _GEN_2014;
    end else begin
      PRFValidList_62 <= _GEN_2014;
    end
    if (reset) begin // @[decode.scala 193:29]
      PRFValidList_63 <= 1'h0; // @[decode.scala 193:29]
    end else if (writeAddrPRF_exec3Valid) begin // @[decode.scala 753:33]
      PRFValidList_63 <= 6'h3f == writeAddrPRF_exec3Addr | _GEN_8962;
    end else if (writeAddrPRF_exec2Valid) begin // @[decode.scala 752:33]
      PRFValidList_63 <= 6'h3f == writeAddrPRF_exec2Addr | _GEN_8834;
    end else if (writeAddrPRF_exec1Valid) begin // @[decode.scala 751:33]
      PRFValidList_63 <= 6'h3f == writeAddrPRF_exec1Addr | _GEN_2015;
    end else begin
      PRFValidList_63 <= _GEN_2015;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_31 <= 6'h1f; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_31 <= reservedRegMap1_31; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_31 <= _GEN_1201;
      end
    end else begin
      frontEndRegMap_31 <= _GEN_1201;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_30 <= 6'h1e; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_30 <= reservedRegMap1_30; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_30 <= _GEN_1200;
      end
    end else begin
      frontEndRegMap_30 <= _GEN_1200;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_29 <= 6'h1d; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_29 <= reservedRegMap1_29; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_29 <= _GEN_1199;
      end
    end else begin
      frontEndRegMap_29 <= _GEN_1199;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_28 <= 6'h1c; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_28 <= reservedRegMap1_28; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_28 <= _GEN_1198;
      end
    end else begin
      frontEndRegMap_28 <= _GEN_1198;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_27 <= 6'h1b; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_27 <= reservedRegMap1_27; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_27 <= _GEN_1197;
      end
    end else begin
      frontEndRegMap_27 <= _GEN_1197;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_26 <= 6'h1a; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_26 <= reservedRegMap1_26; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_26 <= _GEN_1196;
      end
    end else begin
      frontEndRegMap_26 <= _GEN_1196;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_25 <= 6'h19; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_25 <= reservedRegMap1_25; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_25 <= _GEN_1195;
      end
    end else begin
      frontEndRegMap_25 <= _GEN_1195;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_24 <= 6'h18; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_24 <= reservedRegMap1_24; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_24 <= _GEN_1194;
      end
    end else begin
      frontEndRegMap_24 <= _GEN_1194;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_23 <= 6'h17; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_23 <= reservedRegMap1_23; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_23 <= _GEN_1193;
      end
    end else begin
      frontEndRegMap_23 <= _GEN_1193;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_22 <= 6'h16; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_22 <= reservedRegMap1_22; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_22 <= _GEN_1192;
      end
    end else begin
      frontEndRegMap_22 <= _GEN_1192;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_21 <= 6'h15; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_21 <= reservedRegMap1_21; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_21 <= _GEN_1191;
      end
    end else begin
      frontEndRegMap_21 <= _GEN_1191;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_20 <= 6'h14; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_20 <= reservedRegMap1_20; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_20 <= _GEN_1190;
      end
    end else begin
      frontEndRegMap_20 <= _GEN_1190;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_19 <= 6'h13; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_19 <= reservedRegMap1_19; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_19 <= _GEN_1189;
      end
    end else begin
      frontEndRegMap_19 <= _GEN_1189;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_18 <= 6'h12; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_18 <= reservedRegMap1_18; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_18 <= _GEN_1188;
      end
    end else begin
      frontEndRegMap_18 <= _GEN_1188;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_17 <= 6'h11; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_17 <= reservedRegMap1_17; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_17 <= _GEN_1187;
      end
    end else begin
      frontEndRegMap_17 <= _GEN_1187;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_16 <= 6'h10; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_16 <= reservedRegMap1_16; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_16 <= _GEN_1186;
      end
    end else begin
      frontEndRegMap_16 <= _GEN_1186;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_15 <= 6'hf; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_15 <= reservedRegMap1_15; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_15 <= _GEN_1185;
      end
    end else begin
      frontEndRegMap_15 <= _GEN_1185;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_14 <= 6'he; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_14 <= reservedRegMap1_14; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_14 <= _GEN_1184;
      end
    end else begin
      frontEndRegMap_14 <= _GEN_1184;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_13 <= 6'hd; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_13 <= reservedRegMap1_13; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_13 <= _GEN_1183;
      end
    end else begin
      frontEndRegMap_13 <= _GEN_1183;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_12 <= 6'hc; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_12 <= reservedRegMap1_12; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_12 <= _GEN_1182;
      end
    end else begin
      frontEndRegMap_12 <= _GEN_1182;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_11 <= 6'hb; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_11 <= reservedRegMap1_11; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_11 <= _GEN_1181;
      end
    end else begin
      frontEndRegMap_11 <= _GEN_1181;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_10 <= 6'ha; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_10 <= reservedRegMap1_10; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_10 <= _GEN_1180;
      end
    end else begin
      frontEndRegMap_10 <= _GEN_1180;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_9 <= 6'h9; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_9 <= reservedRegMap1_9; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_9 <= _GEN_1179;
      end
    end else begin
      frontEndRegMap_9 <= _GEN_1179;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_8 <= 6'h8; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_8 <= reservedRegMap1_8; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_8 <= _GEN_1178;
      end
    end else begin
      frontEndRegMap_8 <= _GEN_1178;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_7 <= 6'h7; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_7 <= reservedRegMap1_7; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_7 <= _GEN_1177;
      end
    end else begin
      frontEndRegMap_7 <= _GEN_1177;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_6 <= 6'h6; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_6 <= reservedRegMap1_6; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_6 <= _GEN_1176;
      end
    end else begin
      frontEndRegMap_6 <= _GEN_1176;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_5 <= 6'h5; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_5 <= reservedRegMap1_5; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_5 <= _GEN_1175;
      end
    end else begin
      frontEndRegMap_5 <= _GEN_1175;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_4 <= 6'h4; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_4 <= reservedRegMap1_4; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_4 <= _GEN_1174;
      end
    end else begin
      frontEndRegMap_4 <= _GEN_1174;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_3 <= 6'h3; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_3 <= reservedRegMap1_3; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_3 <= _GEN_1173;
      end
    end else begin
      frontEndRegMap_3 <= _GEN_1173;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_2 <= 6'h2; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_2 <= reservedRegMap1_2; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_2 <= _GEN_1172;
      end
    end else begin
      frontEndRegMap_2 <= _GEN_1172;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_1 <= 6'h1; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_1 <= reservedRegMap1_1; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_1 <= _GEN_1171;
      end
    end else begin
      frontEndRegMap_1 <= _GEN_1171;
    end
    if (reset) begin // @[decode.scala 301:36]
      frontEndRegMap_0 <= 6'h0; // @[decode.scala 301:36]
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        frontEndRegMap_0 <= reservedRegMap1_0; // @[decode.scala 365:22]
      end else begin
        frontEndRegMap_0 <= _GEN_1170;
      end
    end else begin
      frontEndRegMap_0 <= _GEN_1170;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_0 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_0 <= _GEN_9198;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_0 <= reservedFreeList1_0 | PRFFreeList_0; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_0 <= _GEN_1042;
      end
    end else begin
      PRFFreeList_0 <= _GEN_1042;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_1 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_1 <= _GEN_9199;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_1 <= reservedFreeList1_1 | PRFFreeList_1; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_1 <= _GEN_1043;
      end
    end else begin
      PRFFreeList_1 <= _GEN_1043;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_2 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_2 <= _GEN_9200;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_2 <= reservedFreeList1_2 | PRFFreeList_2; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_2 <= _GEN_1044;
      end
    end else begin
      PRFFreeList_2 <= _GEN_1044;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_3 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_3 <= _GEN_9201;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_3 <= reservedFreeList1_3 | PRFFreeList_3; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_3 <= _GEN_1045;
      end
    end else begin
      PRFFreeList_3 <= _GEN_1045;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_4 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_4 <= _GEN_9202;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_4 <= reservedFreeList1_4 | PRFFreeList_4; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_4 <= _GEN_1046;
      end
    end else begin
      PRFFreeList_4 <= _GEN_1046;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_5 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_5 <= _GEN_9203;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_5 <= reservedFreeList1_5 | PRFFreeList_5; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_5 <= _GEN_1047;
      end
    end else begin
      PRFFreeList_5 <= _GEN_1047;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_6 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_6 <= _GEN_9204;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_6 <= reservedFreeList1_6 | PRFFreeList_6; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_6 <= _GEN_1048;
      end
    end else begin
      PRFFreeList_6 <= _GEN_1048;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_7 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_7 <= _GEN_9205;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_7 <= reservedFreeList1_7 | PRFFreeList_7; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_7 <= _GEN_1049;
      end
    end else begin
      PRFFreeList_7 <= _GEN_1049;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_8 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_8 <= _GEN_9206;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_8 <= reservedFreeList1_8 | PRFFreeList_8; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_8 <= _GEN_1050;
      end
    end else begin
      PRFFreeList_8 <= _GEN_1050;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_9 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_9 <= _GEN_9207;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_9 <= reservedFreeList1_9 | PRFFreeList_9; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_9 <= _GEN_1051;
      end
    end else begin
      PRFFreeList_9 <= _GEN_1051;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_10 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_10 <= _GEN_9208;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_10 <= reservedFreeList1_10 | PRFFreeList_10; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_10 <= _GEN_1052;
      end
    end else begin
      PRFFreeList_10 <= _GEN_1052;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_11 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_11 <= _GEN_9209;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_11 <= reservedFreeList1_11 | PRFFreeList_11; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_11 <= _GEN_1053;
      end
    end else begin
      PRFFreeList_11 <= _GEN_1053;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_12 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_12 <= _GEN_9210;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_12 <= reservedFreeList1_12 | PRFFreeList_12; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_12 <= _GEN_1054;
      end
    end else begin
      PRFFreeList_12 <= _GEN_1054;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_13 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_13 <= _GEN_9211;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_13 <= reservedFreeList1_13 | PRFFreeList_13; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_13 <= _GEN_1055;
      end
    end else begin
      PRFFreeList_13 <= _GEN_1055;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_14 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_14 <= _GEN_9212;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_14 <= reservedFreeList1_14 | PRFFreeList_14; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_14 <= _GEN_1056;
      end
    end else begin
      PRFFreeList_14 <= _GEN_1056;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_15 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_15 <= _GEN_9213;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_15 <= reservedFreeList1_15 | PRFFreeList_15; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_15 <= _GEN_1057;
      end
    end else begin
      PRFFreeList_15 <= _GEN_1057;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_16 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_16 <= _GEN_9214;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_16 <= reservedFreeList1_16 | PRFFreeList_16; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_16 <= _GEN_1058;
      end
    end else begin
      PRFFreeList_16 <= _GEN_1058;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_17 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_17 <= _GEN_9215;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_17 <= reservedFreeList1_17 | PRFFreeList_17; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_17 <= _GEN_1059;
      end
    end else begin
      PRFFreeList_17 <= _GEN_1059;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_18 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_18 <= _GEN_9216;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_18 <= reservedFreeList1_18 | PRFFreeList_18; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_18 <= _GEN_1060;
      end
    end else begin
      PRFFreeList_18 <= _GEN_1060;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_19 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_19 <= _GEN_9217;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_19 <= reservedFreeList1_19 | PRFFreeList_19; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_19 <= _GEN_1061;
      end
    end else begin
      PRFFreeList_19 <= _GEN_1061;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_20 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_20 <= _GEN_9218;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_20 <= reservedFreeList1_20 | PRFFreeList_20; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_20 <= _GEN_1062;
      end
    end else begin
      PRFFreeList_20 <= _GEN_1062;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_21 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_21 <= _GEN_9219;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_21 <= reservedFreeList1_21 | PRFFreeList_21; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_21 <= _GEN_1063;
      end
    end else begin
      PRFFreeList_21 <= _GEN_1063;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_22 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_22 <= _GEN_9220;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_22 <= reservedFreeList1_22 | PRFFreeList_22; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_22 <= _GEN_1064;
      end
    end else begin
      PRFFreeList_22 <= _GEN_1064;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_23 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_23 <= _GEN_9221;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_23 <= reservedFreeList1_23 | PRFFreeList_23; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_23 <= _GEN_1065;
      end
    end else begin
      PRFFreeList_23 <= _GEN_1065;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_24 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_24 <= _GEN_9222;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_24 <= reservedFreeList1_24 | PRFFreeList_24; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_24 <= _GEN_1066;
      end
    end else begin
      PRFFreeList_24 <= _GEN_1066;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_25 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_25 <= _GEN_9223;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_25 <= reservedFreeList1_25 | PRFFreeList_25; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_25 <= _GEN_1067;
      end
    end else begin
      PRFFreeList_25 <= _GEN_1067;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_26 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_26 <= _GEN_9224;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_26 <= reservedFreeList1_26 | PRFFreeList_26; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_26 <= _GEN_1068;
      end
    end else begin
      PRFFreeList_26 <= _GEN_1068;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_27 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_27 <= _GEN_9225;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_27 <= reservedFreeList1_27 | PRFFreeList_27; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_27 <= _GEN_1069;
      end
    end else begin
      PRFFreeList_27 <= _GEN_1069;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_28 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_28 <= _GEN_9226;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_28 <= reservedFreeList1_28 | PRFFreeList_28; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_28 <= _GEN_1070;
      end
    end else begin
      PRFFreeList_28 <= _GEN_1070;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_29 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_29 <= _GEN_9227;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_29 <= reservedFreeList1_29 | PRFFreeList_29; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_29 <= _GEN_1071;
      end
    end else begin
      PRFFreeList_29 <= _GEN_1071;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_30 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_30 <= _GEN_9228;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_30 <= reservedFreeList1_30 | PRFFreeList_30; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_30 <= _GEN_1072;
      end
    end else begin
      PRFFreeList_30 <= _GEN_1072;
    end
    if (reset) begin // @[decode.scala 303:36]
      PRFFreeList_31 <= 1'h0; // @[decode.scala 303:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      PRFFreeList_31 <= _GEN_9229;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        PRFFreeList_31 <= reservedFreeList1_31 | PRFFreeList_31; // @[decode.scala 366:22]
      end else begin
        PRFFreeList_31 <= _GEN_1073;
      end
    end else begin
      PRFFreeList_31 <= _GEN_1073;
    end
    PRFFreeList_32 <= reset | _GEN_9582; // @[decode.scala 303:{36,36}]
    PRFFreeList_33 <= reset | _GEN_9583; // @[decode.scala 303:{36,36}]
    PRFFreeList_34 <= reset | _GEN_9584; // @[decode.scala 303:{36,36}]
    PRFFreeList_35 <= reset | _GEN_9585; // @[decode.scala 303:{36,36}]
    PRFFreeList_36 <= reset | _GEN_9586; // @[decode.scala 303:{36,36}]
    PRFFreeList_37 <= reset | _GEN_9587; // @[decode.scala 303:{36,36}]
    PRFFreeList_38 <= reset | _GEN_9588; // @[decode.scala 303:{36,36}]
    PRFFreeList_39 <= reset | _GEN_9589; // @[decode.scala 303:{36,36}]
    PRFFreeList_40 <= reset | _GEN_9590; // @[decode.scala 303:{36,36}]
    PRFFreeList_41 <= reset | _GEN_9591; // @[decode.scala 303:{36,36}]
    PRFFreeList_42 <= reset | _GEN_9592; // @[decode.scala 303:{36,36}]
    PRFFreeList_43 <= reset | _GEN_9593; // @[decode.scala 303:{36,36}]
    PRFFreeList_44 <= reset | _GEN_9594; // @[decode.scala 303:{36,36}]
    PRFFreeList_45 <= reset | _GEN_9595; // @[decode.scala 303:{36,36}]
    PRFFreeList_46 <= reset | _GEN_9596; // @[decode.scala 303:{36,36}]
    PRFFreeList_47 <= reset | _GEN_9597; // @[decode.scala 303:{36,36}]
    PRFFreeList_48 <= reset | _GEN_9598; // @[decode.scala 303:{36,36}]
    PRFFreeList_49 <= reset | _GEN_9599; // @[decode.scala 303:{36,36}]
    PRFFreeList_50 <= reset | _GEN_9600; // @[decode.scala 303:{36,36}]
    PRFFreeList_51 <= reset | _GEN_9601; // @[decode.scala 303:{36,36}]
    PRFFreeList_52 <= reset | _GEN_9602; // @[decode.scala 303:{36,36}]
    PRFFreeList_53 <= reset | _GEN_9603; // @[decode.scala 303:{36,36}]
    PRFFreeList_54 <= reset | _GEN_9604; // @[decode.scala 303:{36,36}]
    PRFFreeList_55 <= reset | _GEN_9605; // @[decode.scala 303:{36,36}]
    PRFFreeList_56 <= reset | _GEN_9606; // @[decode.scala 303:{36,36}]
    PRFFreeList_57 <= reset | _GEN_9607; // @[decode.scala 303:{36,36}]
    PRFFreeList_58 <= reset | _GEN_9608; // @[decode.scala 303:{36,36}]
    PRFFreeList_59 <= reset | _GEN_9609; // @[decode.scala 303:{36,36}]
    PRFFreeList_60 <= reset | _GEN_9610; // @[decode.scala 303:{36,36}]
    PRFFreeList_61 <= reset | _GEN_9611; // @[decode.scala 303:{36,36}]
    PRFFreeList_62 <= reset | _GEN_9612; // @[decode.scala 303:{36,36}]
    if (reset) begin // @[decode.scala 219:29]
      branchPCMask <= 4'h0; // @[decode.scala 219:29]
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (_GEN_9879) begin // @[decode.scala 393:27]
          branchPCMask <= 4'h1; // @[decode.scala 394:32]
        end else begin
          branchPCMask <= _GEN_2502;
        end
      end
    end
    if (reset) begin // @[decode.scala 220:29]
      branchReg <= 1'h0; // @[decode.scala 220:29]
    end else if (_T_3) begin // @[decode.scala 388:41]
      branchReg <= _T_181;
    end else if (branchEvalIn_fired) begin // @[decode.scala 352:28]
      if (_T_424) begin // @[decode.scala 356:34]
        branchReg <= 1'h0; // @[decode.scala 357:17]
      end
    end
    if (reset) begin // @[decode.scala 234:31]
      csrReadDataReg <= 64'h0; // @[decode.scala 234:31]
    end else if (opcode == 7'h73 & fun3 != 3'h0 & validInputBuf & readyOutputBuf) begin // @[decode.scala 501:80]
      if (64'h0 == _T_219) begin // @[decode.scala 502:34]
        csrReadDataReg <= ustatus; // @[decode.scala 503:37]
      end else if (64'h5 == _T_219) begin // @[decode.scala 502:34]
        csrReadDataReg <= utvec; // @[decode.scala 504:37]
      end else begin
        csrReadDataReg <= _GEN_6710;
      end
    end
    csrAddrReg <= _GEN_10391[11:0]; // @[decode.scala 236:{27,27}]
    if (reset) begin // @[decode.scala 237:26]
      csrImmReg <= 64'h0; // @[decode.scala 237:26]
    end else if (isCSR) begin // @[decode.scala 492:15]
      csrImmReg <= {{59'd0}, outputBuffer_instruction[19:15]}; // @[decode.scala 496:19]
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_0 <= 6'h0; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h0 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_0 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_1 <= 6'h1; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h1 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_1 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_2 <= 6'h2; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h2 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_2 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_3 <= 6'h3; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h3 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_3 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_4 <= 6'h4; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h4 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_4 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_5 <= 6'h5; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h5 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_5 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_6 <= 6'h6; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h6 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_6 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_7 <= 6'h7; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h7 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_7 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_8 <= 6'h8; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h8 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_8 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_9 <= 6'h9; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h9 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_9 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_10 <= 6'ha; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'ha == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_10 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_11 <= 6'hb; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'hb == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_11 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_12 <= 6'hc; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'hc == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_12 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_13 <= 6'hd; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'hd == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_13 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_14 <= 6'he; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'he == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_14 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_15 <= 6'hf; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'hf == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_15 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_16 <= 6'h10; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h10 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_16 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_17 <= 6'h11; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h11 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_17 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_18 <= 6'h12; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h12 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_18 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_19 <= 6'h13; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h13 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_19 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_20 <= 6'h14; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h14 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_20 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_21 <= 6'h15; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h15 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_21 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_22 <= 6'h16; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h16 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_22 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_23 <= 6'h17; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h17 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_23 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_24 <= 6'h18; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h18 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_24 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_25 <= 6'h19; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h19 == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_25 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_26 <= 6'h1a; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h1a == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_26 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_27 <= 6'h1b; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h1b == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_27 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_28 <= 6'h1c; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h1c == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_28 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_29 <= 6'h1d; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h1d == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_29 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_30 <= 6'h1e; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h1e == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_30 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (reset) begin // @[decode.scala 302:36]
      architecturalRegMap_31 <= 6'h1f; // @[decode.scala 302:36]
    end else if (_T_464) begin // @[decode.scala 856:5]
      if (5'h1f == writeBackResult_rdAddr) begin // @[decode.scala 857:62]
        architecturalRegMap_31 <= writeBackResult_PRFDest; // @[decode.scala 857:62]
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_0 <= _GEN_850;
          end else begin
            reservedRegMap1_0 <= frontEndRegMap_0; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_0 <= _GEN_2016;
        end
      end else begin
        reservedRegMap1_0 <= _GEN_2016;
      end
    end else begin
      reservedRegMap1_0 <= _GEN_2016;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_1 <= _GEN_851;
          end else begin
            reservedRegMap1_1 <= frontEndRegMap_1; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_1 <= _GEN_2017;
        end
      end else begin
        reservedRegMap1_1 <= _GEN_2017;
      end
    end else begin
      reservedRegMap1_1 <= _GEN_2017;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_2 <= _GEN_852;
          end else begin
            reservedRegMap1_2 <= frontEndRegMap_2; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_2 <= _GEN_2018;
        end
      end else begin
        reservedRegMap1_2 <= _GEN_2018;
      end
    end else begin
      reservedRegMap1_2 <= _GEN_2018;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_3 <= _GEN_853;
          end else begin
            reservedRegMap1_3 <= frontEndRegMap_3; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_3 <= _GEN_2019;
        end
      end else begin
        reservedRegMap1_3 <= _GEN_2019;
      end
    end else begin
      reservedRegMap1_3 <= _GEN_2019;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_4 <= _GEN_854;
          end else begin
            reservedRegMap1_4 <= frontEndRegMap_4; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_4 <= _GEN_2020;
        end
      end else begin
        reservedRegMap1_4 <= _GEN_2020;
      end
    end else begin
      reservedRegMap1_4 <= _GEN_2020;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_5 <= _GEN_855;
          end else begin
            reservedRegMap1_5 <= frontEndRegMap_5; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_5 <= _GEN_2021;
        end
      end else begin
        reservedRegMap1_5 <= _GEN_2021;
      end
    end else begin
      reservedRegMap1_5 <= _GEN_2021;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_6 <= _GEN_856;
          end else begin
            reservedRegMap1_6 <= frontEndRegMap_6; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_6 <= _GEN_2022;
        end
      end else begin
        reservedRegMap1_6 <= _GEN_2022;
      end
    end else begin
      reservedRegMap1_6 <= _GEN_2022;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_7 <= _GEN_857;
          end else begin
            reservedRegMap1_7 <= frontEndRegMap_7; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_7 <= _GEN_2023;
        end
      end else begin
        reservedRegMap1_7 <= _GEN_2023;
      end
    end else begin
      reservedRegMap1_7 <= _GEN_2023;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_8 <= _GEN_858;
          end else begin
            reservedRegMap1_8 <= frontEndRegMap_8; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_8 <= _GEN_2024;
        end
      end else begin
        reservedRegMap1_8 <= _GEN_2024;
      end
    end else begin
      reservedRegMap1_8 <= _GEN_2024;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_9 <= _GEN_859;
          end else begin
            reservedRegMap1_9 <= frontEndRegMap_9; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_9 <= _GEN_2025;
        end
      end else begin
        reservedRegMap1_9 <= _GEN_2025;
      end
    end else begin
      reservedRegMap1_9 <= _GEN_2025;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_10 <= _GEN_860;
          end else begin
            reservedRegMap1_10 <= frontEndRegMap_10; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_10 <= _GEN_2026;
        end
      end else begin
        reservedRegMap1_10 <= _GEN_2026;
      end
    end else begin
      reservedRegMap1_10 <= _GEN_2026;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_11 <= _GEN_861;
          end else begin
            reservedRegMap1_11 <= frontEndRegMap_11; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_11 <= _GEN_2027;
        end
      end else begin
        reservedRegMap1_11 <= _GEN_2027;
      end
    end else begin
      reservedRegMap1_11 <= _GEN_2027;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_12 <= _GEN_862;
          end else begin
            reservedRegMap1_12 <= frontEndRegMap_12; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_12 <= _GEN_2028;
        end
      end else begin
        reservedRegMap1_12 <= _GEN_2028;
      end
    end else begin
      reservedRegMap1_12 <= _GEN_2028;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_13 <= _GEN_863;
          end else begin
            reservedRegMap1_13 <= frontEndRegMap_13; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_13 <= _GEN_2029;
        end
      end else begin
        reservedRegMap1_13 <= _GEN_2029;
      end
    end else begin
      reservedRegMap1_13 <= _GEN_2029;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_14 <= _GEN_864;
          end else begin
            reservedRegMap1_14 <= frontEndRegMap_14; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_14 <= _GEN_2030;
        end
      end else begin
        reservedRegMap1_14 <= _GEN_2030;
      end
    end else begin
      reservedRegMap1_14 <= _GEN_2030;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_15 <= _GEN_865;
          end else begin
            reservedRegMap1_15 <= frontEndRegMap_15; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_15 <= _GEN_2031;
        end
      end else begin
        reservedRegMap1_15 <= _GEN_2031;
      end
    end else begin
      reservedRegMap1_15 <= _GEN_2031;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_16 <= _GEN_866;
          end else begin
            reservedRegMap1_16 <= frontEndRegMap_16; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_16 <= _GEN_2032;
        end
      end else begin
        reservedRegMap1_16 <= _GEN_2032;
      end
    end else begin
      reservedRegMap1_16 <= _GEN_2032;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_17 <= _GEN_867;
          end else begin
            reservedRegMap1_17 <= frontEndRegMap_17; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_17 <= _GEN_2033;
        end
      end else begin
        reservedRegMap1_17 <= _GEN_2033;
      end
    end else begin
      reservedRegMap1_17 <= _GEN_2033;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_18 <= _GEN_868;
          end else begin
            reservedRegMap1_18 <= frontEndRegMap_18; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_18 <= _GEN_2034;
        end
      end else begin
        reservedRegMap1_18 <= _GEN_2034;
      end
    end else begin
      reservedRegMap1_18 <= _GEN_2034;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_19 <= _GEN_869;
          end else begin
            reservedRegMap1_19 <= frontEndRegMap_19; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_19 <= _GEN_2035;
        end
      end else begin
        reservedRegMap1_19 <= _GEN_2035;
      end
    end else begin
      reservedRegMap1_19 <= _GEN_2035;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_20 <= _GEN_870;
          end else begin
            reservedRegMap1_20 <= frontEndRegMap_20; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_20 <= _GEN_2036;
        end
      end else begin
        reservedRegMap1_20 <= _GEN_2036;
      end
    end else begin
      reservedRegMap1_20 <= _GEN_2036;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_21 <= _GEN_871;
          end else begin
            reservedRegMap1_21 <= frontEndRegMap_21; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_21 <= _GEN_2037;
        end
      end else begin
        reservedRegMap1_21 <= _GEN_2037;
      end
    end else begin
      reservedRegMap1_21 <= _GEN_2037;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_22 <= _GEN_872;
          end else begin
            reservedRegMap1_22 <= frontEndRegMap_22; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_22 <= _GEN_2038;
        end
      end else begin
        reservedRegMap1_22 <= _GEN_2038;
      end
    end else begin
      reservedRegMap1_22 <= _GEN_2038;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_23 <= _GEN_873;
          end else begin
            reservedRegMap1_23 <= frontEndRegMap_23; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_23 <= _GEN_2039;
        end
      end else begin
        reservedRegMap1_23 <= _GEN_2039;
      end
    end else begin
      reservedRegMap1_23 <= _GEN_2039;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_24 <= _GEN_874;
          end else begin
            reservedRegMap1_24 <= frontEndRegMap_24; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_24 <= _GEN_2040;
        end
      end else begin
        reservedRegMap1_24 <= _GEN_2040;
      end
    end else begin
      reservedRegMap1_24 <= _GEN_2040;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_25 <= _GEN_875;
          end else begin
            reservedRegMap1_25 <= frontEndRegMap_25; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_25 <= _GEN_2041;
        end
      end else begin
        reservedRegMap1_25 <= _GEN_2041;
      end
    end else begin
      reservedRegMap1_25 <= _GEN_2041;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_26 <= _GEN_876;
          end else begin
            reservedRegMap1_26 <= frontEndRegMap_26; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_26 <= _GEN_2042;
        end
      end else begin
        reservedRegMap1_26 <= _GEN_2042;
      end
    end else begin
      reservedRegMap1_26 <= _GEN_2042;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_27 <= _GEN_877;
          end else begin
            reservedRegMap1_27 <= frontEndRegMap_27; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_27 <= _GEN_2043;
        end
      end else begin
        reservedRegMap1_27 <= _GEN_2043;
      end
    end else begin
      reservedRegMap1_27 <= _GEN_2043;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_28 <= _GEN_878;
          end else begin
            reservedRegMap1_28 <= frontEndRegMap_28; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_28 <= _GEN_2044;
        end
      end else begin
        reservedRegMap1_28 <= _GEN_2044;
      end
    end else begin
      reservedRegMap1_28 <= _GEN_2044;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_29 <= _GEN_879;
          end else begin
            reservedRegMap1_29 <= frontEndRegMap_29; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_29 <= _GEN_2045;
        end
      end else begin
        reservedRegMap1_29 <= _GEN_2045;
      end
    end else begin
      reservedRegMap1_29 <= _GEN_2045;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_30 <= _GEN_880;
          end else begin
            reservedRegMap1_30 <= frontEndRegMap_30; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_30 <= _GEN_2046;
        end
      end else begin
        reservedRegMap1_30 <= _GEN_2046;
      end
    end else begin
      reservedRegMap1_30 <= _GEN_2046;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedRegMap1_31 <= _GEN_881;
          end else begin
            reservedRegMap1_31 <= frontEndRegMap_31; // @[decode.scala 402:30]
          end
        end else begin
          reservedRegMap1_31 <= _GEN_2047;
        end
      end else begin
        reservedRegMap1_31 <= _GEN_2047;
      end
    end else begin
      reservedRegMap1_31 <= _GEN_2047;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_0 <= _GEN_2048;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_0 <= _GEN_2664;
        end else begin
          reservedRegMap2_0 <= _GEN_2048;
        end
      end else begin
        reservedRegMap2_0 <= _GEN_2048;
      end
    end else begin
      reservedRegMap2_0 <= _GEN_2048;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_1 <= _GEN_2049;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_1 <= _GEN_2665;
        end else begin
          reservedRegMap2_1 <= _GEN_2049;
        end
      end else begin
        reservedRegMap2_1 <= _GEN_2049;
      end
    end else begin
      reservedRegMap2_1 <= _GEN_2049;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_2 <= _GEN_2050;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_2 <= _GEN_2666;
        end else begin
          reservedRegMap2_2 <= _GEN_2050;
        end
      end else begin
        reservedRegMap2_2 <= _GEN_2050;
      end
    end else begin
      reservedRegMap2_2 <= _GEN_2050;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_3 <= _GEN_2051;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_3 <= _GEN_2667;
        end else begin
          reservedRegMap2_3 <= _GEN_2051;
        end
      end else begin
        reservedRegMap2_3 <= _GEN_2051;
      end
    end else begin
      reservedRegMap2_3 <= _GEN_2051;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_4 <= _GEN_2052;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_4 <= _GEN_2668;
        end else begin
          reservedRegMap2_4 <= _GEN_2052;
        end
      end else begin
        reservedRegMap2_4 <= _GEN_2052;
      end
    end else begin
      reservedRegMap2_4 <= _GEN_2052;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_5 <= _GEN_2053;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_5 <= _GEN_2669;
        end else begin
          reservedRegMap2_5 <= _GEN_2053;
        end
      end else begin
        reservedRegMap2_5 <= _GEN_2053;
      end
    end else begin
      reservedRegMap2_5 <= _GEN_2053;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_6 <= _GEN_2054;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_6 <= _GEN_2670;
        end else begin
          reservedRegMap2_6 <= _GEN_2054;
        end
      end else begin
        reservedRegMap2_6 <= _GEN_2054;
      end
    end else begin
      reservedRegMap2_6 <= _GEN_2054;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_7 <= _GEN_2055;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_7 <= _GEN_2671;
        end else begin
          reservedRegMap2_7 <= _GEN_2055;
        end
      end else begin
        reservedRegMap2_7 <= _GEN_2055;
      end
    end else begin
      reservedRegMap2_7 <= _GEN_2055;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_8 <= _GEN_2056;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_8 <= _GEN_2672;
        end else begin
          reservedRegMap2_8 <= _GEN_2056;
        end
      end else begin
        reservedRegMap2_8 <= _GEN_2056;
      end
    end else begin
      reservedRegMap2_8 <= _GEN_2056;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_9 <= _GEN_2057;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_9 <= _GEN_2673;
        end else begin
          reservedRegMap2_9 <= _GEN_2057;
        end
      end else begin
        reservedRegMap2_9 <= _GEN_2057;
      end
    end else begin
      reservedRegMap2_9 <= _GEN_2057;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_10 <= _GEN_2058;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_10 <= _GEN_2674;
        end else begin
          reservedRegMap2_10 <= _GEN_2058;
        end
      end else begin
        reservedRegMap2_10 <= _GEN_2058;
      end
    end else begin
      reservedRegMap2_10 <= _GEN_2058;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_11 <= _GEN_2059;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_11 <= _GEN_2675;
        end else begin
          reservedRegMap2_11 <= _GEN_2059;
        end
      end else begin
        reservedRegMap2_11 <= _GEN_2059;
      end
    end else begin
      reservedRegMap2_11 <= _GEN_2059;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_12 <= _GEN_2060;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_12 <= _GEN_2676;
        end else begin
          reservedRegMap2_12 <= _GEN_2060;
        end
      end else begin
        reservedRegMap2_12 <= _GEN_2060;
      end
    end else begin
      reservedRegMap2_12 <= _GEN_2060;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_13 <= _GEN_2061;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_13 <= _GEN_2677;
        end else begin
          reservedRegMap2_13 <= _GEN_2061;
        end
      end else begin
        reservedRegMap2_13 <= _GEN_2061;
      end
    end else begin
      reservedRegMap2_13 <= _GEN_2061;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_14 <= _GEN_2062;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_14 <= _GEN_2678;
        end else begin
          reservedRegMap2_14 <= _GEN_2062;
        end
      end else begin
        reservedRegMap2_14 <= _GEN_2062;
      end
    end else begin
      reservedRegMap2_14 <= _GEN_2062;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_15 <= _GEN_2063;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_15 <= _GEN_2679;
        end else begin
          reservedRegMap2_15 <= _GEN_2063;
        end
      end else begin
        reservedRegMap2_15 <= _GEN_2063;
      end
    end else begin
      reservedRegMap2_15 <= _GEN_2063;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_16 <= _GEN_2064;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_16 <= _GEN_2680;
        end else begin
          reservedRegMap2_16 <= _GEN_2064;
        end
      end else begin
        reservedRegMap2_16 <= _GEN_2064;
      end
    end else begin
      reservedRegMap2_16 <= _GEN_2064;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_17 <= _GEN_2065;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_17 <= _GEN_2681;
        end else begin
          reservedRegMap2_17 <= _GEN_2065;
        end
      end else begin
        reservedRegMap2_17 <= _GEN_2065;
      end
    end else begin
      reservedRegMap2_17 <= _GEN_2065;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_18 <= _GEN_2066;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_18 <= _GEN_2682;
        end else begin
          reservedRegMap2_18 <= _GEN_2066;
        end
      end else begin
        reservedRegMap2_18 <= _GEN_2066;
      end
    end else begin
      reservedRegMap2_18 <= _GEN_2066;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_19 <= _GEN_2067;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_19 <= _GEN_2683;
        end else begin
          reservedRegMap2_19 <= _GEN_2067;
        end
      end else begin
        reservedRegMap2_19 <= _GEN_2067;
      end
    end else begin
      reservedRegMap2_19 <= _GEN_2067;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_20 <= _GEN_2068;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_20 <= _GEN_2684;
        end else begin
          reservedRegMap2_20 <= _GEN_2068;
        end
      end else begin
        reservedRegMap2_20 <= _GEN_2068;
      end
    end else begin
      reservedRegMap2_20 <= _GEN_2068;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_21 <= _GEN_2069;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_21 <= _GEN_2685;
        end else begin
          reservedRegMap2_21 <= _GEN_2069;
        end
      end else begin
        reservedRegMap2_21 <= _GEN_2069;
      end
    end else begin
      reservedRegMap2_21 <= _GEN_2069;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_22 <= _GEN_2070;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_22 <= _GEN_2686;
        end else begin
          reservedRegMap2_22 <= _GEN_2070;
        end
      end else begin
        reservedRegMap2_22 <= _GEN_2070;
      end
    end else begin
      reservedRegMap2_22 <= _GEN_2070;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_23 <= _GEN_2071;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_23 <= _GEN_2687;
        end else begin
          reservedRegMap2_23 <= _GEN_2071;
        end
      end else begin
        reservedRegMap2_23 <= _GEN_2071;
      end
    end else begin
      reservedRegMap2_23 <= _GEN_2071;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_24 <= _GEN_2072;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_24 <= _GEN_2688;
        end else begin
          reservedRegMap2_24 <= _GEN_2072;
        end
      end else begin
        reservedRegMap2_24 <= _GEN_2072;
      end
    end else begin
      reservedRegMap2_24 <= _GEN_2072;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_25 <= _GEN_2073;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_25 <= _GEN_2689;
        end else begin
          reservedRegMap2_25 <= _GEN_2073;
        end
      end else begin
        reservedRegMap2_25 <= _GEN_2073;
      end
    end else begin
      reservedRegMap2_25 <= _GEN_2073;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_26 <= _GEN_2074;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_26 <= _GEN_2690;
        end else begin
          reservedRegMap2_26 <= _GEN_2074;
        end
      end else begin
        reservedRegMap2_26 <= _GEN_2074;
      end
    end else begin
      reservedRegMap2_26 <= _GEN_2074;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_27 <= _GEN_2075;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_27 <= _GEN_2691;
        end else begin
          reservedRegMap2_27 <= _GEN_2075;
        end
      end else begin
        reservedRegMap2_27 <= _GEN_2075;
      end
    end else begin
      reservedRegMap2_27 <= _GEN_2075;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_28 <= _GEN_2076;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_28 <= _GEN_2692;
        end else begin
          reservedRegMap2_28 <= _GEN_2076;
        end
      end else begin
        reservedRegMap2_28 <= _GEN_2076;
      end
    end else begin
      reservedRegMap2_28 <= _GEN_2076;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_29 <= _GEN_2077;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_29 <= _GEN_2693;
        end else begin
          reservedRegMap2_29 <= _GEN_2077;
        end
      end else begin
        reservedRegMap2_29 <= _GEN_2077;
      end
    end else begin
      reservedRegMap2_29 <= _GEN_2077;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_30 <= _GEN_2078;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_30 <= _GEN_2694;
        end else begin
          reservedRegMap2_30 <= _GEN_2078;
        end
      end else begin
        reservedRegMap2_30 <= _GEN_2078;
      end
    end else begin
      reservedRegMap2_30 <= _GEN_2078;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_31 <= _GEN_2079;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap2_31 <= _GEN_2695;
        end else begin
          reservedRegMap2_31 <= _GEN_2079;
        end
      end else begin
        reservedRegMap2_31 <= _GEN_2079;
      end
    end else begin
      reservedRegMap2_31 <= _GEN_2079;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_0 <= _GEN_2080;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_0 <= _GEN_2080;
        end else begin
          reservedRegMap3_0 <= _GEN_3944;
        end
      end else begin
        reservedRegMap3_0 <= _GEN_2080;
      end
    end else begin
      reservedRegMap3_0 <= _GEN_2080;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_1 <= _GEN_2081;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_1 <= _GEN_2081;
        end else begin
          reservedRegMap3_1 <= _GEN_3945;
        end
      end else begin
        reservedRegMap3_1 <= _GEN_2081;
      end
    end else begin
      reservedRegMap3_1 <= _GEN_2081;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_2 <= _GEN_2082;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_2 <= _GEN_2082;
        end else begin
          reservedRegMap3_2 <= _GEN_3946;
        end
      end else begin
        reservedRegMap3_2 <= _GEN_2082;
      end
    end else begin
      reservedRegMap3_2 <= _GEN_2082;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_3 <= _GEN_2083;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_3 <= _GEN_2083;
        end else begin
          reservedRegMap3_3 <= _GEN_3947;
        end
      end else begin
        reservedRegMap3_3 <= _GEN_2083;
      end
    end else begin
      reservedRegMap3_3 <= _GEN_2083;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_4 <= _GEN_2084;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_4 <= _GEN_2084;
        end else begin
          reservedRegMap3_4 <= _GEN_3948;
        end
      end else begin
        reservedRegMap3_4 <= _GEN_2084;
      end
    end else begin
      reservedRegMap3_4 <= _GEN_2084;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_5 <= _GEN_2085;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_5 <= _GEN_2085;
        end else begin
          reservedRegMap3_5 <= _GEN_3949;
        end
      end else begin
        reservedRegMap3_5 <= _GEN_2085;
      end
    end else begin
      reservedRegMap3_5 <= _GEN_2085;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_6 <= _GEN_2086;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_6 <= _GEN_2086;
        end else begin
          reservedRegMap3_6 <= _GEN_3950;
        end
      end else begin
        reservedRegMap3_6 <= _GEN_2086;
      end
    end else begin
      reservedRegMap3_6 <= _GEN_2086;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_7 <= _GEN_2087;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_7 <= _GEN_2087;
        end else begin
          reservedRegMap3_7 <= _GEN_3951;
        end
      end else begin
        reservedRegMap3_7 <= _GEN_2087;
      end
    end else begin
      reservedRegMap3_7 <= _GEN_2087;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_8 <= _GEN_2088;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_8 <= _GEN_2088;
        end else begin
          reservedRegMap3_8 <= _GEN_3952;
        end
      end else begin
        reservedRegMap3_8 <= _GEN_2088;
      end
    end else begin
      reservedRegMap3_8 <= _GEN_2088;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_9 <= _GEN_2089;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_9 <= _GEN_2089;
        end else begin
          reservedRegMap3_9 <= _GEN_3953;
        end
      end else begin
        reservedRegMap3_9 <= _GEN_2089;
      end
    end else begin
      reservedRegMap3_9 <= _GEN_2089;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_10 <= _GEN_2090;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_10 <= _GEN_2090;
        end else begin
          reservedRegMap3_10 <= _GEN_3954;
        end
      end else begin
        reservedRegMap3_10 <= _GEN_2090;
      end
    end else begin
      reservedRegMap3_10 <= _GEN_2090;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_11 <= _GEN_2091;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_11 <= _GEN_2091;
        end else begin
          reservedRegMap3_11 <= _GEN_3955;
        end
      end else begin
        reservedRegMap3_11 <= _GEN_2091;
      end
    end else begin
      reservedRegMap3_11 <= _GEN_2091;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_12 <= _GEN_2092;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_12 <= _GEN_2092;
        end else begin
          reservedRegMap3_12 <= _GEN_3956;
        end
      end else begin
        reservedRegMap3_12 <= _GEN_2092;
      end
    end else begin
      reservedRegMap3_12 <= _GEN_2092;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_13 <= _GEN_2093;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_13 <= _GEN_2093;
        end else begin
          reservedRegMap3_13 <= _GEN_3957;
        end
      end else begin
        reservedRegMap3_13 <= _GEN_2093;
      end
    end else begin
      reservedRegMap3_13 <= _GEN_2093;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_14 <= _GEN_2094;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_14 <= _GEN_2094;
        end else begin
          reservedRegMap3_14 <= _GEN_3958;
        end
      end else begin
        reservedRegMap3_14 <= _GEN_2094;
      end
    end else begin
      reservedRegMap3_14 <= _GEN_2094;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_15 <= _GEN_2095;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_15 <= _GEN_2095;
        end else begin
          reservedRegMap3_15 <= _GEN_3959;
        end
      end else begin
        reservedRegMap3_15 <= _GEN_2095;
      end
    end else begin
      reservedRegMap3_15 <= _GEN_2095;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_16 <= _GEN_2096;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_16 <= _GEN_2096;
        end else begin
          reservedRegMap3_16 <= _GEN_3960;
        end
      end else begin
        reservedRegMap3_16 <= _GEN_2096;
      end
    end else begin
      reservedRegMap3_16 <= _GEN_2096;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_17 <= _GEN_2097;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_17 <= _GEN_2097;
        end else begin
          reservedRegMap3_17 <= _GEN_3961;
        end
      end else begin
        reservedRegMap3_17 <= _GEN_2097;
      end
    end else begin
      reservedRegMap3_17 <= _GEN_2097;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_18 <= _GEN_2098;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_18 <= _GEN_2098;
        end else begin
          reservedRegMap3_18 <= _GEN_3962;
        end
      end else begin
        reservedRegMap3_18 <= _GEN_2098;
      end
    end else begin
      reservedRegMap3_18 <= _GEN_2098;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_19 <= _GEN_2099;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_19 <= _GEN_2099;
        end else begin
          reservedRegMap3_19 <= _GEN_3963;
        end
      end else begin
        reservedRegMap3_19 <= _GEN_2099;
      end
    end else begin
      reservedRegMap3_19 <= _GEN_2099;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_20 <= _GEN_2100;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_20 <= _GEN_2100;
        end else begin
          reservedRegMap3_20 <= _GEN_3964;
        end
      end else begin
        reservedRegMap3_20 <= _GEN_2100;
      end
    end else begin
      reservedRegMap3_20 <= _GEN_2100;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_21 <= _GEN_2101;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_21 <= _GEN_2101;
        end else begin
          reservedRegMap3_21 <= _GEN_3965;
        end
      end else begin
        reservedRegMap3_21 <= _GEN_2101;
      end
    end else begin
      reservedRegMap3_21 <= _GEN_2101;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_22 <= _GEN_2102;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_22 <= _GEN_2102;
        end else begin
          reservedRegMap3_22 <= _GEN_3966;
        end
      end else begin
        reservedRegMap3_22 <= _GEN_2102;
      end
    end else begin
      reservedRegMap3_22 <= _GEN_2102;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_23 <= _GEN_2103;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_23 <= _GEN_2103;
        end else begin
          reservedRegMap3_23 <= _GEN_3967;
        end
      end else begin
        reservedRegMap3_23 <= _GEN_2103;
      end
    end else begin
      reservedRegMap3_23 <= _GEN_2103;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_24 <= _GEN_2104;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_24 <= _GEN_2104;
        end else begin
          reservedRegMap3_24 <= _GEN_3968;
        end
      end else begin
        reservedRegMap3_24 <= _GEN_2104;
      end
    end else begin
      reservedRegMap3_24 <= _GEN_2104;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_25 <= _GEN_2105;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_25 <= _GEN_2105;
        end else begin
          reservedRegMap3_25 <= _GEN_3969;
        end
      end else begin
        reservedRegMap3_25 <= _GEN_2105;
      end
    end else begin
      reservedRegMap3_25 <= _GEN_2105;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_26 <= _GEN_2106;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_26 <= _GEN_2106;
        end else begin
          reservedRegMap3_26 <= _GEN_3970;
        end
      end else begin
        reservedRegMap3_26 <= _GEN_2106;
      end
    end else begin
      reservedRegMap3_26 <= _GEN_2106;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_27 <= _GEN_2107;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_27 <= _GEN_2107;
        end else begin
          reservedRegMap3_27 <= _GEN_3971;
        end
      end else begin
        reservedRegMap3_27 <= _GEN_2107;
      end
    end else begin
      reservedRegMap3_27 <= _GEN_2107;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_28 <= _GEN_2108;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_28 <= _GEN_2108;
        end else begin
          reservedRegMap3_28 <= _GEN_3972;
        end
      end else begin
        reservedRegMap3_28 <= _GEN_2108;
      end
    end else begin
      reservedRegMap3_28 <= _GEN_2108;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_29 <= _GEN_2109;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_29 <= _GEN_2109;
        end else begin
          reservedRegMap3_29 <= _GEN_3973;
        end
      end else begin
        reservedRegMap3_29 <= _GEN_2109;
      end
    end else begin
      reservedRegMap3_29 <= _GEN_2109;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_30 <= _GEN_2110;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_30 <= _GEN_2110;
        end else begin
          reservedRegMap3_30 <= _GEN_3974;
        end
      end else begin
        reservedRegMap3_30 <= _GEN_2110;
      end
    end else begin
      reservedRegMap3_30 <= _GEN_2110;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_31 <= _GEN_2111;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedRegMap3_31 <= _GEN_2111;
        end else begin
          reservedRegMap3_31 <= _GEN_3975;
        end
      end else begin
        reservedRegMap3_31 <= _GEN_2111;
      end
    end else begin
      reservedRegMap3_31 <= _GEN_2111;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_0 <= _GEN_4104;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_1 <= _GEN_4105;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_2 <= _GEN_4106;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_3 <= _GEN_4107;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_4 <= _GEN_4108;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_5 <= _GEN_4109;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_6 <= _GEN_4110;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_7 <= _GEN_4111;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_8 <= _GEN_4112;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_9 <= _GEN_4113;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_10 <= _GEN_4114;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_11 <= _GEN_4115;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_12 <= _GEN_4116;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_13 <= _GEN_4117;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_14 <= _GEN_4118;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_15 <= _GEN_4119;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_16 <= _GEN_4120;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_17 <= _GEN_4121;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_18 <= _GEN_4122;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_19 <= _GEN_4123;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_20 <= _GEN_4124;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_21 <= _GEN_4125;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_22 <= _GEN_4126;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_23 <= _GEN_4127;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_24 <= _GEN_4128;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_25 <= _GEN_4129;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_26 <= _GEN_4130;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_27 <= _GEN_4131;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_28 <= _GEN_4132;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_29 <= _GEN_4133;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_30 <= _GEN_4134;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedRegMap4_31 <= _GEN_4135;
          end
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_0 <= _GEN_9262;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_0 <= _GEN_2696;
        end else begin
          reservedFreeList1_0 <= _GEN_2112;
        end
      end else begin
        reservedFreeList1_0 <= _GEN_2112;
      end
    end else begin
      reservedFreeList1_0 <= _GEN_2112;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_1 <= _GEN_9263;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_1 <= _GEN_2697;
        end else begin
          reservedFreeList1_1 <= _GEN_2113;
        end
      end else begin
        reservedFreeList1_1 <= _GEN_2113;
      end
    end else begin
      reservedFreeList1_1 <= _GEN_2113;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_2 <= _GEN_9264;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_2 <= _GEN_2698;
        end else begin
          reservedFreeList1_2 <= _GEN_2114;
        end
      end else begin
        reservedFreeList1_2 <= _GEN_2114;
      end
    end else begin
      reservedFreeList1_2 <= _GEN_2114;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_3 <= _GEN_9265;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_3 <= _GEN_2699;
        end else begin
          reservedFreeList1_3 <= _GEN_2115;
        end
      end else begin
        reservedFreeList1_3 <= _GEN_2115;
      end
    end else begin
      reservedFreeList1_3 <= _GEN_2115;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_4 <= _GEN_9266;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_4 <= _GEN_2700;
        end else begin
          reservedFreeList1_4 <= _GEN_2116;
        end
      end else begin
        reservedFreeList1_4 <= _GEN_2116;
      end
    end else begin
      reservedFreeList1_4 <= _GEN_2116;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_5 <= _GEN_9267;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_5 <= _GEN_2701;
        end else begin
          reservedFreeList1_5 <= _GEN_2117;
        end
      end else begin
        reservedFreeList1_5 <= _GEN_2117;
      end
    end else begin
      reservedFreeList1_5 <= _GEN_2117;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_6 <= _GEN_9268;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_6 <= _GEN_2702;
        end else begin
          reservedFreeList1_6 <= _GEN_2118;
        end
      end else begin
        reservedFreeList1_6 <= _GEN_2118;
      end
    end else begin
      reservedFreeList1_6 <= _GEN_2118;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_7 <= _GEN_9269;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_7 <= _GEN_2703;
        end else begin
          reservedFreeList1_7 <= _GEN_2119;
        end
      end else begin
        reservedFreeList1_7 <= _GEN_2119;
      end
    end else begin
      reservedFreeList1_7 <= _GEN_2119;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_8 <= _GEN_9270;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_8 <= _GEN_2704;
        end else begin
          reservedFreeList1_8 <= _GEN_2120;
        end
      end else begin
        reservedFreeList1_8 <= _GEN_2120;
      end
    end else begin
      reservedFreeList1_8 <= _GEN_2120;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_9 <= _GEN_9271;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_9 <= _GEN_2705;
        end else begin
          reservedFreeList1_9 <= _GEN_2121;
        end
      end else begin
        reservedFreeList1_9 <= _GEN_2121;
      end
    end else begin
      reservedFreeList1_9 <= _GEN_2121;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_10 <= _GEN_9272;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_10 <= _GEN_2706;
        end else begin
          reservedFreeList1_10 <= _GEN_2122;
        end
      end else begin
        reservedFreeList1_10 <= _GEN_2122;
      end
    end else begin
      reservedFreeList1_10 <= _GEN_2122;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_11 <= _GEN_9273;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_11 <= _GEN_2707;
        end else begin
          reservedFreeList1_11 <= _GEN_2123;
        end
      end else begin
        reservedFreeList1_11 <= _GEN_2123;
      end
    end else begin
      reservedFreeList1_11 <= _GEN_2123;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_12 <= _GEN_9274;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_12 <= _GEN_2708;
        end else begin
          reservedFreeList1_12 <= _GEN_2124;
        end
      end else begin
        reservedFreeList1_12 <= _GEN_2124;
      end
    end else begin
      reservedFreeList1_12 <= _GEN_2124;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_13 <= _GEN_9275;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_13 <= _GEN_2709;
        end else begin
          reservedFreeList1_13 <= _GEN_2125;
        end
      end else begin
        reservedFreeList1_13 <= _GEN_2125;
      end
    end else begin
      reservedFreeList1_13 <= _GEN_2125;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_14 <= _GEN_9276;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_14 <= _GEN_2710;
        end else begin
          reservedFreeList1_14 <= _GEN_2126;
        end
      end else begin
        reservedFreeList1_14 <= _GEN_2126;
      end
    end else begin
      reservedFreeList1_14 <= _GEN_2126;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_15 <= _GEN_9277;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_15 <= _GEN_2711;
        end else begin
          reservedFreeList1_15 <= _GEN_2127;
        end
      end else begin
        reservedFreeList1_15 <= _GEN_2127;
      end
    end else begin
      reservedFreeList1_15 <= _GEN_2127;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_16 <= _GEN_9278;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_16 <= _GEN_2712;
        end else begin
          reservedFreeList1_16 <= _GEN_2128;
        end
      end else begin
        reservedFreeList1_16 <= _GEN_2128;
      end
    end else begin
      reservedFreeList1_16 <= _GEN_2128;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_17 <= _GEN_9279;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_17 <= _GEN_2713;
        end else begin
          reservedFreeList1_17 <= _GEN_2129;
        end
      end else begin
        reservedFreeList1_17 <= _GEN_2129;
      end
    end else begin
      reservedFreeList1_17 <= _GEN_2129;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_18 <= _GEN_9280;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_18 <= _GEN_2714;
        end else begin
          reservedFreeList1_18 <= _GEN_2130;
        end
      end else begin
        reservedFreeList1_18 <= _GEN_2130;
      end
    end else begin
      reservedFreeList1_18 <= _GEN_2130;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_19 <= _GEN_9281;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_19 <= _GEN_2715;
        end else begin
          reservedFreeList1_19 <= _GEN_2131;
        end
      end else begin
        reservedFreeList1_19 <= _GEN_2131;
      end
    end else begin
      reservedFreeList1_19 <= _GEN_2131;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_20 <= _GEN_9282;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_20 <= _GEN_2716;
        end else begin
          reservedFreeList1_20 <= _GEN_2132;
        end
      end else begin
        reservedFreeList1_20 <= _GEN_2132;
      end
    end else begin
      reservedFreeList1_20 <= _GEN_2132;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_21 <= _GEN_9283;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_21 <= _GEN_2717;
        end else begin
          reservedFreeList1_21 <= _GEN_2133;
        end
      end else begin
        reservedFreeList1_21 <= _GEN_2133;
      end
    end else begin
      reservedFreeList1_21 <= _GEN_2133;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_22 <= _GEN_9284;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_22 <= _GEN_2718;
        end else begin
          reservedFreeList1_22 <= _GEN_2134;
        end
      end else begin
        reservedFreeList1_22 <= _GEN_2134;
      end
    end else begin
      reservedFreeList1_22 <= _GEN_2134;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_23 <= _GEN_9285;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_23 <= _GEN_2719;
        end else begin
          reservedFreeList1_23 <= _GEN_2135;
        end
      end else begin
        reservedFreeList1_23 <= _GEN_2135;
      end
    end else begin
      reservedFreeList1_23 <= _GEN_2135;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_24 <= _GEN_9286;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_24 <= _GEN_2720;
        end else begin
          reservedFreeList1_24 <= _GEN_2136;
        end
      end else begin
        reservedFreeList1_24 <= _GEN_2136;
      end
    end else begin
      reservedFreeList1_24 <= _GEN_2136;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_25 <= _GEN_9287;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_25 <= _GEN_2721;
        end else begin
          reservedFreeList1_25 <= _GEN_2137;
        end
      end else begin
        reservedFreeList1_25 <= _GEN_2137;
      end
    end else begin
      reservedFreeList1_25 <= _GEN_2137;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_26 <= _GEN_9288;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_26 <= _GEN_2722;
        end else begin
          reservedFreeList1_26 <= _GEN_2138;
        end
      end else begin
        reservedFreeList1_26 <= _GEN_2138;
      end
    end else begin
      reservedFreeList1_26 <= _GEN_2138;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_27 <= _GEN_9289;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_27 <= _GEN_2723;
        end else begin
          reservedFreeList1_27 <= _GEN_2139;
        end
      end else begin
        reservedFreeList1_27 <= _GEN_2139;
      end
    end else begin
      reservedFreeList1_27 <= _GEN_2139;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_28 <= _GEN_9290;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_28 <= _GEN_2724;
        end else begin
          reservedFreeList1_28 <= _GEN_2140;
        end
      end else begin
        reservedFreeList1_28 <= _GEN_2140;
      end
    end else begin
      reservedFreeList1_28 <= _GEN_2140;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_29 <= _GEN_9291;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_29 <= _GEN_2725;
        end else begin
          reservedFreeList1_29 <= _GEN_2141;
        end
      end else begin
        reservedFreeList1_29 <= _GEN_2141;
      end
    end else begin
      reservedFreeList1_29 <= _GEN_2141;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_30 <= _GEN_9292;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_30 <= _GEN_2726;
        end else begin
          reservedFreeList1_30 <= _GEN_2142;
        end
      end else begin
        reservedFreeList1_30 <= _GEN_2142;
      end
    end else begin
      reservedFreeList1_30 <= _GEN_2142;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_31 <= _GEN_9293;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_31 <= _GEN_2727;
        end else begin
          reservedFreeList1_31 <= _GEN_2143;
        end
      end else begin
        reservedFreeList1_31 <= _GEN_2143;
      end
    end else begin
      reservedFreeList1_31 <= _GEN_2143;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_32 <= _GEN_9294;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_32 <= _GEN_2728;
        end else begin
          reservedFreeList1_32 <= _GEN_2144;
        end
      end else begin
        reservedFreeList1_32 <= _GEN_2144;
      end
    end else begin
      reservedFreeList1_32 <= _GEN_2144;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_33 <= _GEN_9295;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_33 <= _GEN_2729;
        end else begin
          reservedFreeList1_33 <= _GEN_2145;
        end
      end else begin
        reservedFreeList1_33 <= _GEN_2145;
      end
    end else begin
      reservedFreeList1_33 <= _GEN_2145;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_34 <= _GEN_9296;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_34 <= _GEN_2730;
        end else begin
          reservedFreeList1_34 <= _GEN_2146;
        end
      end else begin
        reservedFreeList1_34 <= _GEN_2146;
      end
    end else begin
      reservedFreeList1_34 <= _GEN_2146;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_35 <= _GEN_9297;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_35 <= _GEN_2731;
        end else begin
          reservedFreeList1_35 <= _GEN_2147;
        end
      end else begin
        reservedFreeList1_35 <= _GEN_2147;
      end
    end else begin
      reservedFreeList1_35 <= _GEN_2147;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_36 <= _GEN_9298;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_36 <= _GEN_2732;
        end else begin
          reservedFreeList1_36 <= _GEN_2148;
        end
      end else begin
        reservedFreeList1_36 <= _GEN_2148;
      end
    end else begin
      reservedFreeList1_36 <= _GEN_2148;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_37 <= _GEN_9299;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_37 <= _GEN_2733;
        end else begin
          reservedFreeList1_37 <= _GEN_2149;
        end
      end else begin
        reservedFreeList1_37 <= _GEN_2149;
      end
    end else begin
      reservedFreeList1_37 <= _GEN_2149;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_38 <= _GEN_9300;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_38 <= _GEN_2734;
        end else begin
          reservedFreeList1_38 <= _GEN_2150;
        end
      end else begin
        reservedFreeList1_38 <= _GEN_2150;
      end
    end else begin
      reservedFreeList1_38 <= _GEN_2150;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_39 <= _GEN_9301;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_39 <= _GEN_2735;
        end else begin
          reservedFreeList1_39 <= _GEN_2151;
        end
      end else begin
        reservedFreeList1_39 <= _GEN_2151;
      end
    end else begin
      reservedFreeList1_39 <= _GEN_2151;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_40 <= _GEN_9302;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_40 <= _GEN_2736;
        end else begin
          reservedFreeList1_40 <= _GEN_2152;
        end
      end else begin
        reservedFreeList1_40 <= _GEN_2152;
      end
    end else begin
      reservedFreeList1_40 <= _GEN_2152;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_41 <= _GEN_9303;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_41 <= _GEN_2737;
        end else begin
          reservedFreeList1_41 <= _GEN_2153;
        end
      end else begin
        reservedFreeList1_41 <= _GEN_2153;
      end
    end else begin
      reservedFreeList1_41 <= _GEN_2153;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_42 <= _GEN_9304;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_42 <= _GEN_2738;
        end else begin
          reservedFreeList1_42 <= _GEN_2154;
        end
      end else begin
        reservedFreeList1_42 <= _GEN_2154;
      end
    end else begin
      reservedFreeList1_42 <= _GEN_2154;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_43 <= _GEN_9305;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_43 <= _GEN_2739;
        end else begin
          reservedFreeList1_43 <= _GEN_2155;
        end
      end else begin
        reservedFreeList1_43 <= _GEN_2155;
      end
    end else begin
      reservedFreeList1_43 <= _GEN_2155;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_44 <= _GEN_9306;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_44 <= _GEN_2740;
        end else begin
          reservedFreeList1_44 <= _GEN_2156;
        end
      end else begin
        reservedFreeList1_44 <= _GEN_2156;
      end
    end else begin
      reservedFreeList1_44 <= _GEN_2156;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_45 <= _GEN_9307;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_45 <= _GEN_2741;
        end else begin
          reservedFreeList1_45 <= _GEN_2157;
        end
      end else begin
        reservedFreeList1_45 <= _GEN_2157;
      end
    end else begin
      reservedFreeList1_45 <= _GEN_2157;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_46 <= _GEN_9308;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_46 <= _GEN_2742;
        end else begin
          reservedFreeList1_46 <= _GEN_2158;
        end
      end else begin
        reservedFreeList1_46 <= _GEN_2158;
      end
    end else begin
      reservedFreeList1_46 <= _GEN_2158;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_47 <= _GEN_9309;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_47 <= _GEN_2743;
        end else begin
          reservedFreeList1_47 <= _GEN_2159;
        end
      end else begin
        reservedFreeList1_47 <= _GEN_2159;
      end
    end else begin
      reservedFreeList1_47 <= _GEN_2159;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_48 <= _GEN_9310;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_48 <= _GEN_2744;
        end else begin
          reservedFreeList1_48 <= _GEN_2160;
        end
      end else begin
        reservedFreeList1_48 <= _GEN_2160;
      end
    end else begin
      reservedFreeList1_48 <= _GEN_2160;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_49 <= _GEN_9311;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_49 <= _GEN_2745;
        end else begin
          reservedFreeList1_49 <= _GEN_2161;
        end
      end else begin
        reservedFreeList1_49 <= _GEN_2161;
      end
    end else begin
      reservedFreeList1_49 <= _GEN_2161;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_50 <= _GEN_9312;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_50 <= _GEN_2746;
        end else begin
          reservedFreeList1_50 <= _GEN_2162;
        end
      end else begin
        reservedFreeList1_50 <= _GEN_2162;
      end
    end else begin
      reservedFreeList1_50 <= _GEN_2162;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_51 <= _GEN_9313;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_51 <= _GEN_2747;
        end else begin
          reservedFreeList1_51 <= _GEN_2163;
        end
      end else begin
        reservedFreeList1_51 <= _GEN_2163;
      end
    end else begin
      reservedFreeList1_51 <= _GEN_2163;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_52 <= _GEN_9314;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_52 <= _GEN_2748;
        end else begin
          reservedFreeList1_52 <= _GEN_2164;
        end
      end else begin
        reservedFreeList1_52 <= _GEN_2164;
      end
    end else begin
      reservedFreeList1_52 <= _GEN_2164;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_53 <= _GEN_9315;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_53 <= _GEN_2749;
        end else begin
          reservedFreeList1_53 <= _GEN_2165;
        end
      end else begin
        reservedFreeList1_53 <= _GEN_2165;
      end
    end else begin
      reservedFreeList1_53 <= _GEN_2165;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_54 <= _GEN_9316;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_54 <= _GEN_2750;
        end else begin
          reservedFreeList1_54 <= _GEN_2166;
        end
      end else begin
        reservedFreeList1_54 <= _GEN_2166;
      end
    end else begin
      reservedFreeList1_54 <= _GEN_2166;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_55 <= _GEN_9317;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_55 <= _GEN_2751;
        end else begin
          reservedFreeList1_55 <= _GEN_2167;
        end
      end else begin
        reservedFreeList1_55 <= _GEN_2167;
      end
    end else begin
      reservedFreeList1_55 <= _GEN_2167;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_56 <= _GEN_9318;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_56 <= _GEN_2752;
        end else begin
          reservedFreeList1_56 <= _GEN_2168;
        end
      end else begin
        reservedFreeList1_56 <= _GEN_2168;
      end
    end else begin
      reservedFreeList1_56 <= _GEN_2168;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_57 <= _GEN_9319;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_57 <= _GEN_2753;
        end else begin
          reservedFreeList1_57 <= _GEN_2169;
        end
      end else begin
        reservedFreeList1_57 <= _GEN_2169;
      end
    end else begin
      reservedFreeList1_57 <= _GEN_2169;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_58 <= _GEN_9320;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_58 <= _GEN_2754;
        end else begin
          reservedFreeList1_58 <= _GEN_2170;
        end
      end else begin
        reservedFreeList1_58 <= _GEN_2170;
      end
    end else begin
      reservedFreeList1_58 <= _GEN_2170;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_59 <= _GEN_9321;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_59 <= _GEN_2755;
        end else begin
          reservedFreeList1_59 <= _GEN_2171;
        end
      end else begin
        reservedFreeList1_59 <= _GEN_2171;
      end
    end else begin
      reservedFreeList1_59 <= _GEN_2171;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_60 <= _GEN_9322;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_60 <= _GEN_2756;
        end else begin
          reservedFreeList1_60 <= _GEN_2172;
        end
      end else begin
        reservedFreeList1_60 <= _GEN_2172;
      end
    end else begin
      reservedFreeList1_60 <= _GEN_2172;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_61 <= _GEN_9323;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_61 <= _GEN_2757;
        end else begin
          reservedFreeList1_61 <= _GEN_2173;
        end
      end else begin
        reservedFreeList1_61 <= _GEN_2173;
      end
    end else begin
      reservedFreeList1_61 <= _GEN_2173;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList1_62 <= _GEN_9324;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList1_62 <= _GEN_2758;
        end else begin
          reservedFreeList1_62 <= _GEN_2174;
        end
      end else begin
        reservedFreeList1_62 <= _GEN_2174;
      end
    end else begin
      reservedFreeList1_62 <= _GEN_2174;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_0 <= _GEN_9326;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_0 <= _GEN_2176;
        end else begin
          reservedFreeList2_0 <= _GEN_4296;
        end
      end else begin
        reservedFreeList2_0 <= _GEN_2176;
      end
    end else begin
      reservedFreeList2_0 <= _GEN_2176;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_1 <= _GEN_9327;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_1 <= _GEN_2177;
        end else begin
          reservedFreeList2_1 <= _GEN_4297;
        end
      end else begin
        reservedFreeList2_1 <= _GEN_2177;
      end
    end else begin
      reservedFreeList2_1 <= _GEN_2177;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_2 <= _GEN_9328;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_2 <= _GEN_2178;
        end else begin
          reservedFreeList2_2 <= _GEN_4298;
        end
      end else begin
        reservedFreeList2_2 <= _GEN_2178;
      end
    end else begin
      reservedFreeList2_2 <= _GEN_2178;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_3 <= _GEN_9329;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_3 <= _GEN_2179;
        end else begin
          reservedFreeList2_3 <= _GEN_4299;
        end
      end else begin
        reservedFreeList2_3 <= _GEN_2179;
      end
    end else begin
      reservedFreeList2_3 <= _GEN_2179;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_4 <= _GEN_9330;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_4 <= _GEN_2180;
        end else begin
          reservedFreeList2_4 <= _GEN_4300;
        end
      end else begin
        reservedFreeList2_4 <= _GEN_2180;
      end
    end else begin
      reservedFreeList2_4 <= _GEN_2180;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_5 <= _GEN_9331;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_5 <= _GEN_2181;
        end else begin
          reservedFreeList2_5 <= _GEN_4301;
        end
      end else begin
        reservedFreeList2_5 <= _GEN_2181;
      end
    end else begin
      reservedFreeList2_5 <= _GEN_2181;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_6 <= _GEN_9332;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_6 <= _GEN_2182;
        end else begin
          reservedFreeList2_6 <= _GEN_4302;
        end
      end else begin
        reservedFreeList2_6 <= _GEN_2182;
      end
    end else begin
      reservedFreeList2_6 <= _GEN_2182;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_7 <= _GEN_9333;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_7 <= _GEN_2183;
        end else begin
          reservedFreeList2_7 <= _GEN_4303;
        end
      end else begin
        reservedFreeList2_7 <= _GEN_2183;
      end
    end else begin
      reservedFreeList2_7 <= _GEN_2183;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_8 <= _GEN_9334;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_8 <= _GEN_2184;
        end else begin
          reservedFreeList2_8 <= _GEN_4304;
        end
      end else begin
        reservedFreeList2_8 <= _GEN_2184;
      end
    end else begin
      reservedFreeList2_8 <= _GEN_2184;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_9 <= _GEN_9335;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_9 <= _GEN_2185;
        end else begin
          reservedFreeList2_9 <= _GEN_4305;
        end
      end else begin
        reservedFreeList2_9 <= _GEN_2185;
      end
    end else begin
      reservedFreeList2_9 <= _GEN_2185;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_10 <= _GEN_9336;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_10 <= _GEN_2186;
        end else begin
          reservedFreeList2_10 <= _GEN_4306;
        end
      end else begin
        reservedFreeList2_10 <= _GEN_2186;
      end
    end else begin
      reservedFreeList2_10 <= _GEN_2186;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_11 <= _GEN_9337;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_11 <= _GEN_2187;
        end else begin
          reservedFreeList2_11 <= _GEN_4307;
        end
      end else begin
        reservedFreeList2_11 <= _GEN_2187;
      end
    end else begin
      reservedFreeList2_11 <= _GEN_2187;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_12 <= _GEN_9338;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_12 <= _GEN_2188;
        end else begin
          reservedFreeList2_12 <= _GEN_4308;
        end
      end else begin
        reservedFreeList2_12 <= _GEN_2188;
      end
    end else begin
      reservedFreeList2_12 <= _GEN_2188;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_13 <= _GEN_9339;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_13 <= _GEN_2189;
        end else begin
          reservedFreeList2_13 <= _GEN_4309;
        end
      end else begin
        reservedFreeList2_13 <= _GEN_2189;
      end
    end else begin
      reservedFreeList2_13 <= _GEN_2189;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_14 <= _GEN_9340;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_14 <= _GEN_2190;
        end else begin
          reservedFreeList2_14 <= _GEN_4310;
        end
      end else begin
        reservedFreeList2_14 <= _GEN_2190;
      end
    end else begin
      reservedFreeList2_14 <= _GEN_2190;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_15 <= _GEN_9341;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_15 <= _GEN_2191;
        end else begin
          reservedFreeList2_15 <= _GEN_4311;
        end
      end else begin
        reservedFreeList2_15 <= _GEN_2191;
      end
    end else begin
      reservedFreeList2_15 <= _GEN_2191;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_16 <= _GEN_9342;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_16 <= _GEN_2192;
        end else begin
          reservedFreeList2_16 <= _GEN_4312;
        end
      end else begin
        reservedFreeList2_16 <= _GEN_2192;
      end
    end else begin
      reservedFreeList2_16 <= _GEN_2192;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_17 <= _GEN_9343;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_17 <= _GEN_2193;
        end else begin
          reservedFreeList2_17 <= _GEN_4313;
        end
      end else begin
        reservedFreeList2_17 <= _GEN_2193;
      end
    end else begin
      reservedFreeList2_17 <= _GEN_2193;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_18 <= _GEN_9344;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_18 <= _GEN_2194;
        end else begin
          reservedFreeList2_18 <= _GEN_4314;
        end
      end else begin
        reservedFreeList2_18 <= _GEN_2194;
      end
    end else begin
      reservedFreeList2_18 <= _GEN_2194;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_19 <= _GEN_9345;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_19 <= _GEN_2195;
        end else begin
          reservedFreeList2_19 <= _GEN_4315;
        end
      end else begin
        reservedFreeList2_19 <= _GEN_2195;
      end
    end else begin
      reservedFreeList2_19 <= _GEN_2195;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_20 <= _GEN_9346;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_20 <= _GEN_2196;
        end else begin
          reservedFreeList2_20 <= _GEN_4316;
        end
      end else begin
        reservedFreeList2_20 <= _GEN_2196;
      end
    end else begin
      reservedFreeList2_20 <= _GEN_2196;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_21 <= _GEN_9347;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_21 <= _GEN_2197;
        end else begin
          reservedFreeList2_21 <= _GEN_4317;
        end
      end else begin
        reservedFreeList2_21 <= _GEN_2197;
      end
    end else begin
      reservedFreeList2_21 <= _GEN_2197;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_22 <= _GEN_9348;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_22 <= _GEN_2198;
        end else begin
          reservedFreeList2_22 <= _GEN_4318;
        end
      end else begin
        reservedFreeList2_22 <= _GEN_2198;
      end
    end else begin
      reservedFreeList2_22 <= _GEN_2198;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_23 <= _GEN_9349;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_23 <= _GEN_2199;
        end else begin
          reservedFreeList2_23 <= _GEN_4319;
        end
      end else begin
        reservedFreeList2_23 <= _GEN_2199;
      end
    end else begin
      reservedFreeList2_23 <= _GEN_2199;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_24 <= _GEN_9350;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_24 <= _GEN_2200;
        end else begin
          reservedFreeList2_24 <= _GEN_4320;
        end
      end else begin
        reservedFreeList2_24 <= _GEN_2200;
      end
    end else begin
      reservedFreeList2_24 <= _GEN_2200;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_25 <= _GEN_9351;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_25 <= _GEN_2201;
        end else begin
          reservedFreeList2_25 <= _GEN_4321;
        end
      end else begin
        reservedFreeList2_25 <= _GEN_2201;
      end
    end else begin
      reservedFreeList2_25 <= _GEN_2201;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_26 <= _GEN_9352;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_26 <= _GEN_2202;
        end else begin
          reservedFreeList2_26 <= _GEN_4322;
        end
      end else begin
        reservedFreeList2_26 <= _GEN_2202;
      end
    end else begin
      reservedFreeList2_26 <= _GEN_2202;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_27 <= _GEN_9353;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_27 <= _GEN_2203;
        end else begin
          reservedFreeList2_27 <= _GEN_4323;
        end
      end else begin
        reservedFreeList2_27 <= _GEN_2203;
      end
    end else begin
      reservedFreeList2_27 <= _GEN_2203;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_28 <= _GEN_9354;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_28 <= _GEN_2204;
        end else begin
          reservedFreeList2_28 <= _GEN_4324;
        end
      end else begin
        reservedFreeList2_28 <= _GEN_2204;
      end
    end else begin
      reservedFreeList2_28 <= _GEN_2204;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_29 <= _GEN_9355;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_29 <= _GEN_2205;
        end else begin
          reservedFreeList2_29 <= _GEN_4325;
        end
      end else begin
        reservedFreeList2_29 <= _GEN_2205;
      end
    end else begin
      reservedFreeList2_29 <= _GEN_2205;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_30 <= _GEN_9356;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_30 <= _GEN_2206;
        end else begin
          reservedFreeList2_30 <= _GEN_4326;
        end
      end else begin
        reservedFreeList2_30 <= _GEN_2206;
      end
    end else begin
      reservedFreeList2_30 <= _GEN_2206;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_31 <= _GEN_9357;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_31 <= _GEN_2207;
        end else begin
          reservedFreeList2_31 <= _GEN_4327;
        end
      end else begin
        reservedFreeList2_31 <= _GEN_2207;
      end
    end else begin
      reservedFreeList2_31 <= _GEN_2207;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_32 <= _GEN_9358;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_32 <= _GEN_2208;
        end else begin
          reservedFreeList2_32 <= _GEN_4328;
        end
      end else begin
        reservedFreeList2_32 <= _GEN_2208;
      end
    end else begin
      reservedFreeList2_32 <= _GEN_2208;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_33 <= _GEN_9359;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_33 <= _GEN_2209;
        end else begin
          reservedFreeList2_33 <= _GEN_4329;
        end
      end else begin
        reservedFreeList2_33 <= _GEN_2209;
      end
    end else begin
      reservedFreeList2_33 <= _GEN_2209;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_34 <= _GEN_9360;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_34 <= _GEN_2210;
        end else begin
          reservedFreeList2_34 <= _GEN_4330;
        end
      end else begin
        reservedFreeList2_34 <= _GEN_2210;
      end
    end else begin
      reservedFreeList2_34 <= _GEN_2210;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_35 <= _GEN_9361;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_35 <= _GEN_2211;
        end else begin
          reservedFreeList2_35 <= _GEN_4331;
        end
      end else begin
        reservedFreeList2_35 <= _GEN_2211;
      end
    end else begin
      reservedFreeList2_35 <= _GEN_2211;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_36 <= _GEN_9362;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_36 <= _GEN_2212;
        end else begin
          reservedFreeList2_36 <= _GEN_4332;
        end
      end else begin
        reservedFreeList2_36 <= _GEN_2212;
      end
    end else begin
      reservedFreeList2_36 <= _GEN_2212;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_37 <= _GEN_9363;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_37 <= _GEN_2213;
        end else begin
          reservedFreeList2_37 <= _GEN_4333;
        end
      end else begin
        reservedFreeList2_37 <= _GEN_2213;
      end
    end else begin
      reservedFreeList2_37 <= _GEN_2213;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_38 <= _GEN_9364;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_38 <= _GEN_2214;
        end else begin
          reservedFreeList2_38 <= _GEN_4334;
        end
      end else begin
        reservedFreeList2_38 <= _GEN_2214;
      end
    end else begin
      reservedFreeList2_38 <= _GEN_2214;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_39 <= _GEN_9365;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_39 <= _GEN_2215;
        end else begin
          reservedFreeList2_39 <= _GEN_4335;
        end
      end else begin
        reservedFreeList2_39 <= _GEN_2215;
      end
    end else begin
      reservedFreeList2_39 <= _GEN_2215;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_40 <= _GEN_9366;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_40 <= _GEN_2216;
        end else begin
          reservedFreeList2_40 <= _GEN_4336;
        end
      end else begin
        reservedFreeList2_40 <= _GEN_2216;
      end
    end else begin
      reservedFreeList2_40 <= _GEN_2216;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_41 <= _GEN_9367;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_41 <= _GEN_2217;
        end else begin
          reservedFreeList2_41 <= _GEN_4337;
        end
      end else begin
        reservedFreeList2_41 <= _GEN_2217;
      end
    end else begin
      reservedFreeList2_41 <= _GEN_2217;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_42 <= _GEN_9368;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_42 <= _GEN_2218;
        end else begin
          reservedFreeList2_42 <= _GEN_4338;
        end
      end else begin
        reservedFreeList2_42 <= _GEN_2218;
      end
    end else begin
      reservedFreeList2_42 <= _GEN_2218;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_43 <= _GEN_9369;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_43 <= _GEN_2219;
        end else begin
          reservedFreeList2_43 <= _GEN_4339;
        end
      end else begin
        reservedFreeList2_43 <= _GEN_2219;
      end
    end else begin
      reservedFreeList2_43 <= _GEN_2219;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_44 <= _GEN_9370;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_44 <= _GEN_2220;
        end else begin
          reservedFreeList2_44 <= _GEN_4340;
        end
      end else begin
        reservedFreeList2_44 <= _GEN_2220;
      end
    end else begin
      reservedFreeList2_44 <= _GEN_2220;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_45 <= _GEN_9371;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_45 <= _GEN_2221;
        end else begin
          reservedFreeList2_45 <= _GEN_4341;
        end
      end else begin
        reservedFreeList2_45 <= _GEN_2221;
      end
    end else begin
      reservedFreeList2_45 <= _GEN_2221;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_46 <= _GEN_9372;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_46 <= _GEN_2222;
        end else begin
          reservedFreeList2_46 <= _GEN_4342;
        end
      end else begin
        reservedFreeList2_46 <= _GEN_2222;
      end
    end else begin
      reservedFreeList2_46 <= _GEN_2222;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_47 <= _GEN_9373;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_47 <= _GEN_2223;
        end else begin
          reservedFreeList2_47 <= _GEN_4343;
        end
      end else begin
        reservedFreeList2_47 <= _GEN_2223;
      end
    end else begin
      reservedFreeList2_47 <= _GEN_2223;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_48 <= _GEN_9374;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_48 <= _GEN_2224;
        end else begin
          reservedFreeList2_48 <= _GEN_4344;
        end
      end else begin
        reservedFreeList2_48 <= _GEN_2224;
      end
    end else begin
      reservedFreeList2_48 <= _GEN_2224;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_49 <= _GEN_9375;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_49 <= _GEN_2225;
        end else begin
          reservedFreeList2_49 <= _GEN_4345;
        end
      end else begin
        reservedFreeList2_49 <= _GEN_2225;
      end
    end else begin
      reservedFreeList2_49 <= _GEN_2225;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_50 <= _GEN_9376;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_50 <= _GEN_2226;
        end else begin
          reservedFreeList2_50 <= _GEN_4346;
        end
      end else begin
        reservedFreeList2_50 <= _GEN_2226;
      end
    end else begin
      reservedFreeList2_50 <= _GEN_2226;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_51 <= _GEN_9377;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_51 <= _GEN_2227;
        end else begin
          reservedFreeList2_51 <= _GEN_4347;
        end
      end else begin
        reservedFreeList2_51 <= _GEN_2227;
      end
    end else begin
      reservedFreeList2_51 <= _GEN_2227;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_52 <= _GEN_9378;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_52 <= _GEN_2228;
        end else begin
          reservedFreeList2_52 <= _GEN_4348;
        end
      end else begin
        reservedFreeList2_52 <= _GEN_2228;
      end
    end else begin
      reservedFreeList2_52 <= _GEN_2228;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_53 <= _GEN_9379;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_53 <= _GEN_2229;
        end else begin
          reservedFreeList2_53 <= _GEN_4349;
        end
      end else begin
        reservedFreeList2_53 <= _GEN_2229;
      end
    end else begin
      reservedFreeList2_53 <= _GEN_2229;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_54 <= _GEN_9380;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_54 <= _GEN_2230;
        end else begin
          reservedFreeList2_54 <= _GEN_4350;
        end
      end else begin
        reservedFreeList2_54 <= _GEN_2230;
      end
    end else begin
      reservedFreeList2_54 <= _GEN_2230;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_55 <= _GEN_9381;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_55 <= _GEN_2231;
        end else begin
          reservedFreeList2_55 <= _GEN_4351;
        end
      end else begin
        reservedFreeList2_55 <= _GEN_2231;
      end
    end else begin
      reservedFreeList2_55 <= _GEN_2231;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_56 <= _GEN_9382;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_56 <= _GEN_2232;
        end else begin
          reservedFreeList2_56 <= _GEN_4352;
        end
      end else begin
        reservedFreeList2_56 <= _GEN_2232;
      end
    end else begin
      reservedFreeList2_56 <= _GEN_2232;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_57 <= _GEN_9383;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_57 <= _GEN_2233;
        end else begin
          reservedFreeList2_57 <= _GEN_4353;
        end
      end else begin
        reservedFreeList2_57 <= _GEN_2233;
      end
    end else begin
      reservedFreeList2_57 <= _GEN_2233;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_58 <= _GEN_9384;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_58 <= _GEN_2234;
        end else begin
          reservedFreeList2_58 <= _GEN_4354;
        end
      end else begin
        reservedFreeList2_58 <= _GEN_2234;
      end
    end else begin
      reservedFreeList2_58 <= _GEN_2234;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_59 <= _GEN_9385;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_59 <= _GEN_2235;
        end else begin
          reservedFreeList2_59 <= _GEN_4355;
        end
      end else begin
        reservedFreeList2_59 <= _GEN_2235;
      end
    end else begin
      reservedFreeList2_59 <= _GEN_2235;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_60 <= _GEN_9386;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_60 <= _GEN_2236;
        end else begin
          reservedFreeList2_60 <= _GEN_4356;
        end
      end else begin
        reservedFreeList2_60 <= _GEN_2236;
      end
    end else begin
      reservedFreeList2_60 <= _GEN_2236;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_61 <= _GEN_9387;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_61 <= _GEN_2237;
        end else begin
          reservedFreeList2_61 <= _GEN_4357;
        end
      end else begin
        reservedFreeList2_61 <= _GEN_2237;
      end
    end else begin
      reservedFreeList2_61 <= _GEN_2237;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList2_62 <= _GEN_9388;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList2_62 <= _GEN_2238;
        end else begin
          reservedFreeList2_62 <= _GEN_4358;
        end
      end else begin
        reservedFreeList2_62 <= _GEN_2238;
      end
    end else begin
      reservedFreeList2_62 <= _GEN_2238;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_0 <= _GEN_9390;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_0 <= _GEN_2240;
        end else begin
          reservedFreeList3_0 <= _GEN_4456;
        end
      end else begin
        reservedFreeList3_0 <= _GEN_2240;
      end
    end else begin
      reservedFreeList3_0 <= _GEN_2240;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_1 <= _GEN_9391;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_1 <= _GEN_2241;
        end else begin
          reservedFreeList3_1 <= _GEN_4457;
        end
      end else begin
        reservedFreeList3_1 <= _GEN_2241;
      end
    end else begin
      reservedFreeList3_1 <= _GEN_2241;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_2 <= _GEN_9392;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_2 <= _GEN_2242;
        end else begin
          reservedFreeList3_2 <= _GEN_4458;
        end
      end else begin
        reservedFreeList3_2 <= _GEN_2242;
      end
    end else begin
      reservedFreeList3_2 <= _GEN_2242;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_3 <= _GEN_9393;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_3 <= _GEN_2243;
        end else begin
          reservedFreeList3_3 <= _GEN_4459;
        end
      end else begin
        reservedFreeList3_3 <= _GEN_2243;
      end
    end else begin
      reservedFreeList3_3 <= _GEN_2243;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_4 <= _GEN_9394;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_4 <= _GEN_2244;
        end else begin
          reservedFreeList3_4 <= _GEN_4460;
        end
      end else begin
        reservedFreeList3_4 <= _GEN_2244;
      end
    end else begin
      reservedFreeList3_4 <= _GEN_2244;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_5 <= _GEN_9395;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_5 <= _GEN_2245;
        end else begin
          reservedFreeList3_5 <= _GEN_4461;
        end
      end else begin
        reservedFreeList3_5 <= _GEN_2245;
      end
    end else begin
      reservedFreeList3_5 <= _GEN_2245;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_6 <= _GEN_9396;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_6 <= _GEN_2246;
        end else begin
          reservedFreeList3_6 <= _GEN_4462;
        end
      end else begin
        reservedFreeList3_6 <= _GEN_2246;
      end
    end else begin
      reservedFreeList3_6 <= _GEN_2246;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_7 <= _GEN_9397;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_7 <= _GEN_2247;
        end else begin
          reservedFreeList3_7 <= _GEN_4463;
        end
      end else begin
        reservedFreeList3_7 <= _GEN_2247;
      end
    end else begin
      reservedFreeList3_7 <= _GEN_2247;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_8 <= _GEN_9398;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_8 <= _GEN_2248;
        end else begin
          reservedFreeList3_8 <= _GEN_4464;
        end
      end else begin
        reservedFreeList3_8 <= _GEN_2248;
      end
    end else begin
      reservedFreeList3_8 <= _GEN_2248;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_9 <= _GEN_9399;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_9 <= _GEN_2249;
        end else begin
          reservedFreeList3_9 <= _GEN_4465;
        end
      end else begin
        reservedFreeList3_9 <= _GEN_2249;
      end
    end else begin
      reservedFreeList3_9 <= _GEN_2249;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_10 <= _GEN_9400;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_10 <= _GEN_2250;
        end else begin
          reservedFreeList3_10 <= _GEN_4466;
        end
      end else begin
        reservedFreeList3_10 <= _GEN_2250;
      end
    end else begin
      reservedFreeList3_10 <= _GEN_2250;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_11 <= _GEN_9401;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_11 <= _GEN_2251;
        end else begin
          reservedFreeList3_11 <= _GEN_4467;
        end
      end else begin
        reservedFreeList3_11 <= _GEN_2251;
      end
    end else begin
      reservedFreeList3_11 <= _GEN_2251;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_12 <= _GEN_9402;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_12 <= _GEN_2252;
        end else begin
          reservedFreeList3_12 <= _GEN_4468;
        end
      end else begin
        reservedFreeList3_12 <= _GEN_2252;
      end
    end else begin
      reservedFreeList3_12 <= _GEN_2252;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_13 <= _GEN_9403;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_13 <= _GEN_2253;
        end else begin
          reservedFreeList3_13 <= _GEN_4469;
        end
      end else begin
        reservedFreeList3_13 <= _GEN_2253;
      end
    end else begin
      reservedFreeList3_13 <= _GEN_2253;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_14 <= _GEN_9404;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_14 <= _GEN_2254;
        end else begin
          reservedFreeList3_14 <= _GEN_4470;
        end
      end else begin
        reservedFreeList3_14 <= _GEN_2254;
      end
    end else begin
      reservedFreeList3_14 <= _GEN_2254;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_15 <= _GEN_9405;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_15 <= _GEN_2255;
        end else begin
          reservedFreeList3_15 <= _GEN_4471;
        end
      end else begin
        reservedFreeList3_15 <= _GEN_2255;
      end
    end else begin
      reservedFreeList3_15 <= _GEN_2255;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_16 <= _GEN_9406;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_16 <= _GEN_2256;
        end else begin
          reservedFreeList3_16 <= _GEN_4472;
        end
      end else begin
        reservedFreeList3_16 <= _GEN_2256;
      end
    end else begin
      reservedFreeList3_16 <= _GEN_2256;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_17 <= _GEN_9407;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_17 <= _GEN_2257;
        end else begin
          reservedFreeList3_17 <= _GEN_4473;
        end
      end else begin
        reservedFreeList3_17 <= _GEN_2257;
      end
    end else begin
      reservedFreeList3_17 <= _GEN_2257;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_18 <= _GEN_9408;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_18 <= _GEN_2258;
        end else begin
          reservedFreeList3_18 <= _GEN_4474;
        end
      end else begin
        reservedFreeList3_18 <= _GEN_2258;
      end
    end else begin
      reservedFreeList3_18 <= _GEN_2258;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_19 <= _GEN_9409;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_19 <= _GEN_2259;
        end else begin
          reservedFreeList3_19 <= _GEN_4475;
        end
      end else begin
        reservedFreeList3_19 <= _GEN_2259;
      end
    end else begin
      reservedFreeList3_19 <= _GEN_2259;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_20 <= _GEN_9410;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_20 <= _GEN_2260;
        end else begin
          reservedFreeList3_20 <= _GEN_4476;
        end
      end else begin
        reservedFreeList3_20 <= _GEN_2260;
      end
    end else begin
      reservedFreeList3_20 <= _GEN_2260;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_21 <= _GEN_9411;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_21 <= _GEN_2261;
        end else begin
          reservedFreeList3_21 <= _GEN_4477;
        end
      end else begin
        reservedFreeList3_21 <= _GEN_2261;
      end
    end else begin
      reservedFreeList3_21 <= _GEN_2261;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_22 <= _GEN_9412;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_22 <= _GEN_2262;
        end else begin
          reservedFreeList3_22 <= _GEN_4478;
        end
      end else begin
        reservedFreeList3_22 <= _GEN_2262;
      end
    end else begin
      reservedFreeList3_22 <= _GEN_2262;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_23 <= _GEN_9413;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_23 <= _GEN_2263;
        end else begin
          reservedFreeList3_23 <= _GEN_4479;
        end
      end else begin
        reservedFreeList3_23 <= _GEN_2263;
      end
    end else begin
      reservedFreeList3_23 <= _GEN_2263;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_24 <= _GEN_9414;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_24 <= _GEN_2264;
        end else begin
          reservedFreeList3_24 <= _GEN_4480;
        end
      end else begin
        reservedFreeList3_24 <= _GEN_2264;
      end
    end else begin
      reservedFreeList3_24 <= _GEN_2264;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_25 <= _GEN_9415;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_25 <= _GEN_2265;
        end else begin
          reservedFreeList3_25 <= _GEN_4481;
        end
      end else begin
        reservedFreeList3_25 <= _GEN_2265;
      end
    end else begin
      reservedFreeList3_25 <= _GEN_2265;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_26 <= _GEN_9416;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_26 <= _GEN_2266;
        end else begin
          reservedFreeList3_26 <= _GEN_4482;
        end
      end else begin
        reservedFreeList3_26 <= _GEN_2266;
      end
    end else begin
      reservedFreeList3_26 <= _GEN_2266;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_27 <= _GEN_9417;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_27 <= _GEN_2267;
        end else begin
          reservedFreeList3_27 <= _GEN_4483;
        end
      end else begin
        reservedFreeList3_27 <= _GEN_2267;
      end
    end else begin
      reservedFreeList3_27 <= _GEN_2267;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_28 <= _GEN_9418;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_28 <= _GEN_2268;
        end else begin
          reservedFreeList3_28 <= _GEN_4484;
        end
      end else begin
        reservedFreeList3_28 <= _GEN_2268;
      end
    end else begin
      reservedFreeList3_28 <= _GEN_2268;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_29 <= _GEN_9419;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_29 <= _GEN_2269;
        end else begin
          reservedFreeList3_29 <= _GEN_4485;
        end
      end else begin
        reservedFreeList3_29 <= _GEN_2269;
      end
    end else begin
      reservedFreeList3_29 <= _GEN_2269;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_30 <= _GEN_9420;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_30 <= _GEN_2270;
        end else begin
          reservedFreeList3_30 <= _GEN_4486;
        end
      end else begin
        reservedFreeList3_30 <= _GEN_2270;
      end
    end else begin
      reservedFreeList3_30 <= _GEN_2270;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_31 <= _GEN_9421;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_31 <= _GEN_2271;
        end else begin
          reservedFreeList3_31 <= _GEN_4487;
        end
      end else begin
        reservedFreeList3_31 <= _GEN_2271;
      end
    end else begin
      reservedFreeList3_31 <= _GEN_2271;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_32 <= _GEN_9422;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_32 <= _GEN_2272;
        end else begin
          reservedFreeList3_32 <= _GEN_4488;
        end
      end else begin
        reservedFreeList3_32 <= _GEN_2272;
      end
    end else begin
      reservedFreeList3_32 <= _GEN_2272;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_33 <= _GEN_9423;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_33 <= _GEN_2273;
        end else begin
          reservedFreeList3_33 <= _GEN_4489;
        end
      end else begin
        reservedFreeList3_33 <= _GEN_2273;
      end
    end else begin
      reservedFreeList3_33 <= _GEN_2273;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_34 <= _GEN_9424;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_34 <= _GEN_2274;
        end else begin
          reservedFreeList3_34 <= _GEN_4490;
        end
      end else begin
        reservedFreeList3_34 <= _GEN_2274;
      end
    end else begin
      reservedFreeList3_34 <= _GEN_2274;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_35 <= _GEN_9425;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_35 <= _GEN_2275;
        end else begin
          reservedFreeList3_35 <= _GEN_4491;
        end
      end else begin
        reservedFreeList3_35 <= _GEN_2275;
      end
    end else begin
      reservedFreeList3_35 <= _GEN_2275;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_36 <= _GEN_9426;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_36 <= _GEN_2276;
        end else begin
          reservedFreeList3_36 <= _GEN_4492;
        end
      end else begin
        reservedFreeList3_36 <= _GEN_2276;
      end
    end else begin
      reservedFreeList3_36 <= _GEN_2276;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_37 <= _GEN_9427;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_37 <= _GEN_2277;
        end else begin
          reservedFreeList3_37 <= _GEN_4493;
        end
      end else begin
        reservedFreeList3_37 <= _GEN_2277;
      end
    end else begin
      reservedFreeList3_37 <= _GEN_2277;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_38 <= _GEN_9428;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_38 <= _GEN_2278;
        end else begin
          reservedFreeList3_38 <= _GEN_4494;
        end
      end else begin
        reservedFreeList3_38 <= _GEN_2278;
      end
    end else begin
      reservedFreeList3_38 <= _GEN_2278;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_39 <= _GEN_9429;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_39 <= _GEN_2279;
        end else begin
          reservedFreeList3_39 <= _GEN_4495;
        end
      end else begin
        reservedFreeList3_39 <= _GEN_2279;
      end
    end else begin
      reservedFreeList3_39 <= _GEN_2279;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_40 <= _GEN_9430;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_40 <= _GEN_2280;
        end else begin
          reservedFreeList3_40 <= _GEN_4496;
        end
      end else begin
        reservedFreeList3_40 <= _GEN_2280;
      end
    end else begin
      reservedFreeList3_40 <= _GEN_2280;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_41 <= _GEN_9431;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_41 <= _GEN_2281;
        end else begin
          reservedFreeList3_41 <= _GEN_4497;
        end
      end else begin
        reservedFreeList3_41 <= _GEN_2281;
      end
    end else begin
      reservedFreeList3_41 <= _GEN_2281;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_42 <= _GEN_9432;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_42 <= _GEN_2282;
        end else begin
          reservedFreeList3_42 <= _GEN_4498;
        end
      end else begin
        reservedFreeList3_42 <= _GEN_2282;
      end
    end else begin
      reservedFreeList3_42 <= _GEN_2282;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_43 <= _GEN_9433;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_43 <= _GEN_2283;
        end else begin
          reservedFreeList3_43 <= _GEN_4499;
        end
      end else begin
        reservedFreeList3_43 <= _GEN_2283;
      end
    end else begin
      reservedFreeList3_43 <= _GEN_2283;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_44 <= _GEN_9434;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_44 <= _GEN_2284;
        end else begin
          reservedFreeList3_44 <= _GEN_4500;
        end
      end else begin
        reservedFreeList3_44 <= _GEN_2284;
      end
    end else begin
      reservedFreeList3_44 <= _GEN_2284;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_45 <= _GEN_9435;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_45 <= _GEN_2285;
        end else begin
          reservedFreeList3_45 <= _GEN_4501;
        end
      end else begin
        reservedFreeList3_45 <= _GEN_2285;
      end
    end else begin
      reservedFreeList3_45 <= _GEN_2285;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_46 <= _GEN_9436;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_46 <= _GEN_2286;
        end else begin
          reservedFreeList3_46 <= _GEN_4502;
        end
      end else begin
        reservedFreeList3_46 <= _GEN_2286;
      end
    end else begin
      reservedFreeList3_46 <= _GEN_2286;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_47 <= _GEN_9437;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_47 <= _GEN_2287;
        end else begin
          reservedFreeList3_47 <= _GEN_4503;
        end
      end else begin
        reservedFreeList3_47 <= _GEN_2287;
      end
    end else begin
      reservedFreeList3_47 <= _GEN_2287;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_48 <= _GEN_9438;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_48 <= _GEN_2288;
        end else begin
          reservedFreeList3_48 <= _GEN_4504;
        end
      end else begin
        reservedFreeList3_48 <= _GEN_2288;
      end
    end else begin
      reservedFreeList3_48 <= _GEN_2288;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_49 <= _GEN_9439;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_49 <= _GEN_2289;
        end else begin
          reservedFreeList3_49 <= _GEN_4505;
        end
      end else begin
        reservedFreeList3_49 <= _GEN_2289;
      end
    end else begin
      reservedFreeList3_49 <= _GEN_2289;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_50 <= _GEN_9440;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_50 <= _GEN_2290;
        end else begin
          reservedFreeList3_50 <= _GEN_4506;
        end
      end else begin
        reservedFreeList3_50 <= _GEN_2290;
      end
    end else begin
      reservedFreeList3_50 <= _GEN_2290;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_51 <= _GEN_9441;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_51 <= _GEN_2291;
        end else begin
          reservedFreeList3_51 <= _GEN_4507;
        end
      end else begin
        reservedFreeList3_51 <= _GEN_2291;
      end
    end else begin
      reservedFreeList3_51 <= _GEN_2291;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_52 <= _GEN_9442;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_52 <= _GEN_2292;
        end else begin
          reservedFreeList3_52 <= _GEN_4508;
        end
      end else begin
        reservedFreeList3_52 <= _GEN_2292;
      end
    end else begin
      reservedFreeList3_52 <= _GEN_2292;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_53 <= _GEN_9443;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_53 <= _GEN_2293;
        end else begin
          reservedFreeList3_53 <= _GEN_4509;
        end
      end else begin
        reservedFreeList3_53 <= _GEN_2293;
      end
    end else begin
      reservedFreeList3_53 <= _GEN_2293;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_54 <= _GEN_9444;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_54 <= _GEN_2294;
        end else begin
          reservedFreeList3_54 <= _GEN_4510;
        end
      end else begin
        reservedFreeList3_54 <= _GEN_2294;
      end
    end else begin
      reservedFreeList3_54 <= _GEN_2294;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_55 <= _GEN_9445;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_55 <= _GEN_2295;
        end else begin
          reservedFreeList3_55 <= _GEN_4511;
        end
      end else begin
        reservedFreeList3_55 <= _GEN_2295;
      end
    end else begin
      reservedFreeList3_55 <= _GEN_2295;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_56 <= _GEN_9446;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_56 <= _GEN_2296;
        end else begin
          reservedFreeList3_56 <= _GEN_4512;
        end
      end else begin
        reservedFreeList3_56 <= _GEN_2296;
      end
    end else begin
      reservedFreeList3_56 <= _GEN_2296;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_57 <= _GEN_9447;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_57 <= _GEN_2297;
        end else begin
          reservedFreeList3_57 <= _GEN_4513;
        end
      end else begin
        reservedFreeList3_57 <= _GEN_2297;
      end
    end else begin
      reservedFreeList3_57 <= _GEN_2297;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_58 <= _GEN_9448;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_58 <= _GEN_2298;
        end else begin
          reservedFreeList3_58 <= _GEN_4514;
        end
      end else begin
        reservedFreeList3_58 <= _GEN_2298;
      end
    end else begin
      reservedFreeList3_58 <= _GEN_2298;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_59 <= _GEN_9449;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_59 <= _GEN_2299;
        end else begin
          reservedFreeList3_59 <= _GEN_4515;
        end
      end else begin
        reservedFreeList3_59 <= _GEN_2299;
      end
    end else begin
      reservedFreeList3_59 <= _GEN_2299;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_60 <= _GEN_9450;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_60 <= _GEN_2300;
        end else begin
          reservedFreeList3_60 <= _GEN_4516;
        end
      end else begin
        reservedFreeList3_60 <= _GEN_2300;
      end
    end else begin
      reservedFreeList3_60 <= _GEN_2300;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_61 <= _GEN_9451;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_61 <= _GEN_2301;
        end else begin
          reservedFreeList3_61 <= _GEN_4517;
        end
      end else begin
        reservedFreeList3_61 <= _GEN_2301;
      end
    end else begin
      reservedFreeList3_61 <= _GEN_2301;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList3_62 <= _GEN_9452;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedFreeList3_62 <= _GEN_2302;
        end else begin
          reservedFreeList3_62 <= _GEN_4518;
        end
      end else begin
        reservedFreeList3_62 <= _GEN_2302;
      end
    end else begin
      reservedFreeList3_62 <= _GEN_2302;
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_0 <= _GEN_9454;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_0 <= _GEN_4616;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_1 <= _GEN_9455;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_1 <= _GEN_4617;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_2 <= _GEN_9456;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_2 <= _GEN_4618;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_3 <= _GEN_9457;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_3 <= _GEN_4619;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_4 <= _GEN_9458;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_4 <= _GEN_4620;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_5 <= _GEN_9459;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_5 <= _GEN_4621;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_6 <= _GEN_9460;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_6 <= _GEN_4622;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_7 <= _GEN_9461;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_7 <= _GEN_4623;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_8 <= _GEN_9462;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_8 <= _GEN_4624;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_9 <= _GEN_9463;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_9 <= _GEN_4625;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_10 <= _GEN_9464;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_10 <= _GEN_4626;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_11 <= _GEN_9465;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_11 <= _GEN_4627;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_12 <= _GEN_9466;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_12 <= _GEN_4628;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_13 <= _GEN_9467;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_13 <= _GEN_4629;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_14 <= _GEN_9468;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_14 <= _GEN_4630;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_15 <= _GEN_9469;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_15 <= _GEN_4631;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_16 <= _GEN_9470;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_16 <= _GEN_4632;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_17 <= _GEN_9471;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_17 <= _GEN_4633;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_18 <= _GEN_9472;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_18 <= _GEN_4634;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_19 <= _GEN_9473;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_19 <= _GEN_4635;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_20 <= _GEN_9474;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_20 <= _GEN_4636;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_21 <= _GEN_9475;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_21 <= _GEN_4637;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_22 <= _GEN_9476;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_22 <= _GEN_4638;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_23 <= _GEN_9477;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_23 <= _GEN_4639;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_24 <= _GEN_9478;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_24 <= _GEN_4640;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_25 <= _GEN_9479;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_25 <= _GEN_4641;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_26 <= _GEN_9480;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_26 <= _GEN_4642;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_27 <= _GEN_9481;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_27 <= _GEN_4643;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_28 <= _GEN_9482;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_28 <= _GEN_4644;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_29 <= _GEN_9483;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_29 <= _GEN_4645;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_30 <= _GEN_9484;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_30 <= _GEN_4646;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_31 <= _GEN_9485;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_31 <= _GEN_4647;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_32 <= _GEN_9486;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_32 <= _GEN_4648;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_33 <= _GEN_9487;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_33 <= _GEN_4649;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_34 <= _GEN_9488;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_34 <= _GEN_4650;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_35 <= _GEN_9489;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_35 <= _GEN_4651;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_36 <= _GEN_9490;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_36 <= _GEN_4652;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_37 <= _GEN_9491;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_37 <= _GEN_4653;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_38 <= _GEN_9492;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_38 <= _GEN_4654;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_39 <= _GEN_9493;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_39 <= _GEN_4655;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_40 <= _GEN_9494;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_40 <= _GEN_4656;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_41 <= _GEN_9495;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_41 <= _GEN_4657;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_42 <= _GEN_9496;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_42 <= _GEN_4658;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_43 <= _GEN_9497;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_43 <= _GEN_4659;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_44 <= _GEN_9498;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_44 <= _GEN_4660;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_45 <= _GEN_9499;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_45 <= _GEN_4661;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_46 <= _GEN_9500;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_46 <= _GEN_4662;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_47 <= _GEN_9501;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_47 <= _GEN_4663;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_48 <= _GEN_9502;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_48 <= _GEN_4664;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_49 <= _GEN_9503;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_49 <= _GEN_4665;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_50 <= _GEN_9504;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_50 <= _GEN_4666;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_51 <= _GEN_9505;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_51 <= _GEN_4667;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_52 <= _GEN_9506;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_52 <= _GEN_4668;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_53 <= _GEN_9507;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_53 <= _GEN_4669;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_54 <= _GEN_9508;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_54 <= _GEN_4670;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_55 <= _GEN_9509;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_55 <= _GEN_4671;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_56 <= _GEN_9510;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_56 <= _GEN_4672;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_57 <= _GEN_9511;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_57 <= _GEN_4673;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_58 <= _GEN_9512;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_58 <= _GEN_4674;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_59 <= _GEN_9513;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_59 <= _GEN_4675;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_60 <= _GEN_9514;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_60 <= _GEN_4676;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_61 <= _GEN_9515;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_61 <= _GEN_4677;
        end
      end
    end
    if (_T_464) begin // @[decode.scala 856:5]
      reservedFreeList4_62 <= _GEN_9516;
    end else if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          reservedFreeList4_62 <= _GEN_4678;
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_0 <= _GEN_2600;
          end else begin
            reservedValidList1_0 <= PRFValidList_0; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_0 <= _GEN_2304;
        end
      end else begin
        reservedValidList1_0 <= _GEN_2304;
      end
    end else begin
      reservedValidList1_0 <= _GEN_2304;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_1 <= _GEN_2601;
          end else begin
            reservedValidList1_1 <= PRFValidList_1; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_1 <= _GEN_2305;
        end
      end else begin
        reservedValidList1_1 <= _GEN_2305;
      end
    end else begin
      reservedValidList1_1 <= _GEN_2305;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_2 <= _GEN_2602;
          end else begin
            reservedValidList1_2 <= PRFValidList_2; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_2 <= _GEN_2306;
        end
      end else begin
        reservedValidList1_2 <= _GEN_2306;
      end
    end else begin
      reservedValidList1_2 <= _GEN_2306;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_3 <= _GEN_2603;
          end else begin
            reservedValidList1_3 <= PRFValidList_3; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_3 <= _GEN_2307;
        end
      end else begin
        reservedValidList1_3 <= _GEN_2307;
      end
    end else begin
      reservedValidList1_3 <= _GEN_2307;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_4 <= _GEN_2604;
          end else begin
            reservedValidList1_4 <= PRFValidList_4; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_4 <= _GEN_2308;
        end
      end else begin
        reservedValidList1_4 <= _GEN_2308;
      end
    end else begin
      reservedValidList1_4 <= _GEN_2308;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_5 <= _GEN_2605;
          end else begin
            reservedValidList1_5 <= PRFValidList_5; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_5 <= _GEN_2309;
        end
      end else begin
        reservedValidList1_5 <= _GEN_2309;
      end
    end else begin
      reservedValidList1_5 <= _GEN_2309;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_6 <= _GEN_2606;
          end else begin
            reservedValidList1_6 <= PRFValidList_6; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_6 <= _GEN_2310;
        end
      end else begin
        reservedValidList1_6 <= _GEN_2310;
      end
    end else begin
      reservedValidList1_6 <= _GEN_2310;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_7 <= _GEN_2607;
          end else begin
            reservedValidList1_7 <= PRFValidList_7; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_7 <= _GEN_2311;
        end
      end else begin
        reservedValidList1_7 <= _GEN_2311;
      end
    end else begin
      reservedValidList1_7 <= _GEN_2311;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_8 <= _GEN_2608;
          end else begin
            reservedValidList1_8 <= PRFValidList_8; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_8 <= _GEN_2312;
        end
      end else begin
        reservedValidList1_8 <= _GEN_2312;
      end
    end else begin
      reservedValidList1_8 <= _GEN_2312;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_9 <= _GEN_2609;
          end else begin
            reservedValidList1_9 <= PRFValidList_9; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_9 <= _GEN_2313;
        end
      end else begin
        reservedValidList1_9 <= _GEN_2313;
      end
    end else begin
      reservedValidList1_9 <= _GEN_2313;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_10 <= _GEN_2610;
          end else begin
            reservedValidList1_10 <= PRFValidList_10; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_10 <= _GEN_2314;
        end
      end else begin
        reservedValidList1_10 <= _GEN_2314;
      end
    end else begin
      reservedValidList1_10 <= _GEN_2314;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_11 <= _GEN_2611;
          end else begin
            reservedValidList1_11 <= PRFValidList_11; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_11 <= _GEN_2315;
        end
      end else begin
        reservedValidList1_11 <= _GEN_2315;
      end
    end else begin
      reservedValidList1_11 <= _GEN_2315;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_12 <= _GEN_2612;
          end else begin
            reservedValidList1_12 <= PRFValidList_12; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_12 <= _GEN_2316;
        end
      end else begin
        reservedValidList1_12 <= _GEN_2316;
      end
    end else begin
      reservedValidList1_12 <= _GEN_2316;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_13 <= _GEN_2613;
          end else begin
            reservedValidList1_13 <= PRFValidList_13; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_13 <= _GEN_2317;
        end
      end else begin
        reservedValidList1_13 <= _GEN_2317;
      end
    end else begin
      reservedValidList1_13 <= _GEN_2317;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_14 <= _GEN_2614;
          end else begin
            reservedValidList1_14 <= PRFValidList_14; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_14 <= _GEN_2318;
        end
      end else begin
        reservedValidList1_14 <= _GEN_2318;
      end
    end else begin
      reservedValidList1_14 <= _GEN_2318;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_15 <= _GEN_2615;
          end else begin
            reservedValidList1_15 <= PRFValidList_15; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_15 <= _GEN_2319;
        end
      end else begin
        reservedValidList1_15 <= _GEN_2319;
      end
    end else begin
      reservedValidList1_15 <= _GEN_2319;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_16 <= _GEN_2616;
          end else begin
            reservedValidList1_16 <= PRFValidList_16; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_16 <= _GEN_2320;
        end
      end else begin
        reservedValidList1_16 <= _GEN_2320;
      end
    end else begin
      reservedValidList1_16 <= _GEN_2320;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_17 <= _GEN_2617;
          end else begin
            reservedValidList1_17 <= PRFValidList_17; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_17 <= _GEN_2321;
        end
      end else begin
        reservedValidList1_17 <= _GEN_2321;
      end
    end else begin
      reservedValidList1_17 <= _GEN_2321;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_18 <= _GEN_2618;
          end else begin
            reservedValidList1_18 <= PRFValidList_18; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_18 <= _GEN_2322;
        end
      end else begin
        reservedValidList1_18 <= _GEN_2322;
      end
    end else begin
      reservedValidList1_18 <= _GEN_2322;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_19 <= _GEN_2619;
          end else begin
            reservedValidList1_19 <= PRFValidList_19; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_19 <= _GEN_2323;
        end
      end else begin
        reservedValidList1_19 <= _GEN_2323;
      end
    end else begin
      reservedValidList1_19 <= _GEN_2323;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_20 <= _GEN_2620;
          end else begin
            reservedValidList1_20 <= PRFValidList_20; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_20 <= _GEN_2324;
        end
      end else begin
        reservedValidList1_20 <= _GEN_2324;
      end
    end else begin
      reservedValidList1_20 <= _GEN_2324;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_21 <= _GEN_2621;
          end else begin
            reservedValidList1_21 <= PRFValidList_21; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_21 <= _GEN_2325;
        end
      end else begin
        reservedValidList1_21 <= _GEN_2325;
      end
    end else begin
      reservedValidList1_21 <= _GEN_2325;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_22 <= _GEN_2622;
          end else begin
            reservedValidList1_22 <= PRFValidList_22; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_22 <= _GEN_2326;
        end
      end else begin
        reservedValidList1_22 <= _GEN_2326;
      end
    end else begin
      reservedValidList1_22 <= _GEN_2326;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_23 <= _GEN_2623;
          end else begin
            reservedValidList1_23 <= PRFValidList_23; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_23 <= _GEN_2327;
        end
      end else begin
        reservedValidList1_23 <= _GEN_2327;
      end
    end else begin
      reservedValidList1_23 <= _GEN_2327;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_24 <= _GEN_2624;
          end else begin
            reservedValidList1_24 <= PRFValidList_24; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_24 <= _GEN_2328;
        end
      end else begin
        reservedValidList1_24 <= _GEN_2328;
      end
    end else begin
      reservedValidList1_24 <= _GEN_2328;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_25 <= _GEN_2625;
          end else begin
            reservedValidList1_25 <= PRFValidList_25; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_25 <= _GEN_2329;
        end
      end else begin
        reservedValidList1_25 <= _GEN_2329;
      end
    end else begin
      reservedValidList1_25 <= _GEN_2329;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_26 <= _GEN_2626;
          end else begin
            reservedValidList1_26 <= PRFValidList_26; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_26 <= _GEN_2330;
        end
      end else begin
        reservedValidList1_26 <= _GEN_2330;
      end
    end else begin
      reservedValidList1_26 <= _GEN_2330;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_27 <= _GEN_2627;
          end else begin
            reservedValidList1_27 <= PRFValidList_27; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_27 <= _GEN_2331;
        end
      end else begin
        reservedValidList1_27 <= _GEN_2331;
      end
    end else begin
      reservedValidList1_27 <= _GEN_2331;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_28 <= _GEN_2628;
          end else begin
            reservedValidList1_28 <= PRFValidList_28; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_28 <= _GEN_2332;
        end
      end else begin
        reservedValidList1_28 <= _GEN_2332;
      end
    end else begin
      reservedValidList1_28 <= _GEN_2332;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_29 <= _GEN_2629;
          end else begin
            reservedValidList1_29 <= PRFValidList_29; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_29 <= _GEN_2333;
        end
      end else begin
        reservedValidList1_29 <= _GEN_2333;
      end
    end else begin
      reservedValidList1_29 <= _GEN_2333;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_30 <= _GEN_2630;
          end else begin
            reservedValidList1_30 <= PRFValidList_30; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_30 <= _GEN_2334;
        end
      end else begin
        reservedValidList1_30 <= _GEN_2334;
      end
    end else begin
      reservedValidList1_30 <= _GEN_2334;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_31 <= _GEN_2631;
          end else begin
            reservedValidList1_31 <= PRFValidList_31; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_31 <= _GEN_2335;
        end
      end else begin
        reservedValidList1_31 <= _GEN_2335;
      end
    end else begin
      reservedValidList1_31 <= _GEN_2335;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_32 <= _GEN_2632;
          end else begin
            reservedValidList1_32 <= PRFValidList_32; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_32 <= _GEN_2336;
        end
      end else begin
        reservedValidList1_32 <= _GEN_2336;
      end
    end else begin
      reservedValidList1_32 <= _GEN_2336;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_33 <= _GEN_2633;
          end else begin
            reservedValidList1_33 <= PRFValidList_33; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_33 <= _GEN_2337;
        end
      end else begin
        reservedValidList1_33 <= _GEN_2337;
      end
    end else begin
      reservedValidList1_33 <= _GEN_2337;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_34 <= _GEN_2634;
          end else begin
            reservedValidList1_34 <= PRFValidList_34; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_34 <= _GEN_2338;
        end
      end else begin
        reservedValidList1_34 <= _GEN_2338;
      end
    end else begin
      reservedValidList1_34 <= _GEN_2338;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_35 <= _GEN_2635;
          end else begin
            reservedValidList1_35 <= PRFValidList_35; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_35 <= _GEN_2339;
        end
      end else begin
        reservedValidList1_35 <= _GEN_2339;
      end
    end else begin
      reservedValidList1_35 <= _GEN_2339;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_36 <= _GEN_2636;
          end else begin
            reservedValidList1_36 <= PRFValidList_36; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_36 <= _GEN_2340;
        end
      end else begin
        reservedValidList1_36 <= _GEN_2340;
      end
    end else begin
      reservedValidList1_36 <= _GEN_2340;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_37 <= _GEN_2637;
          end else begin
            reservedValidList1_37 <= PRFValidList_37; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_37 <= _GEN_2341;
        end
      end else begin
        reservedValidList1_37 <= _GEN_2341;
      end
    end else begin
      reservedValidList1_37 <= _GEN_2341;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_38 <= _GEN_2638;
          end else begin
            reservedValidList1_38 <= PRFValidList_38; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_38 <= _GEN_2342;
        end
      end else begin
        reservedValidList1_38 <= _GEN_2342;
      end
    end else begin
      reservedValidList1_38 <= _GEN_2342;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_39 <= _GEN_2639;
          end else begin
            reservedValidList1_39 <= PRFValidList_39; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_39 <= _GEN_2343;
        end
      end else begin
        reservedValidList1_39 <= _GEN_2343;
      end
    end else begin
      reservedValidList1_39 <= _GEN_2343;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_40 <= _GEN_2640;
          end else begin
            reservedValidList1_40 <= PRFValidList_40; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_40 <= _GEN_2344;
        end
      end else begin
        reservedValidList1_40 <= _GEN_2344;
      end
    end else begin
      reservedValidList1_40 <= _GEN_2344;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_41 <= _GEN_2641;
          end else begin
            reservedValidList1_41 <= PRFValidList_41; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_41 <= _GEN_2345;
        end
      end else begin
        reservedValidList1_41 <= _GEN_2345;
      end
    end else begin
      reservedValidList1_41 <= _GEN_2345;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_42 <= _GEN_2642;
          end else begin
            reservedValidList1_42 <= PRFValidList_42; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_42 <= _GEN_2346;
        end
      end else begin
        reservedValidList1_42 <= _GEN_2346;
      end
    end else begin
      reservedValidList1_42 <= _GEN_2346;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_43 <= _GEN_2643;
          end else begin
            reservedValidList1_43 <= PRFValidList_43; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_43 <= _GEN_2347;
        end
      end else begin
        reservedValidList1_43 <= _GEN_2347;
      end
    end else begin
      reservedValidList1_43 <= _GEN_2347;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_44 <= _GEN_2644;
          end else begin
            reservedValidList1_44 <= PRFValidList_44; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_44 <= _GEN_2348;
        end
      end else begin
        reservedValidList1_44 <= _GEN_2348;
      end
    end else begin
      reservedValidList1_44 <= _GEN_2348;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_45 <= _GEN_2645;
          end else begin
            reservedValidList1_45 <= PRFValidList_45; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_45 <= _GEN_2349;
        end
      end else begin
        reservedValidList1_45 <= _GEN_2349;
      end
    end else begin
      reservedValidList1_45 <= _GEN_2349;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_46 <= _GEN_2646;
          end else begin
            reservedValidList1_46 <= PRFValidList_46; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_46 <= _GEN_2350;
        end
      end else begin
        reservedValidList1_46 <= _GEN_2350;
      end
    end else begin
      reservedValidList1_46 <= _GEN_2350;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_47 <= _GEN_2647;
          end else begin
            reservedValidList1_47 <= PRFValidList_47; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_47 <= _GEN_2351;
        end
      end else begin
        reservedValidList1_47 <= _GEN_2351;
      end
    end else begin
      reservedValidList1_47 <= _GEN_2351;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_48 <= _GEN_2648;
          end else begin
            reservedValidList1_48 <= PRFValidList_48; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_48 <= _GEN_2352;
        end
      end else begin
        reservedValidList1_48 <= _GEN_2352;
      end
    end else begin
      reservedValidList1_48 <= _GEN_2352;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_49 <= _GEN_2649;
          end else begin
            reservedValidList1_49 <= PRFValidList_49; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_49 <= _GEN_2353;
        end
      end else begin
        reservedValidList1_49 <= _GEN_2353;
      end
    end else begin
      reservedValidList1_49 <= _GEN_2353;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_50 <= _GEN_2650;
          end else begin
            reservedValidList1_50 <= PRFValidList_50; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_50 <= _GEN_2354;
        end
      end else begin
        reservedValidList1_50 <= _GEN_2354;
      end
    end else begin
      reservedValidList1_50 <= _GEN_2354;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_51 <= _GEN_2651;
          end else begin
            reservedValidList1_51 <= PRFValidList_51; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_51 <= _GEN_2355;
        end
      end else begin
        reservedValidList1_51 <= _GEN_2355;
      end
    end else begin
      reservedValidList1_51 <= _GEN_2355;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_52 <= _GEN_2652;
          end else begin
            reservedValidList1_52 <= PRFValidList_52; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_52 <= _GEN_2356;
        end
      end else begin
        reservedValidList1_52 <= _GEN_2356;
      end
    end else begin
      reservedValidList1_52 <= _GEN_2356;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_53 <= _GEN_2653;
          end else begin
            reservedValidList1_53 <= PRFValidList_53; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_53 <= _GEN_2357;
        end
      end else begin
        reservedValidList1_53 <= _GEN_2357;
      end
    end else begin
      reservedValidList1_53 <= _GEN_2357;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_54 <= _GEN_2654;
          end else begin
            reservedValidList1_54 <= PRFValidList_54; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_54 <= _GEN_2358;
        end
      end else begin
        reservedValidList1_54 <= _GEN_2358;
      end
    end else begin
      reservedValidList1_54 <= _GEN_2358;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_55 <= _GEN_2655;
          end else begin
            reservedValidList1_55 <= PRFValidList_55; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_55 <= _GEN_2359;
        end
      end else begin
        reservedValidList1_55 <= _GEN_2359;
      end
    end else begin
      reservedValidList1_55 <= _GEN_2359;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_56 <= _GEN_2656;
          end else begin
            reservedValidList1_56 <= PRFValidList_56; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_56 <= _GEN_2360;
        end
      end else begin
        reservedValidList1_56 <= _GEN_2360;
      end
    end else begin
      reservedValidList1_56 <= _GEN_2360;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_57 <= _GEN_2657;
          end else begin
            reservedValidList1_57 <= PRFValidList_57; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_57 <= _GEN_2361;
        end
      end else begin
        reservedValidList1_57 <= _GEN_2361;
      end
    end else begin
      reservedValidList1_57 <= _GEN_2361;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_58 <= _GEN_2658;
          end else begin
            reservedValidList1_58 <= PRFValidList_58; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_58 <= _GEN_2362;
        end
      end else begin
        reservedValidList1_58 <= _GEN_2362;
      end
    end else begin
      reservedValidList1_58 <= _GEN_2362;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_59 <= _GEN_2659;
          end else begin
            reservedValidList1_59 <= PRFValidList_59; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_59 <= _GEN_2363;
        end
      end else begin
        reservedValidList1_59 <= _GEN_2363;
      end
    end else begin
      reservedValidList1_59 <= _GEN_2363;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_60 <= _GEN_2660;
          end else begin
            reservedValidList1_60 <= PRFValidList_60; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_60 <= _GEN_2364;
        end
      end else begin
        reservedValidList1_60 <= _GEN_2364;
      end
    end else begin
      reservedValidList1_60 <= _GEN_2364;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_61 <= _GEN_2661;
          end else begin
            reservedValidList1_61 <= PRFValidList_61; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_61 <= _GEN_2365;
        end
      end else begin
        reservedValidList1_61 <= _GEN_2365;
      end
    end else begin
      reservedValidList1_61 <= _GEN_2365;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_62 <= _GEN_2662;
          end else begin
            reservedValidList1_62 <= PRFValidList_62; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_62 <= _GEN_2366;
        end
      end else begin
        reservedValidList1_62 <= _GEN_2366;
      end
    end else begin
      reservedValidList1_62 <= _GEN_2366;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          if (opcode[2] & |inputBuffer_instruction[11:7]) begin // @[decode.scala 405:44]
            reservedValidList1_63 <= _GEN_2663;
          end else begin
            reservedValidList1_63 <= PRFValidList_63; // @[decode.scala 404:30]
          end
        end else begin
          reservedValidList1_63 <= _GEN_2367;
        end
      end else begin
        reservedValidList1_63 <= _GEN_2367;
      end
    end else begin
      reservedValidList1_63 <= _GEN_2367;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_0 <= _GEN_2368;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_0 <= _GEN_2760;
        end else begin
          reservedValidList2_0 <= _GEN_2368;
        end
      end else begin
        reservedValidList2_0 <= _GEN_2368;
      end
    end else begin
      reservedValidList2_0 <= _GEN_2368;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_1 <= _GEN_2369;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_1 <= _GEN_2761;
        end else begin
          reservedValidList2_1 <= _GEN_2369;
        end
      end else begin
        reservedValidList2_1 <= _GEN_2369;
      end
    end else begin
      reservedValidList2_1 <= _GEN_2369;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_2 <= _GEN_2370;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_2 <= _GEN_2762;
        end else begin
          reservedValidList2_2 <= _GEN_2370;
        end
      end else begin
        reservedValidList2_2 <= _GEN_2370;
      end
    end else begin
      reservedValidList2_2 <= _GEN_2370;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_3 <= _GEN_2371;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_3 <= _GEN_2763;
        end else begin
          reservedValidList2_3 <= _GEN_2371;
        end
      end else begin
        reservedValidList2_3 <= _GEN_2371;
      end
    end else begin
      reservedValidList2_3 <= _GEN_2371;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_4 <= _GEN_2372;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_4 <= _GEN_2764;
        end else begin
          reservedValidList2_4 <= _GEN_2372;
        end
      end else begin
        reservedValidList2_4 <= _GEN_2372;
      end
    end else begin
      reservedValidList2_4 <= _GEN_2372;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_5 <= _GEN_2373;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_5 <= _GEN_2765;
        end else begin
          reservedValidList2_5 <= _GEN_2373;
        end
      end else begin
        reservedValidList2_5 <= _GEN_2373;
      end
    end else begin
      reservedValidList2_5 <= _GEN_2373;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_6 <= _GEN_2374;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_6 <= _GEN_2766;
        end else begin
          reservedValidList2_6 <= _GEN_2374;
        end
      end else begin
        reservedValidList2_6 <= _GEN_2374;
      end
    end else begin
      reservedValidList2_6 <= _GEN_2374;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_7 <= _GEN_2375;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_7 <= _GEN_2767;
        end else begin
          reservedValidList2_7 <= _GEN_2375;
        end
      end else begin
        reservedValidList2_7 <= _GEN_2375;
      end
    end else begin
      reservedValidList2_7 <= _GEN_2375;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_8 <= _GEN_2376;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_8 <= _GEN_2768;
        end else begin
          reservedValidList2_8 <= _GEN_2376;
        end
      end else begin
        reservedValidList2_8 <= _GEN_2376;
      end
    end else begin
      reservedValidList2_8 <= _GEN_2376;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_9 <= _GEN_2377;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_9 <= _GEN_2769;
        end else begin
          reservedValidList2_9 <= _GEN_2377;
        end
      end else begin
        reservedValidList2_9 <= _GEN_2377;
      end
    end else begin
      reservedValidList2_9 <= _GEN_2377;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_10 <= _GEN_2378;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_10 <= _GEN_2770;
        end else begin
          reservedValidList2_10 <= _GEN_2378;
        end
      end else begin
        reservedValidList2_10 <= _GEN_2378;
      end
    end else begin
      reservedValidList2_10 <= _GEN_2378;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_11 <= _GEN_2379;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_11 <= _GEN_2771;
        end else begin
          reservedValidList2_11 <= _GEN_2379;
        end
      end else begin
        reservedValidList2_11 <= _GEN_2379;
      end
    end else begin
      reservedValidList2_11 <= _GEN_2379;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_12 <= _GEN_2380;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_12 <= _GEN_2772;
        end else begin
          reservedValidList2_12 <= _GEN_2380;
        end
      end else begin
        reservedValidList2_12 <= _GEN_2380;
      end
    end else begin
      reservedValidList2_12 <= _GEN_2380;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_13 <= _GEN_2381;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_13 <= _GEN_2773;
        end else begin
          reservedValidList2_13 <= _GEN_2381;
        end
      end else begin
        reservedValidList2_13 <= _GEN_2381;
      end
    end else begin
      reservedValidList2_13 <= _GEN_2381;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_14 <= _GEN_2382;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_14 <= _GEN_2774;
        end else begin
          reservedValidList2_14 <= _GEN_2382;
        end
      end else begin
        reservedValidList2_14 <= _GEN_2382;
      end
    end else begin
      reservedValidList2_14 <= _GEN_2382;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_15 <= _GEN_2383;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_15 <= _GEN_2775;
        end else begin
          reservedValidList2_15 <= _GEN_2383;
        end
      end else begin
        reservedValidList2_15 <= _GEN_2383;
      end
    end else begin
      reservedValidList2_15 <= _GEN_2383;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_16 <= _GEN_2384;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_16 <= _GEN_2776;
        end else begin
          reservedValidList2_16 <= _GEN_2384;
        end
      end else begin
        reservedValidList2_16 <= _GEN_2384;
      end
    end else begin
      reservedValidList2_16 <= _GEN_2384;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_17 <= _GEN_2385;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_17 <= _GEN_2777;
        end else begin
          reservedValidList2_17 <= _GEN_2385;
        end
      end else begin
        reservedValidList2_17 <= _GEN_2385;
      end
    end else begin
      reservedValidList2_17 <= _GEN_2385;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_18 <= _GEN_2386;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_18 <= _GEN_2778;
        end else begin
          reservedValidList2_18 <= _GEN_2386;
        end
      end else begin
        reservedValidList2_18 <= _GEN_2386;
      end
    end else begin
      reservedValidList2_18 <= _GEN_2386;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_19 <= _GEN_2387;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_19 <= _GEN_2779;
        end else begin
          reservedValidList2_19 <= _GEN_2387;
        end
      end else begin
        reservedValidList2_19 <= _GEN_2387;
      end
    end else begin
      reservedValidList2_19 <= _GEN_2387;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_20 <= _GEN_2388;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_20 <= _GEN_2780;
        end else begin
          reservedValidList2_20 <= _GEN_2388;
        end
      end else begin
        reservedValidList2_20 <= _GEN_2388;
      end
    end else begin
      reservedValidList2_20 <= _GEN_2388;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_21 <= _GEN_2389;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_21 <= _GEN_2781;
        end else begin
          reservedValidList2_21 <= _GEN_2389;
        end
      end else begin
        reservedValidList2_21 <= _GEN_2389;
      end
    end else begin
      reservedValidList2_21 <= _GEN_2389;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_22 <= _GEN_2390;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_22 <= _GEN_2782;
        end else begin
          reservedValidList2_22 <= _GEN_2390;
        end
      end else begin
        reservedValidList2_22 <= _GEN_2390;
      end
    end else begin
      reservedValidList2_22 <= _GEN_2390;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_23 <= _GEN_2391;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_23 <= _GEN_2783;
        end else begin
          reservedValidList2_23 <= _GEN_2391;
        end
      end else begin
        reservedValidList2_23 <= _GEN_2391;
      end
    end else begin
      reservedValidList2_23 <= _GEN_2391;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_24 <= _GEN_2392;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_24 <= _GEN_2784;
        end else begin
          reservedValidList2_24 <= _GEN_2392;
        end
      end else begin
        reservedValidList2_24 <= _GEN_2392;
      end
    end else begin
      reservedValidList2_24 <= _GEN_2392;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_25 <= _GEN_2393;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_25 <= _GEN_2785;
        end else begin
          reservedValidList2_25 <= _GEN_2393;
        end
      end else begin
        reservedValidList2_25 <= _GEN_2393;
      end
    end else begin
      reservedValidList2_25 <= _GEN_2393;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_26 <= _GEN_2394;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_26 <= _GEN_2786;
        end else begin
          reservedValidList2_26 <= _GEN_2394;
        end
      end else begin
        reservedValidList2_26 <= _GEN_2394;
      end
    end else begin
      reservedValidList2_26 <= _GEN_2394;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_27 <= _GEN_2395;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_27 <= _GEN_2787;
        end else begin
          reservedValidList2_27 <= _GEN_2395;
        end
      end else begin
        reservedValidList2_27 <= _GEN_2395;
      end
    end else begin
      reservedValidList2_27 <= _GEN_2395;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_28 <= _GEN_2396;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_28 <= _GEN_2788;
        end else begin
          reservedValidList2_28 <= _GEN_2396;
        end
      end else begin
        reservedValidList2_28 <= _GEN_2396;
      end
    end else begin
      reservedValidList2_28 <= _GEN_2396;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_29 <= _GEN_2397;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_29 <= _GEN_2789;
        end else begin
          reservedValidList2_29 <= _GEN_2397;
        end
      end else begin
        reservedValidList2_29 <= _GEN_2397;
      end
    end else begin
      reservedValidList2_29 <= _GEN_2397;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_30 <= _GEN_2398;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_30 <= _GEN_2790;
        end else begin
          reservedValidList2_30 <= _GEN_2398;
        end
      end else begin
        reservedValidList2_30 <= _GEN_2398;
      end
    end else begin
      reservedValidList2_30 <= _GEN_2398;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_31 <= _GEN_2399;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_31 <= _GEN_2791;
        end else begin
          reservedValidList2_31 <= _GEN_2399;
        end
      end else begin
        reservedValidList2_31 <= _GEN_2399;
      end
    end else begin
      reservedValidList2_31 <= _GEN_2399;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_32 <= _GEN_2400;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_32 <= _GEN_2792;
        end else begin
          reservedValidList2_32 <= _GEN_2400;
        end
      end else begin
        reservedValidList2_32 <= _GEN_2400;
      end
    end else begin
      reservedValidList2_32 <= _GEN_2400;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_33 <= _GEN_2401;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_33 <= _GEN_2793;
        end else begin
          reservedValidList2_33 <= _GEN_2401;
        end
      end else begin
        reservedValidList2_33 <= _GEN_2401;
      end
    end else begin
      reservedValidList2_33 <= _GEN_2401;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_34 <= _GEN_2402;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_34 <= _GEN_2794;
        end else begin
          reservedValidList2_34 <= _GEN_2402;
        end
      end else begin
        reservedValidList2_34 <= _GEN_2402;
      end
    end else begin
      reservedValidList2_34 <= _GEN_2402;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_35 <= _GEN_2403;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_35 <= _GEN_2795;
        end else begin
          reservedValidList2_35 <= _GEN_2403;
        end
      end else begin
        reservedValidList2_35 <= _GEN_2403;
      end
    end else begin
      reservedValidList2_35 <= _GEN_2403;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_36 <= _GEN_2404;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_36 <= _GEN_2796;
        end else begin
          reservedValidList2_36 <= _GEN_2404;
        end
      end else begin
        reservedValidList2_36 <= _GEN_2404;
      end
    end else begin
      reservedValidList2_36 <= _GEN_2404;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_37 <= _GEN_2405;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_37 <= _GEN_2797;
        end else begin
          reservedValidList2_37 <= _GEN_2405;
        end
      end else begin
        reservedValidList2_37 <= _GEN_2405;
      end
    end else begin
      reservedValidList2_37 <= _GEN_2405;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_38 <= _GEN_2406;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_38 <= _GEN_2798;
        end else begin
          reservedValidList2_38 <= _GEN_2406;
        end
      end else begin
        reservedValidList2_38 <= _GEN_2406;
      end
    end else begin
      reservedValidList2_38 <= _GEN_2406;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_39 <= _GEN_2407;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_39 <= _GEN_2799;
        end else begin
          reservedValidList2_39 <= _GEN_2407;
        end
      end else begin
        reservedValidList2_39 <= _GEN_2407;
      end
    end else begin
      reservedValidList2_39 <= _GEN_2407;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_40 <= _GEN_2408;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_40 <= _GEN_2800;
        end else begin
          reservedValidList2_40 <= _GEN_2408;
        end
      end else begin
        reservedValidList2_40 <= _GEN_2408;
      end
    end else begin
      reservedValidList2_40 <= _GEN_2408;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_41 <= _GEN_2409;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_41 <= _GEN_2801;
        end else begin
          reservedValidList2_41 <= _GEN_2409;
        end
      end else begin
        reservedValidList2_41 <= _GEN_2409;
      end
    end else begin
      reservedValidList2_41 <= _GEN_2409;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_42 <= _GEN_2410;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_42 <= _GEN_2802;
        end else begin
          reservedValidList2_42 <= _GEN_2410;
        end
      end else begin
        reservedValidList2_42 <= _GEN_2410;
      end
    end else begin
      reservedValidList2_42 <= _GEN_2410;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_43 <= _GEN_2411;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_43 <= _GEN_2803;
        end else begin
          reservedValidList2_43 <= _GEN_2411;
        end
      end else begin
        reservedValidList2_43 <= _GEN_2411;
      end
    end else begin
      reservedValidList2_43 <= _GEN_2411;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_44 <= _GEN_2412;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_44 <= _GEN_2804;
        end else begin
          reservedValidList2_44 <= _GEN_2412;
        end
      end else begin
        reservedValidList2_44 <= _GEN_2412;
      end
    end else begin
      reservedValidList2_44 <= _GEN_2412;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_45 <= _GEN_2413;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_45 <= _GEN_2805;
        end else begin
          reservedValidList2_45 <= _GEN_2413;
        end
      end else begin
        reservedValidList2_45 <= _GEN_2413;
      end
    end else begin
      reservedValidList2_45 <= _GEN_2413;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_46 <= _GEN_2414;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_46 <= _GEN_2806;
        end else begin
          reservedValidList2_46 <= _GEN_2414;
        end
      end else begin
        reservedValidList2_46 <= _GEN_2414;
      end
    end else begin
      reservedValidList2_46 <= _GEN_2414;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_47 <= _GEN_2415;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_47 <= _GEN_2807;
        end else begin
          reservedValidList2_47 <= _GEN_2415;
        end
      end else begin
        reservedValidList2_47 <= _GEN_2415;
      end
    end else begin
      reservedValidList2_47 <= _GEN_2415;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_48 <= _GEN_2416;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_48 <= _GEN_2808;
        end else begin
          reservedValidList2_48 <= _GEN_2416;
        end
      end else begin
        reservedValidList2_48 <= _GEN_2416;
      end
    end else begin
      reservedValidList2_48 <= _GEN_2416;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_49 <= _GEN_2417;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_49 <= _GEN_2809;
        end else begin
          reservedValidList2_49 <= _GEN_2417;
        end
      end else begin
        reservedValidList2_49 <= _GEN_2417;
      end
    end else begin
      reservedValidList2_49 <= _GEN_2417;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_50 <= _GEN_2418;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_50 <= _GEN_2810;
        end else begin
          reservedValidList2_50 <= _GEN_2418;
        end
      end else begin
        reservedValidList2_50 <= _GEN_2418;
      end
    end else begin
      reservedValidList2_50 <= _GEN_2418;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_51 <= _GEN_2419;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_51 <= _GEN_2811;
        end else begin
          reservedValidList2_51 <= _GEN_2419;
        end
      end else begin
        reservedValidList2_51 <= _GEN_2419;
      end
    end else begin
      reservedValidList2_51 <= _GEN_2419;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_52 <= _GEN_2420;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_52 <= _GEN_2812;
        end else begin
          reservedValidList2_52 <= _GEN_2420;
        end
      end else begin
        reservedValidList2_52 <= _GEN_2420;
      end
    end else begin
      reservedValidList2_52 <= _GEN_2420;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_53 <= _GEN_2421;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_53 <= _GEN_2813;
        end else begin
          reservedValidList2_53 <= _GEN_2421;
        end
      end else begin
        reservedValidList2_53 <= _GEN_2421;
      end
    end else begin
      reservedValidList2_53 <= _GEN_2421;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_54 <= _GEN_2422;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_54 <= _GEN_2814;
        end else begin
          reservedValidList2_54 <= _GEN_2422;
        end
      end else begin
        reservedValidList2_54 <= _GEN_2422;
      end
    end else begin
      reservedValidList2_54 <= _GEN_2422;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_55 <= _GEN_2423;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_55 <= _GEN_2815;
        end else begin
          reservedValidList2_55 <= _GEN_2423;
        end
      end else begin
        reservedValidList2_55 <= _GEN_2423;
      end
    end else begin
      reservedValidList2_55 <= _GEN_2423;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_56 <= _GEN_2424;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_56 <= _GEN_2816;
        end else begin
          reservedValidList2_56 <= _GEN_2424;
        end
      end else begin
        reservedValidList2_56 <= _GEN_2424;
      end
    end else begin
      reservedValidList2_56 <= _GEN_2424;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_57 <= _GEN_2425;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_57 <= _GEN_2817;
        end else begin
          reservedValidList2_57 <= _GEN_2425;
        end
      end else begin
        reservedValidList2_57 <= _GEN_2425;
      end
    end else begin
      reservedValidList2_57 <= _GEN_2425;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_58 <= _GEN_2426;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_58 <= _GEN_2818;
        end else begin
          reservedValidList2_58 <= _GEN_2426;
        end
      end else begin
        reservedValidList2_58 <= _GEN_2426;
      end
    end else begin
      reservedValidList2_58 <= _GEN_2426;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_59 <= _GEN_2427;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_59 <= _GEN_2819;
        end else begin
          reservedValidList2_59 <= _GEN_2427;
        end
      end else begin
        reservedValidList2_59 <= _GEN_2427;
      end
    end else begin
      reservedValidList2_59 <= _GEN_2427;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_60 <= _GEN_2428;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_60 <= _GEN_2820;
        end else begin
          reservedValidList2_60 <= _GEN_2428;
        end
      end else begin
        reservedValidList2_60 <= _GEN_2428;
      end
    end else begin
      reservedValidList2_60 <= _GEN_2428;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_61 <= _GEN_2429;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_61 <= _GEN_2821;
        end else begin
          reservedValidList2_61 <= _GEN_2429;
        end
      end else begin
        reservedValidList2_61 <= _GEN_2429;
      end
    end else begin
      reservedValidList2_61 <= _GEN_2429;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_62 <= _GEN_2430;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_62 <= _GEN_2822;
        end else begin
          reservedValidList2_62 <= _GEN_2430;
        end
      end else begin
        reservedValidList2_62 <= _GEN_2430;
      end
    end else begin
      reservedValidList2_62 <= _GEN_2430;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_63 <= _GEN_2431;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList2_63 <= _GEN_2823;
        end else begin
          reservedValidList2_63 <= _GEN_2431;
        end
      end else begin
        reservedValidList2_63 <= _GEN_2431;
      end
    end else begin
      reservedValidList2_63 <= _GEN_2431;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_0 <= _GEN_2432;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_0 <= _GEN_2432;
        end else begin
          reservedValidList3_0 <= _GEN_4040;
        end
      end else begin
        reservedValidList3_0 <= _GEN_2432;
      end
    end else begin
      reservedValidList3_0 <= _GEN_2432;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_1 <= _GEN_2433;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_1 <= _GEN_2433;
        end else begin
          reservedValidList3_1 <= _GEN_4041;
        end
      end else begin
        reservedValidList3_1 <= _GEN_2433;
      end
    end else begin
      reservedValidList3_1 <= _GEN_2433;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_2 <= _GEN_2434;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_2 <= _GEN_2434;
        end else begin
          reservedValidList3_2 <= _GEN_4042;
        end
      end else begin
        reservedValidList3_2 <= _GEN_2434;
      end
    end else begin
      reservedValidList3_2 <= _GEN_2434;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_3 <= _GEN_2435;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_3 <= _GEN_2435;
        end else begin
          reservedValidList3_3 <= _GEN_4043;
        end
      end else begin
        reservedValidList3_3 <= _GEN_2435;
      end
    end else begin
      reservedValidList3_3 <= _GEN_2435;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_4 <= _GEN_2436;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_4 <= _GEN_2436;
        end else begin
          reservedValidList3_4 <= _GEN_4044;
        end
      end else begin
        reservedValidList3_4 <= _GEN_2436;
      end
    end else begin
      reservedValidList3_4 <= _GEN_2436;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_5 <= _GEN_2437;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_5 <= _GEN_2437;
        end else begin
          reservedValidList3_5 <= _GEN_4045;
        end
      end else begin
        reservedValidList3_5 <= _GEN_2437;
      end
    end else begin
      reservedValidList3_5 <= _GEN_2437;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_6 <= _GEN_2438;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_6 <= _GEN_2438;
        end else begin
          reservedValidList3_6 <= _GEN_4046;
        end
      end else begin
        reservedValidList3_6 <= _GEN_2438;
      end
    end else begin
      reservedValidList3_6 <= _GEN_2438;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_7 <= _GEN_2439;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_7 <= _GEN_2439;
        end else begin
          reservedValidList3_7 <= _GEN_4047;
        end
      end else begin
        reservedValidList3_7 <= _GEN_2439;
      end
    end else begin
      reservedValidList3_7 <= _GEN_2439;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_8 <= _GEN_2440;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_8 <= _GEN_2440;
        end else begin
          reservedValidList3_8 <= _GEN_4048;
        end
      end else begin
        reservedValidList3_8 <= _GEN_2440;
      end
    end else begin
      reservedValidList3_8 <= _GEN_2440;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_9 <= _GEN_2441;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_9 <= _GEN_2441;
        end else begin
          reservedValidList3_9 <= _GEN_4049;
        end
      end else begin
        reservedValidList3_9 <= _GEN_2441;
      end
    end else begin
      reservedValidList3_9 <= _GEN_2441;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_10 <= _GEN_2442;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_10 <= _GEN_2442;
        end else begin
          reservedValidList3_10 <= _GEN_4050;
        end
      end else begin
        reservedValidList3_10 <= _GEN_2442;
      end
    end else begin
      reservedValidList3_10 <= _GEN_2442;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_11 <= _GEN_2443;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_11 <= _GEN_2443;
        end else begin
          reservedValidList3_11 <= _GEN_4051;
        end
      end else begin
        reservedValidList3_11 <= _GEN_2443;
      end
    end else begin
      reservedValidList3_11 <= _GEN_2443;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_12 <= _GEN_2444;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_12 <= _GEN_2444;
        end else begin
          reservedValidList3_12 <= _GEN_4052;
        end
      end else begin
        reservedValidList3_12 <= _GEN_2444;
      end
    end else begin
      reservedValidList3_12 <= _GEN_2444;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_13 <= _GEN_2445;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_13 <= _GEN_2445;
        end else begin
          reservedValidList3_13 <= _GEN_4053;
        end
      end else begin
        reservedValidList3_13 <= _GEN_2445;
      end
    end else begin
      reservedValidList3_13 <= _GEN_2445;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_14 <= _GEN_2446;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_14 <= _GEN_2446;
        end else begin
          reservedValidList3_14 <= _GEN_4054;
        end
      end else begin
        reservedValidList3_14 <= _GEN_2446;
      end
    end else begin
      reservedValidList3_14 <= _GEN_2446;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_15 <= _GEN_2447;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_15 <= _GEN_2447;
        end else begin
          reservedValidList3_15 <= _GEN_4055;
        end
      end else begin
        reservedValidList3_15 <= _GEN_2447;
      end
    end else begin
      reservedValidList3_15 <= _GEN_2447;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_16 <= _GEN_2448;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_16 <= _GEN_2448;
        end else begin
          reservedValidList3_16 <= _GEN_4056;
        end
      end else begin
        reservedValidList3_16 <= _GEN_2448;
      end
    end else begin
      reservedValidList3_16 <= _GEN_2448;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_17 <= _GEN_2449;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_17 <= _GEN_2449;
        end else begin
          reservedValidList3_17 <= _GEN_4057;
        end
      end else begin
        reservedValidList3_17 <= _GEN_2449;
      end
    end else begin
      reservedValidList3_17 <= _GEN_2449;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_18 <= _GEN_2450;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_18 <= _GEN_2450;
        end else begin
          reservedValidList3_18 <= _GEN_4058;
        end
      end else begin
        reservedValidList3_18 <= _GEN_2450;
      end
    end else begin
      reservedValidList3_18 <= _GEN_2450;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_19 <= _GEN_2451;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_19 <= _GEN_2451;
        end else begin
          reservedValidList3_19 <= _GEN_4059;
        end
      end else begin
        reservedValidList3_19 <= _GEN_2451;
      end
    end else begin
      reservedValidList3_19 <= _GEN_2451;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_20 <= _GEN_2452;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_20 <= _GEN_2452;
        end else begin
          reservedValidList3_20 <= _GEN_4060;
        end
      end else begin
        reservedValidList3_20 <= _GEN_2452;
      end
    end else begin
      reservedValidList3_20 <= _GEN_2452;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_21 <= _GEN_2453;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_21 <= _GEN_2453;
        end else begin
          reservedValidList3_21 <= _GEN_4061;
        end
      end else begin
        reservedValidList3_21 <= _GEN_2453;
      end
    end else begin
      reservedValidList3_21 <= _GEN_2453;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_22 <= _GEN_2454;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_22 <= _GEN_2454;
        end else begin
          reservedValidList3_22 <= _GEN_4062;
        end
      end else begin
        reservedValidList3_22 <= _GEN_2454;
      end
    end else begin
      reservedValidList3_22 <= _GEN_2454;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_23 <= _GEN_2455;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_23 <= _GEN_2455;
        end else begin
          reservedValidList3_23 <= _GEN_4063;
        end
      end else begin
        reservedValidList3_23 <= _GEN_2455;
      end
    end else begin
      reservedValidList3_23 <= _GEN_2455;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_24 <= _GEN_2456;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_24 <= _GEN_2456;
        end else begin
          reservedValidList3_24 <= _GEN_4064;
        end
      end else begin
        reservedValidList3_24 <= _GEN_2456;
      end
    end else begin
      reservedValidList3_24 <= _GEN_2456;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_25 <= _GEN_2457;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_25 <= _GEN_2457;
        end else begin
          reservedValidList3_25 <= _GEN_4065;
        end
      end else begin
        reservedValidList3_25 <= _GEN_2457;
      end
    end else begin
      reservedValidList3_25 <= _GEN_2457;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_26 <= _GEN_2458;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_26 <= _GEN_2458;
        end else begin
          reservedValidList3_26 <= _GEN_4066;
        end
      end else begin
        reservedValidList3_26 <= _GEN_2458;
      end
    end else begin
      reservedValidList3_26 <= _GEN_2458;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_27 <= _GEN_2459;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_27 <= _GEN_2459;
        end else begin
          reservedValidList3_27 <= _GEN_4067;
        end
      end else begin
        reservedValidList3_27 <= _GEN_2459;
      end
    end else begin
      reservedValidList3_27 <= _GEN_2459;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_28 <= _GEN_2460;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_28 <= _GEN_2460;
        end else begin
          reservedValidList3_28 <= _GEN_4068;
        end
      end else begin
        reservedValidList3_28 <= _GEN_2460;
      end
    end else begin
      reservedValidList3_28 <= _GEN_2460;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_29 <= _GEN_2461;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_29 <= _GEN_2461;
        end else begin
          reservedValidList3_29 <= _GEN_4069;
        end
      end else begin
        reservedValidList3_29 <= _GEN_2461;
      end
    end else begin
      reservedValidList3_29 <= _GEN_2461;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_30 <= _GEN_2462;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_30 <= _GEN_2462;
        end else begin
          reservedValidList3_30 <= _GEN_4070;
        end
      end else begin
        reservedValidList3_30 <= _GEN_2462;
      end
    end else begin
      reservedValidList3_30 <= _GEN_2462;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_31 <= _GEN_2463;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_31 <= _GEN_2463;
        end else begin
          reservedValidList3_31 <= _GEN_4071;
        end
      end else begin
        reservedValidList3_31 <= _GEN_2463;
      end
    end else begin
      reservedValidList3_31 <= _GEN_2463;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_32 <= _GEN_2464;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_32 <= _GEN_2464;
        end else begin
          reservedValidList3_32 <= _GEN_4072;
        end
      end else begin
        reservedValidList3_32 <= _GEN_2464;
      end
    end else begin
      reservedValidList3_32 <= _GEN_2464;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_33 <= _GEN_2465;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_33 <= _GEN_2465;
        end else begin
          reservedValidList3_33 <= _GEN_4073;
        end
      end else begin
        reservedValidList3_33 <= _GEN_2465;
      end
    end else begin
      reservedValidList3_33 <= _GEN_2465;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_34 <= _GEN_2466;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_34 <= _GEN_2466;
        end else begin
          reservedValidList3_34 <= _GEN_4074;
        end
      end else begin
        reservedValidList3_34 <= _GEN_2466;
      end
    end else begin
      reservedValidList3_34 <= _GEN_2466;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_35 <= _GEN_2467;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_35 <= _GEN_2467;
        end else begin
          reservedValidList3_35 <= _GEN_4075;
        end
      end else begin
        reservedValidList3_35 <= _GEN_2467;
      end
    end else begin
      reservedValidList3_35 <= _GEN_2467;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_36 <= _GEN_2468;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_36 <= _GEN_2468;
        end else begin
          reservedValidList3_36 <= _GEN_4076;
        end
      end else begin
        reservedValidList3_36 <= _GEN_2468;
      end
    end else begin
      reservedValidList3_36 <= _GEN_2468;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_37 <= _GEN_2469;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_37 <= _GEN_2469;
        end else begin
          reservedValidList3_37 <= _GEN_4077;
        end
      end else begin
        reservedValidList3_37 <= _GEN_2469;
      end
    end else begin
      reservedValidList3_37 <= _GEN_2469;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_38 <= _GEN_2470;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_38 <= _GEN_2470;
        end else begin
          reservedValidList3_38 <= _GEN_4078;
        end
      end else begin
        reservedValidList3_38 <= _GEN_2470;
      end
    end else begin
      reservedValidList3_38 <= _GEN_2470;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_39 <= _GEN_2471;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_39 <= _GEN_2471;
        end else begin
          reservedValidList3_39 <= _GEN_4079;
        end
      end else begin
        reservedValidList3_39 <= _GEN_2471;
      end
    end else begin
      reservedValidList3_39 <= _GEN_2471;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_40 <= _GEN_2472;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_40 <= _GEN_2472;
        end else begin
          reservedValidList3_40 <= _GEN_4080;
        end
      end else begin
        reservedValidList3_40 <= _GEN_2472;
      end
    end else begin
      reservedValidList3_40 <= _GEN_2472;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_41 <= _GEN_2473;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_41 <= _GEN_2473;
        end else begin
          reservedValidList3_41 <= _GEN_4081;
        end
      end else begin
        reservedValidList3_41 <= _GEN_2473;
      end
    end else begin
      reservedValidList3_41 <= _GEN_2473;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_42 <= _GEN_2474;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_42 <= _GEN_2474;
        end else begin
          reservedValidList3_42 <= _GEN_4082;
        end
      end else begin
        reservedValidList3_42 <= _GEN_2474;
      end
    end else begin
      reservedValidList3_42 <= _GEN_2474;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_43 <= _GEN_2475;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_43 <= _GEN_2475;
        end else begin
          reservedValidList3_43 <= _GEN_4083;
        end
      end else begin
        reservedValidList3_43 <= _GEN_2475;
      end
    end else begin
      reservedValidList3_43 <= _GEN_2475;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_44 <= _GEN_2476;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_44 <= _GEN_2476;
        end else begin
          reservedValidList3_44 <= _GEN_4084;
        end
      end else begin
        reservedValidList3_44 <= _GEN_2476;
      end
    end else begin
      reservedValidList3_44 <= _GEN_2476;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_45 <= _GEN_2477;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_45 <= _GEN_2477;
        end else begin
          reservedValidList3_45 <= _GEN_4085;
        end
      end else begin
        reservedValidList3_45 <= _GEN_2477;
      end
    end else begin
      reservedValidList3_45 <= _GEN_2477;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_46 <= _GEN_2478;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_46 <= _GEN_2478;
        end else begin
          reservedValidList3_46 <= _GEN_4086;
        end
      end else begin
        reservedValidList3_46 <= _GEN_2478;
      end
    end else begin
      reservedValidList3_46 <= _GEN_2478;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_47 <= _GEN_2479;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_47 <= _GEN_2479;
        end else begin
          reservedValidList3_47 <= _GEN_4087;
        end
      end else begin
        reservedValidList3_47 <= _GEN_2479;
      end
    end else begin
      reservedValidList3_47 <= _GEN_2479;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_48 <= _GEN_2480;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_48 <= _GEN_2480;
        end else begin
          reservedValidList3_48 <= _GEN_4088;
        end
      end else begin
        reservedValidList3_48 <= _GEN_2480;
      end
    end else begin
      reservedValidList3_48 <= _GEN_2480;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_49 <= _GEN_2481;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_49 <= _GEN_2481;
        end else begin
          reservedValidList3_49 <= _GEN_4089;
        end
      end else begin
        reservedValidList3_49 <= _GEN_2481;
      end
    end else begin
      reservedValidList3_49 <= _GEN_2481;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_50 <= _GEN_2482;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_50 <= _GEN_2482;
        end else begin
          reservedValidList3_50 <= _GEN_4090;
        end
      end else begin
        reservedValidList3_50 <= _GEN_2482;
      end
    end else begin
      reservedValidList3_50 <= _GEN_2482;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_51 <= _GEN_2483;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_51 <= _GEN_2483;
        end else begin
          reservedValidList3_51 <= _GEN_4091;
        end
      end else begin
        reservedValidList3_51 <= _GEN_2483;
      end
    end else begin
      reservedValidList3_51 <= _GEN_2483;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_52 <= _GEN_2484;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_52 <= _GEN_2484;
        end else begin
          reservedValidList3_52 <= _GEN_4092;
        end
      end else begin
        reservedValidList3_52 <= _GEN_2484;
      end
    end else begin
      reservedValidList3_52 <= _GEN_2484;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_53 <= _GEN_2485;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_53 <= _GEN_2485;
        end else begin
          reservedValidList3_53 <= _GEN_4093;
        end
      end else begin
        reservedValidList3_53 <= _GEN_2485;
      end
    end else begin
      reservedValidList3_53 <= _GEN_2485;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_54 <= _GEN_2486;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_54 <= _GEN_2486;
        end else begin
          reservedValidList3_54 <= _GEN_4094;
        end
      end else begin
        reservedValidList3_54 <= _GEN_2486;
      end
    end else begin
      reservedValidList3_54 <= _GEN_2486;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_55 <= _GEN_2487;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_55 <= _GEN_2487;
        end else begin
          reservedValidList3_55 <= _GEN_4095;
        end
      end else begin
        reservedValidList3_55 <= _GEN_2487;
      end
    end else begin
      reservedValidList3_55 <= _GEN_2487;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_56 <= _GEN_2488;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_56 <= _GEN_2488;
        end else begin
          reservedValidList3_56 <= _GEN_4096;
        end
      end else begin
        reservedValidList3_56 <= _GEN_2488;
      end
    end else begin
      reservedValidList3_56 <= _GEN_2488;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_57 <= _GEN_2489;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_57 <= _GEN_2489;
        end else begin
          reservedValidList3_57 <= _GEN_4097;
        end
      end else begin
        reservedValidList3_57 <= _GEN_2489;
      end
    end else begin
      reservedValidList3_57 <= _GEN_2489;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_58 <= _GEN_2490;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_58 <= _GEN_2490;
        end else begin
          reservedValidList3_58 <= _GEN_4098;
        end
      end else begin
        reservedValidList3_58 <= _GEN_2490;
      end
    end else begin
      reservedValidList3_58 <= _GEN_2490;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_59 <= _GEN_2491;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_59 <= _GEN_2491;
        end else begin
          reservedValidList3_59 <= _GEN_4099;
        end
      end else begin
        reservedValidList3_59 <= _GEN_2491;
      end
    end else begin
      reservedValidList3_59 <= _GEN_2491;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_60 <= _GEN_2492;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_60 <= _GEN_2492;
        end else begin
          reservedValidList3_60 <= _GEN_4100;
        end
      end else begin
        reservedValidList3_60 <= _GEN_2492;
      end
    end else begin
      reservedValidList3_60 <= _GEN_2492;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_61 <= _GEN_2493;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_61 <= _GEN_2493;
        end else begin
          reservedValidList3_61 <= _GEN_4101;
        end
      end else begin
        reservedValidList3_61 <= _GEN_2493;
      end
    end else begin
      reservedValidList3_61 <= _GEN_2493;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_62 <= _GEN_2494;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_62 <= _GEN_2494;
        end else begin
          reservedValidList3_62 <= _GEN_4102;
        end
      end else begin
        reservedValidList3_62 <= _GEN_2494;
      end
    end else begin
      reservedValidList3_62 <= _GEN_2494;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (3'h0 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_63 <= _GEN_2495;
        end else if (3'h1 == branchTracker) begin // @[decode.scala 400:29]
          reservedValidList3_63 <= _GEN_2495;
        end else begin
          reservedValidList3_63 <= _GEN_4103;
        end
      end else begin
        reservedValidList3_63 <= _GEN_2495;
      end
    end else begin
      reservedValidList3_63 <= _GEN_2495;
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_0 <= _GEN_4200;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_1 <= _GEN_4201;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_2 <= _GEN_4202;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_3 <= _GEN_4203;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_4 <= _GEN_4204;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_5 <= _GEN_4205;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_6 <= _GEN_4206;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_7 <= _GEN_4207;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_8 <= _GEN_4208;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_9 <= _GEN_4209;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_10 <= _GEN_4210;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_11 <= _GEN_4211;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_12 <= _GEN_4212;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_13 <= _GEN_4213;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_14 <= _GEN_4214;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_15 <= _GEN_4215;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_16 <= _GEN_4216;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_17 <= _GEN_4217;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_18 <= _GEN_4218;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_19 <= _GEN_4219;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_20 <= _GEN_4220;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_21 <= _GEN_4221;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_22 <= _GEN_4222;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_23 <= _GEN_4223;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_24 <= _GEN_4224;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_25 <= _GEN_4225;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_26 <= _GEN_4226;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_27 <= _GEN_4227;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_28 <= _GEN_4228;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_29 <= _GEN_4229;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_30 <= _GEN_4230;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_31 <= _GEN_4231;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_32 <= _GEN_4232;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_33 <= _GEN_4233;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_34 <= _GEN_4234;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_35 <= _GEN_4235;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_36 <= _GEN_4236;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_37 <= _GEN_4237;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_38 <= _GEN_4238;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_39 <= _GEN_4239;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_40 <= _GEN_4240;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_41 <= _GEN_4241;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_42 <= _GEN_4242;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_43 <= _GEN_4243;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_44 <= _GEN_4244;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_45 <= _GEN_4245;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_46 <= _GEN_4246;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_47 <= _GEN_4247;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_48 <= _GEN_4248;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_49 <= _GEN_4249;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_50 <= _GEN_4250;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_51 <= _GEN_4251;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_52 <= _GEN_4252;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_53 <= _GEN_4253;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_54 <= _GEN_4254;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_55 <= _GEN_4255;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_56 <= _GEN_4256;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_57 <= _GEN_4257;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_58 <= _GEN_4258;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_59 <= _GEN_4259;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_60 <= _GEN_4260;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_61 <= _GEN_4261;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_62 <= _GEN_4262;
          end
        end
      end
    end
    if (_T_3) begin // @[decode.scala 388:41]
      if (_T_432 | _T_434 | _T_431) begin // @[decode.scala 389:73]
        if (!(3'h0 == branchTracker)) begin // @[decode.scala 400:29]
          if (!(3'h1 == branchTracker)) begin // @[decode.scala 400:29]
            reservedValidList4_63 <= _GEN_4263;
          end
        end
      end
    end
    if (reset) begin // @[decode.scala 464:28]
      ustatus <= 64'h0; // @[decode.scala 464:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (12'h0 == csrAddrReg) begin // @[decode.scala 540:39]
          ustatus <= csrWriteData; // @[decode.scala 541:37]
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        ustatus <= _GEN_7291;
      end else begin
        ustatus <= _GEN_8587;
      end
    end
    if (reset) begin // @[decode.scala 465:28]
      utvec <= 64'h0; // @[decode.scala 465:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 540:39]
          utvec <= _GEN_6968;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        utvec <= _GEN_7292;
      end else begin
        utvec <= _GEN_8588;
      end
    end
    if (reset) begin // @[decode.scala 466:28]
      uepc <= 64'h0; // @[decode.scala 466:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 540:39]
          uepc <= _GEN_6969;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        uepc <= _GEN_7293;
      end else begin
        uepc <= _GEN_8589;
      end
    end
    if (reset) begin // @[decode.scala 467:28]
      ucause <= 64'h0; // @[decode.scala 467:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 540:39]
          ucause <= _GEN_6970;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        ucause <= _GEN_7294;
      end else begin
        ucause <= _GEN_8590;
      end
    end
    if (reset) begin // @[decode.scala 468:28]
      scounteren <= 64'h0; // @[decode.scala 468:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 540:39]
          scounteren <= _GEN_6971;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        scounteren <= _GEN_7295;
      end else begin
        scounteren <= _GEN_8591;
      end
    end
    if (reset) begin // @[decode.scala 469:28]
      satp <= 64'h0; // @[decode.scala 469:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 540:39]
          satp <= _GEN_6972;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        satp <= _GEN_7296;
      end else begin
        satp <= _GEN_8592;
      end
    end
    if (reset) begin // @[decode.scala 470:28]
      mstatus <= 64'h0; // @[decode.scala 470:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] == 3'h0) begin // @[decode.scala 711:126]
      if (writeBackResult_instruction[31:20] == 12'h302) begin // @[decode.scala 712:60]
        mstatus <= _mstatus_T_9; // @[decode.scala 716:15]
      end else if (~(|writeBackResult_instruction[31:20])) begin // @[decode.scala 717:58]
        mstatus <= _mstatus_T_14; // @[decode.scala 724:15]
      end else begin
        mstatus <= _GEN_8691;
      end
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        mstatus <= _GEN_6997;
      end else begin
        mstatus <= _GEN_8617;
      end
    end else begin
      mstatus <= _mstatus_T_1; // @[decode.scala 489:11]
    end
    misa <= _GEN_10392[63:0]; // @[decode.scala 471:{28,28}]
    if (reset) begin // @[decode.scala 472:28]
      medeleg <= 64'h0; // @[decode.scala 472:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 540:39]
          medeleg <= _GEN_6975;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        medeleg <= _GEN_7299;
      end else begin
        medeleg <= _GEN_8595;
      end
    end
    if (reset) begin // @[decode.scala 473:28]
      mideleg <= 64'h0; // @[decode.scala 473:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 540:39]
          mideleg <= _GEN_6976;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        mideleg <= _GEN_7300;
      end else begin
        mideleg <= _GEN_8596;
      end
    end
    if (reset) begin // @[decode.scala 474:28]
      mie <= 64'h0; // @[decode.scala 474:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 540:39]
          mie <= _GEN_6977;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        mie <= _GEN_7301;
      end else begin
        mie <= _GEN_8597;
      end
    end
    if (reset) begin // @[decode.scala 475:28]
      mtvec <= 64'h0; // @[decode.scala 475:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 540:39]
          mtvec <= _GEN_6978;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        mtvec <= _GEN_7302;
      end else begin
        mtvec <= _GEN_8598;
      end
    end
    if (reset) begin // @[decode.scala 476:28]
      mcounteren <= 64'h0; // @[decode.scala 476:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 540:39]
          mcounteren <= _GEN_6979;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        mcounteren <= _GEN_7303;
      end else begin
        mcounteren <= _GEN_8599;
      end
    end
    if (reset) begin // @[decode.scala 477:28]
      mscratch <= 64'h0; // @[decode.scala 477:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 540:39]
          mscratch <= _GEN_6980;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        mscratch <= _GEN_7304;
      end else begin
        mscratch <= _GEN_8600;
      end
    end
    if (reset) begin // @[decode.scala 478:28]
      mepc <= 64'h0; // @[decode.scala 478:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] == 3'h0) begin // @[decode.scala 711:126]
      if (writeBackResult_instruction[31:20] == 12'h302) begin // @[decode.scala 712:60]
        mepc <= _GEN_8674;
      end else if (~(|writeBackResult_instruction[31:20])) begin // @[decode.scala 717:58]
        mepc <= ecallPC; // @[decode.scala 719:12]
      end else begin
        mepc <= _GEN_8687;
      end
    end else begin
      mepc <= _GEN_8674;
    end
    if (reset) begin // @[decode.scala 479:28]
      mcause <= 64'h0; // @[decode.scala 479:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] == 3'h0) begin // @[decode.scala 711:126]
      if (writeBackResult_instruction[31:20] == 12'h302) begin // @[decode.scala 712:60]
        mcause <= _GEN_8675;
      end else if (~(|writeBackResult_instruction[31:20])) begin // @[decode.scala 717:58]
        mcause <= {{60'd0}, _GEN_8686};
      end else begin
        mcause <= _GEN_8688;
      end
    end else begin
      mcause <= _GEN_8675;
    end
    if (reset) begin // @[decode.scala 480:28]
      mtval <= 64'h0; // @[decode.scala 480:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 540:39]
          mtval <= _GEN_6983;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        mtval <= _GEN_7307;
      end else begin
        mtval <= _GEN_8603;
      end
    end
    if (reset) begin // @[decode.scala 481:28]
      mip <= 64'h0; // @[decode.scala 481:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 540:39]
          mip <= _GEN_6984;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        mip <= _GEN_7308;
      end else begin
        mip <= _GEN_8604;
      end
    end
    if (reset) begin // @[decode.scala 482:28]
      pmpcfg0 <= 64'h0; // @[decode.scala 482:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 540:39]
          pmpcfg0 <= _GEN_6985;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        pmpcfg0 <= _GEN_7309;
      end else begin
        pmpcfg0 <= _GEN_8605;
      end
    end
    if (reset) begin // @[decode.scala 483:28]
      pmpaddr0 <= 64'h0; // @[decode.scala 483:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 540:39]
          pmpaddr0 <= _GEN_6986;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        pmpaddr0 <= _GEN_7310;
      end else begin
        pmpaddr0 <= _GEN_8606;
      end
    end
    if (reset) begin // @[decode.scala 484:28]
      mvendorid <= 64'h0; // @[decode.scala 484:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 540:39]
          mvendorid <= _GEN_6987;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        mvendorid <= _GEN_7311;
      end else begin
        mvendorid <= _GEN_8607;
      end
    end
    if (reset) begin // @[decode.scala 485:28]
      marchid <= 64'h0; // @[decode.scala 485:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 540:39]
          marchid <= _GEN_6988;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        marchid <= _GEN_7312;
      end else begin
        marchid <= _GEN_8608;
      end
    end
    if (reset) begin // @[decode.scala 486:28]
      mimpid <= 64'h0; // @[decode.scala 486:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 540:39]
          mimpid <= _GEN_6989;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        mimpid <= _GEN_7313;
      end else begin
        mimpid <= _GEN_8609;
      end
    end
    if (reset) begin // @[decode.scala 487:28]
      mhartid <= 64'h0; // @[decode.scala 487:28]
    end else if (_T_246 & writeBackResult_instruction[14:12] != 3'h0) begin // @[decode.scala 535:126]
      if (3'h1 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        if (!(12'h0 == csrAddrReg)) begin // @[decode.scala 540:39]
          mhartid <= _GEN_6990;
        end
      end else if (3'h2 == writeBackResult_instruction[14:12]) begin // @[decode.scala 538:48]
        mhartid <= _GEN_7314;
      end else begin
        mhartid <= _GEN_8610;
      end
    end
    if (reset) begin // @[decode.scala 710:33]
      currentPrivilege <= 64'h2200000000; // @[decode.scala 710:33]
    end else if (_T_246 & writeBackResult_instruction[14:12] == 3'h0) begin // @[decode.scala 711:126]
      if (writeBackResult_instruction[31:20] == 12'h302) begin // @[decode.scala 712:60]
        currentPrivilege <= {{26'd0}, _GEN_8685}; // @[decode.scala 714:24]
      end else if (~(|writeBackResult_instruction[31:20])) begin // @[decode.scala 717:58]
        currentPrivilege <= 64'h2200000000; // @[decode.scala 722:24]
      end else begin
        currentPrivilege <= _GEN_8689;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  inputBuffer_pc = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  inputBuffer_instruction = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  outputBuffer_instruction = _RAND_2[31:0];
  _RAND_3 = {2{`RANDOM}};
  outputBuffer_pc = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  outputBuffer_PRFDest = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  outputBuffer_rs1Addr = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  outputBuffer_rs2Addr = _RAND_6[5:0];
  _RAND_7 = {2{`RANDOM}};
  outputBuffer_immediate = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  branchBuffer_branchPCReady = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  branchBuffer_predictedPCReady = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  branchBuffer_branchPC = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  branchBuffer_predictedPC = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  branchBuffer_branchMask_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  branchBuffer_branchMask_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  branchBuffer_branchMask_2 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  branchBuffer_branchMask_3 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  branchTracker = _RAND_16[2:0];
  _RAND_17 = {2{`RANDOM}};
  expectedPC = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  stateRegInputBuf = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  stateRegOutputBuf = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  stallReg = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  ecallPC = _RAND_21[63:0];
  _RAND_22 = {1{`RANDOM}};
  PRFValidList_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  PRFValidList_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  PRFValidList_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  PRFValidList_3 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  PRFValidList_4 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  PRFValidList_5 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  PRFValidList_6 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  PRFValidList_7 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  PRFValidList_8 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  PRFValidList_9 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  PRFValidList_10 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  PRFValidList_11 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  PRFValidList_12 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  PRFValidList_13 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  PRFValidList_14 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  PRFValidList_15 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  PRFValidList_16 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  PRFValidList_17 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  PRFValidList_18 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  PRFValidList_19 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  PRFValidList_20 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  PRFValidList_21 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  PRFValidList_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  PRFValidList_23 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  PRFValidList_24 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  PRFValidList_25 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  PRFValidList_26 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  PRFValidList_27 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  PRFValidList_28 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  PRFValidList_29 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  PRFValidList_30 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  PRFValidList_31 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  PRFValidList_32 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  PRFValidList_33 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  PRFValidList_34 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  PRFValidList_35 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  PRFValidList_36 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  PRFValidList_37 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  PRFValidList_38 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  PRFValidList_39 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  PRFValidList_40 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  PRFValidList_41 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  PRFValidList_42 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  PRFValidList_43 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  PRFValidList_44 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  PRFValidList_45 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  PRFValidList_46 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  PRFValidList_47 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  PRFValidList_48 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  PRFValidList_49 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  PRFValidList_50 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  PRFValidList_51 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  PRFValidList_52 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  PRFValidList_53 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  PRFValidList_54 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  PRFValidList_55 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  PRFValidList_56 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  PRFValidList_57 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  PRFValidList_58 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  PRFValidList_59 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  PRFValidList_60 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  PRFValidList_61 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  PRFValidList_62 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  PRFValidList_63 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  frontEndRegMap_31 = _RAND_86[5:0];
  _RAND_87 = {1{`RANDOM}};
  frontEndRegMap_30 = _RAND_87[5:0];
  _RAND_88 = {1{`RANDOM}};
  frontEndRegMap_29 = _RAND_88[5:0];
  _RAND_89 = {1{`RANDOM}};
  frontEndRegMap_28 = _RAND_89[5:0];
  _RAND_90 = {1{`RANDOM}};
  frontEndRegMap_27 = _RAND_90[5:0];
  _RAND_91 = {1{`RANDOM}};
  frontEndRegMap_26 = _RAND_91[5:0];
  _RAND_92 = {1{`RANDOM}};
  frontEndRegMap_25 = _RAND_92[5:0];
  _RAND_93 = {1{`RANDOM}};
  frontEndRegMap_24 = _RAND_93[5:0];
  _RAND_94 = {1{`RANDOM}};
  frontEndRegMap_23 = _RAND_94[5:0];
  _RAND_95 = {1{`RANDOM}};
  frontEndRegMap_22 = _RAND_95[5:0];
  _RAND_96 = {1{`RANDOM}};
  frontEndRegMap_21 = _RAND_96[5:0];
  _RAND_97 = {1{`RANDOM}};
  frontEndRegMap_20 = _RAND_97[5:0];
  _RAND_98 = {1{`RANDOM}};
  frontEndRegMap_19 = _RAND_98[5:0];
  _RAND_99 = {1{`RANDOM}};
  frontEndRegMap_18 = _RAND_99[5:0];
  _RAND_100 = {1{`RANDOM}};
  frontEndRegMap_17 = _RAND_100[5:0];
  _RAND_101 = {1{`RANDOM}};
  frontEndRegMap_16 = _RAND_101[5:0];
  _RAND_102 = {1{`RANDOM}};
  frontEndRegMap_15 = _RAND_102[5:0];
  _RAND_103 = {1{`RANDOM}};
  frontEndRegMap_14 = _RAND_103[5:0];
  _RAND_104 = {1{`RANDOM}};
  frontEndRegMap_13 = _RAND_104[5:0];
  _RAND_105 = {1{`RANDOM}};
  frontEndRegMap_12 = _RAND_105[5:0];
  _RAND_106 = {1{`RANDOM}};
  frontEndRegMap_11 = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  frontEndRegMap_10 = _RAND_107[5:0];
  _RAND_108 = {1{`RANDOM}};
  frontEndRegMap_9 = _RAND_108[5:0];
  _RAND_109 = {1{`RANDOM}};
  frontEndRegMap_8 = _RAND_109[5:0];
  _RAND_110 = {1{`RANDOM}};
  frontEndRegMap_7 = _RAND_110[5:0];
  _RAND_111 = {1{`RANDOM}};
  frontEndRegMap_6 = _RAND_111[5:0];
  _RAND_112 = {1{`RANDOM}};
  frontEndRegMap_5 = _RAND_112[5:0];
  _RAND_113 = {1{`RANDOM}};
  frontEndRegMap_4 = _RAND_113[5:0];
  _RAND_114 = {1{`RANDOM}};
  frontEndRegMap_3 = _RAND_114[5:0];
  _RAND_115 = {1{`RANDOM}};
  frontEndRegMap_2 = _RAND_115[5:0];
  _RAND_116 = {1{`RANDOM}};
  frontEndRegMap_1 = _RAND_116[5:0];
  _RAND_117 = {1{`RANDOM}};
  frontEndRegMap_0 = _RAND_117[5:0];
  _RAND_118 = {1{`RANDOM}};
  PRFFreeList_0 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  PRFFreeList_1 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  PRFFreeList_2 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  PRFFreeList_3 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  PRFFreeList_4 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  PRFFreeList_5 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  PRFFreeList_6 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  PRFFreeList_7 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  PRFFreeList_8 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  PRFFreeList_9 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  PRFFreeList_10 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  PRFFreeList_11 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  PRFFreeList_12 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  PRFFreeList_13 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  PRFFreeList_14 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  PRFFreeList_15 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  PRFFreeList_16 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  PRFFreeList_17 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  PRFFreeList_18 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  PRFFreeList_19 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  PRFFreeList_20 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  PRFFreeList_21 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  PRFFreeList_22 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  PRFFreeList_23 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  PRFFreeList_24 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  PRFFreeList_25 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  PRFFreeList_26 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  PRFFreeList_27 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  PRFFreeList_28 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  PRFFreeList_29 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  PRFFreeList_30 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  PRFFreeList_31 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  PRFFreeList_32 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  PRFFreeList_33 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  PRFFreeList_34 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  PRFFreeList_35 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  PRFFreeList_36 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  PRFFreeList_37 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  PRFFreeList_38 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  PRFFreeList_39 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  PRFFreeList_40 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  PRFFreeList_41 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  PRFFreeList_42 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  PRFFreeList_43 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  PRFFreeList_44 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  PRFFreeList_45 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  PRFFreeList_46 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  PRFFreeList_47 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  PRFFreeList_48 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  PRFFreeList_49 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  PRFFreeList_50 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  PRFFreeList_51 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  PRFFreeList_52 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  PRFFreeList_53 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  PRFFreeList_54 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  PRFFreeList_55 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  PRFFreeList_56 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  PRFFreeList_57 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  PRFFreeList_58 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  PRFFreeList_59 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  PRFFreeList_60 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  PRFFreeList_61 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  PRFFreeList_62 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  branchPCMask = _RAND_181[3:0];
  _RAND_182 = {1{`RANDOM}};
  branchReg = _RAND_182[0:0];
  _RAND_183 = {2{`RANDOM}};
  csrReadDataReg = _RAND_183[63:0];
  _RAND_184 = {1{`RANDOM}};
  csrAddrReg = _RAND_184[11:0];
  _RAND_185 = {2{`RANDOM}};
  csrImmReg = _RAND_185[63:0];
  _RAND_186 = {1{`RANDOM}};
  architecturalRegMap_0 = _RAND_186[5:0];
  _RAND_187 = {1{`RANDOM}};
  architecturalRegMap_1 = _RAND_187[5:0];
  _RAND_188 = {1{`RANDOM}};
  architecturalRegMap_2 = _RAND_188[5:0];
  _RAND_189 = {1{`RANDOM}};
  architecturalRegMap_3 = _RAND_189[5:0];
  _RAND_190 = {1{`RANDOM}};
  architecturalRegMap_4 = _RAND_190[5:0];
  _RAND_191 = {1{`RANDOM}};
  architecturalRegMap_5 = _RAND_191[5:0];
  _RAND_192 = {1{`RANDOM}};
  architecturalRegMap_6 = _RAND_192[5:0];
  _RAND_193 = {1{`RANDOM}};
  architecturalRegMap_7 = _RAND_193[5:0];
  _RAND_194 = {1{`RANDOM}};
  architecturalRegMap_8 = _RAND_194[5:0];
  _RAND_195 = {1{`RANDOM}};
  architecturalRegMap_9 = _RAND_195[5:0];
  _RAND_196 = {1{`RANDOM}};
  architecturalRegMap_10 = _RAND_196[5:0];
  _RAND_197 = {1{`RANDOM}};
  architecturalRegMap_11 = _RAND_197[5:0];
  _RAND_198 = {1{`RANDOM}};
  architecturalRegMap_12 = _RAND_198[5:0];
  _RAND_199 = {1{`RANDOM}};
  architecturalRegMap_13 = _RAND_199[5:0];
  _RAND_200 = {1{`RANDOM}};
  architecturalRegMap_14 = _RAND_200[5:0];
  _RAND_201 = {1{`RANDOM}};
  architecturalRegMap_15 = _RAND_201[5:0];
  _RAND_202 = {1{`RANDOM}};
  architecturalRegMap_16 = _RAND_202[5:0];
  _RAND_203 = {1{`RANDOM}};
  architecturalRegMap_17 = _RAND_203[5:0];
  _RAND_204 = {1{`RANDOM}};
  architecturalRegMap_18 = _RAND_204[5:0];
  _RAND_205 = {1{`RANDOM}};
  architecturalRegMap_19 = _RAND_205[5:0];
  _RAND_206 = {1{`RANDOM}};
  architecturalRegMap_20 = _RAND_206[5:0];
  _RAND_207 = {1{`RANDOM}};
  architecturalRegMap_21 = _RAND_207[5:0];
  _RAND_208 = {1{`RANDOM}};
  architecturalRegMap_22 = _RAND_208[5:0];
  _RAND_209 = {1{`RANDOM}};
  architecturalRegMap_23 = _RAND_209[5:0];
  _RAND_210 = {1{`RANDOM}};
  architecturalRegMap_24 = _RAND_210[5:0];
  _RAND_211 = {1{`RANDOM}};
  architecturalRegMap_25 = _RAND_211[5:0];
  _RAND_212 = {1{`RANDOM}};
  architecturalRegMap_26 = _RAND_212[5:0];
  _RAND_213 = {1{`RANDOM}};
  architecturalRegMap_27 = _RAND_213[5:0];
  _RAND_214 = {1{`RANDOM}};
  architecturalRegMap_28 = _RAND_214[5:0];
  _RAND_215 = {1{`RANDOM}};
  architecturalRegMap_29 = _RAND_215[5:0];
  _RAND_216 = {1{`RANDOM}};
  architecturalRegMap_30 = _RAND_216[5:0];
  _RAND_217 = {1{`RANDOM}};
  architecturalRegMap_31 = _RAND_217[5:0];
  _RAND_218 = {1{`RANDOM}};
  reservedRegMap1_0 = _RAND_218[5:0];
  _RAND_219 = {1{`RANDOM}};
  reservedRegMap1_1 = _RAND_219[5:0];
  _RAND_220 = {1{`RANDOM}};
  reservedRegMap1_2 = _RAND_220[5:0];
  _RAND_221 = {1{`RANDOM}};
  reservedRegMap1_3 = _RAND_221[5:0];
  _RAND_222 = {1{`RANDOM}};
  reservedRegMap1_4 = _RAND_222[5:0];
  _RAND_223 = {1{`RANDOM}};
  reservedRegMap1_5 = _RAND_223[5:0];
  _RAND_224 = {1{`RANDOM}};
  reservedRegMap1_6 = _RAND_224[5:0];
  _RAND_225 = {1{`RANDOM}};
  reservedRegMap1_7 = _RAND_225[5:0];
  _RAND_226 = {1{`RANDOM}};
  reservedRegMap1_8 = _RAND_226[5:0];
  _RAND_227 = {1{`RANDOM}};
  reservedRegMap1_9 = _RAND_227[5:0];
  _RAND_228 = {1{`RANDOM}};
  reservedRegMap1_10 = _RAND_228[5:0];
  _RAND_229 = {1{`RANDOM}};
  reservedRegMap1_11 = _RAND_229[5:0];
  _RAND_230 = {1{`RANDOM}};
  reservedRegMap1_12 = _RAND_230[5:0];
  _RAND_231 = {1{`RANDOM}};
  reservedRegMap1_13 = _RAND_231[5:0];
  _RAND_232 = {1{`RANDOM}};
  reservedRegMap1_14 = _RAND_232[5:0];
  _RAND_233 = {1{`RANDOM}};
  reservedRegMap1_15 = _RAND_233[5:0];
  _RAND_234 = {1{`RANDOM}};
  reservedRegMap1_16 = _RAND_234[5:0];
  _RAND_235 = {1{`RANDOM}};
  reservedRegMap1_17 = _RAND_235[5:0];
  _RAND_236 = {1{`RANDOM}};
  reservedRegMap1_18 = _RAND_236[5:0];
  _RAND_237 = {1{`RANDOM}};
  reservedRegMap1_19 = _RAND_237[5:0];
  _RAND_238 = {1{`RANDOM}};
  reservedRegMap1_20 = _RAND_238[5:0];
  _RAND_239 = {1{`RANDOM}};
  reservedRegMap1_21 = _RAND_239[5:0];
  _RAND_240 = {1{`RANDOM}};
  reservedRegMap1_22 = _RAND_240[5:0];
  _RAND_241 = {1{`RANDOM}};
  reservedRegMap1_23 = _RAND_241[5:0];
  _RAND_242 = {1{`RANDOM}};
  reservedRegMap1_24 = _RAND_242[5:0];
  _RAND_243 = {1{`RANDOM}};
  reservedRegMap1_25 = _RAND_243[5:0];
  _RAND_244 = {1{`RANDOM}};
  reservedRegMap1_26 = _RAND_244[5:0];
  _RAND_245 = {1{`RANDOM}};
  reservedRegMap1_27 = _RAND_245[5:0];
  _RAND_246 = {1{`RANDOM}};
  reservedRegMap1_28 = _RAND_246[5:0];
  _RAND_247 = {1{`RANDOM}};
  reservedRegMap1_29 = _RAND_247[5:0];
  _RAND_248 = {1{`RANDOM}};
  reservedRegMap1_30 = _RAND_248[5:0];
  _RAND_249 = {1{`RANDOM}};
  reservedRegMap1_31 = _RAND_249[5:0];
  _RAND_250 = {1{`RANDOM}};
  reservedRegMap2_0 = _RAND_250[5:0];
  _RAND_251 = {1{`RANDOM}};
  reservedRegMap2_1 = _RAND_251[5:0];
  _RAND_252 = {1{`RANDOM}};
  reservedRegMap2_2 = _RAND_252[5:0];
  _RAND_253 = {1{`RANDOM}};
  reservedRegMap2_3 = _RAND_253[5:0];
  _RAND_254 = {1{`RANDOM}};
  reservedRegMap2_4 = _RAND_254[5:0];
  _RAND_255 = {1{`RANDOM}};
  reservedRegMap2_5 = _RAND_255[5:0];
  _RAND_256 = {1{`RANDOM}};
  reservedRegMap2_6 = _RAND_256[5:0];
  _RAND_257 = {1{`RANDOM}};
  reservedRegMap2_7 = _RAND_257[5:0];
  _RAND_258 = {1{`RANDOM}};
  reservedRegMap2_8 = _RAND_258[5:0];
  _RAND_259 = {1{`RANDOM}};
  reservedRegMap2_9 = _RAND_259[5:0];
  _RAND_260 = {1{`RANDOM}};
  reservedRegMap2_10 = _RAND_260[5:0];
  _RAND_261 = {1{`RANDOM}};
  reservedRegMap2_11 = _RAND_261[5:0];
  _RAND_262 = {1{`RANDOM}};
  reservedRegMap2_12 = _RAND_262[5:0];
  _RAND_263 = {1{`RANDOM}};
  reservedRegMap2_13 = _RAND_263[5:0];
  _RAND_264 = {1{`RANDOM}};
  reservedRegMap2_14 = _RAND_264[5:0];
  _RAND_265 = {1{`RANDOM}};
  reservedRegMap2_15 = _RAND_265[5:0];
  _RAND_266 = {1{`RANDOM}};
  reservedRegMap2_16 = _RAND_266[5:0];
  _RAND_267 = {1{`RANDOM}};
  reservedRegMap2_17 = _RAND_267[5:0];
  _RAND_268 = {1{`RANDOM}};
  reservedRegMap2_18 = _RAND_268[5:0];
  _RAND_269 = {1{`RANDOM}};
  reservedRegMap2_19 = _RAND_269[5:0];
  _RAND_270 = {1{`RANDOM}};
  reservedRegMap2_20 = _RAND_270[5:0];
  _RAND_271 = {1{`RANDOM}};
  reservedRegMap2_21 = _RAND_271[5:0];
  _RAND_272 = {1{`RANDOM}};
  reservedRegMap2_22 = _RAND_272[5:0];
  _RAND_273 = {1{`RANDOM}};
  reservedRegMap2_23 = _RAND_273[5:0];
  _RAND_274 = {1{`RANDOM}};
  reservedRegMap2_24 = _RAND_274[5:0];
  _RAND_275 = {1{`RANDOM}};
  reservedRegMap2_25 = _RAND_275[5:0];
  _RAND_276 = {1{`RANDOM}};
  reservedRegMap2_26 = _RAND_276[5:0];
  _RAND_277 = {1{`RANDOM}};
  reservedRegMap2_27 = _RAND_277[5:0];
  _RAND_278 = {1{`RANDOM}};
  reservedRegMap2_28 = _RAND_278[5:0];
  _RAND_279 = {1{`RANDOM}};
  reservedRegMap2_29 = _RAND_279[5:0];
  _RAND_280 = {1{`RANDOM}};
  reservedRegMap2_30 = _RAND_280[5:0];
  _RAND_281 = {1{`RANDOM}};
  reservedRegMap2_31 = _RAND_281[5:0];
  _RAND_282 = {1{`RANDOM}};
  reservedRegMap3_0 = _RAND_282[5:0];
  _RAND_283 = {1{`RANDOM}};
  reservedRegMap3_1 = _RAND_283[5:0];
  _RAND_284 = {1{`RANDOM}};
  reservedRegMap3_2 = _RAND_284[5:0];
  _RAND_285 = {1{`RANDOM}};
  reservedRegMap3_3 = _RAND_285[5:0];
  _RAND_286 = {1{`RANDOM}};
  reservedRegMap3_4 = _RAND_286[5:0];
  _RAND_287 = {1{`RANDOM}};
  reservedRegMap3_5 = _RAND_287[5:0];
  _RAND_288 = {1{`RANDOM}};
  reservedRegMap3_6 = _RAND_288[5:0];
  _RAND_289 = {1{`RANDOM}};
  reservedRegMap3_7 = _RAND_289[5:0];
  _RAND_290 = {1{`RANDOM}};
  reservedRegMap3_8 = _RAND_290[5:0];
  _RAND_291 = {1{`RANDOM}};
  reservedRegMap3_9 = _RAND_291[5:0];
  _RAND_292 = {1{`RANDOM}};
  reservedRegMap3_10 = _RAND_292[5:0];
  _RAND_293 = {1{`RANDOM}};
  reservedRegMap3_11 = _RAND_293[5:0];
  _RAND_294 = {1{`RANDOM}};
  reservedRegMap3_12 = _RAND_294[5:0];
  _RAND_295 = {1{`RANDOM}};
  reservedRegMap3_13 = _RAND_295[5:0];
  _RAND_296 = {1{`RANDOM}};
  reservedRegMap3_14 = _RAND_296[5:0];
  _RAND_297 = {1{`RANDOM}};
  reservedRegMap3_15 = _RAND_297[5:0];
  _RAND_298 = {1{`RANDOM}};
  reservedRegMap3_16 = _RAND_298[5:0];
  _RAND_299 = {1{`RANDOM}};
  reservedRegMap3_17 = _RAND_299[5:0];
  _RAND_300 = {1{`RANDOM}};
  reservedRegMap3_18 = _RAND_300[5:0];
  _RAND_301 = {1{`RANDOM}};
  reservedRegMap3_19 = _RAND_301[5:0];
  _RAND_302 = {1{`RANDOM}};
  reservedRegMap3_20 = _RAND_302[5:0];
  _RAND_303 = {1{`RANDOM}};
  reservedRegMap3_21 = _RAND_303[5:0];
  _RAND_304 = {1{`RANDOM}};
  reservedRegMap3_22 = _RAND_304[5:0];
  _RAND_305 = {1{`RANDOM}};
  reservedRegMap3_23 = _RAND_305[5:0];
  _RAND_306 = {1{`RANDOM}};
  reservedRegMap3_24 = _RAND_306[5:0];
  _RAND_307 = {1{`RANDOM}};
  reservedRegMap3_25 = _RAND_307[5:0];
  _RAND_308 = {1{`RANDOM}};
  reservedRegMap3_26 = _RAND_308[5:0];
  _RAND_309 = {1{`RANDOM}};
  reservedRegMap3_27 = _RAND_309[5:0];
  _RAND_310 = {1{`RANDOM}};
  reservedRegMap3_28 = _RAND_310[5:0];
  _RAND_311 = {1{`RANDOM}};
  reservedRegMap3_29 = _RAND_311[5:0];
  _RAND_312 = {1{`RANDOM}};
  reservedRegMap3_30 = _RAND_312[5:0];
  _RAND_313 = {1{`RANDOM}};
  reservedRegMap3_31 = _RAND_313[5:0];
  _RAND_314 = {1{`RANDOM}};
  reservedRegMap4_0 = _RAND_314[5:0];
  _RAND_315 = {1{`RANDOM}};
  reservedRegMap4_1 = _RAND_315[5:0];
  _RAND_316 = {1{`RANDOM}};
  reservedRegMap4_2 = _RAND_316[5:0];
  _RAND_317 = {1{`RANDOM}};
  reservedRegMap4_3 = _RAND_317[5:0];
  _RAND_318 = {1{`RANDOM}};
  reservedRegMap4_4 = _RAND_318[5:0];
  _RAND_319 = {1{`RANDOM}};
  reservedRegMap4_5 = _RAND_319[5:0];
  _RAND_320 = {1{`RANDOM}};
  reservedRegMap4_6 = _RAND_320[5:0];
  _RAND_321 = {1{`RANDOM}};
  reservedRegMap4_7 = _RAND_321[5:0];
  _RAND_322 = {1{`RANDOM}};
  reservedRegMap4_8 = _RAND_322[5:0];
  _RAND_323 = {1{`RANDOM}};
  reservedRegMap4_9 = _RAND_323[5:0];
  _RAND_324 = {1{`RANDOM}};
  reservedRegMap4_10 = _RAND_324[5:0];
  _RAND_325 = {1{`RANDOM}};
  reservedRegMap4_11 = _RAND_325[5:0];
  _RAND_326 = {1{`RANDOM}};
  reservedRegMap4_12 = _RAND_326[5:0];
  _RAND_327 = {1{`RANDOM}};
  reservedRegMap4_13 = _RAND_327[5:0];
  _RAND_328 = {1{`RANDOM}};
  reservedRegMap4_14 = _RAND_328[5:0];
  _RAND_329 = {1{`RANDOM}};
  reservedRegMap4_15 = _RAND_329[5:0];
  _RAND_330 = {1{`RANDOM}};
  reservedRegMap4_16 = _RAND_330[5:0];
  _RAND_331 = {1{`RANDOM}};
  reservedRegMap4_17 = _RAND_331[5:0];
  _RAND_332 = {1{`RANDOM}};
  reservedRegMap4_18 = _RAND_332[5:0];
  _RAND_333 = {1{`RANDOM}};
  reservedRegMap4_19 = _RAND_333[5:0];
  _RAND_334 = {1{`RANDOM}};
  reservedRegMap4_20 = _RAND_334[5:0];
  _RAND_335 = {1{`RANDOM}};
  reservedRegMap4_21 = _RAND_335[5:0];
  _RAND_336 = {1{`RANDOM}};
  reservedRegMap4_22 = _RAND_336[5:0];
  _RAND_337 = {1{`RANDOM}};
  reservedRegMap4_23 = _RAND_337[5:0];
  _RAND_338 = {1{`RANDOM}};
  reservedRegMap4_24 = _RAND_338[5:0];
  _RAND_339 = {1{`RANDOM}};
  reservedRegMap4_25 = _RAND_339[5:0];
  _RAND_340 = {1{`RANDOM}};
  reservedRegMap4_26 = _RAND_340[5:0];
  _RAND_341 = {1{`RANDOM}};
  reservedRegMap4_27 = _RAND_341[5:0];
  _RAND_342 = {1{`RANDOM}};
  reservedRegMap4_28 = _RAND_342[5:0];
  _RAND_343 = {1{`RANDOM}};
  reservedRegMap4_29 = _RAND_343[5:0];
  _RAND_344 = {1{`RANDOM}};
  reservedRegMap4_30 = _RAND_344[5:0];
  _RAND_345 = {1{`RANDOM}};
  reservedRegMap4_31 = _RAND_345[5:0];
  _RAND_346 = {1{`RANDOM}};
  reservedFreeList1_0 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  reservedFreeList1_1 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  reservedFreeList1_2 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  reservedFreeList1_3 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  reservedFreeList1_4 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  reservedFreeList1_5 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  reservedFreeList1_6 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  reservedFreeList1_7 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  reservedFreeList1_8 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  reservedFreeList1_9 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  reservedFreeList1_10 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  reservedFreeList1_11 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  reservedFreeList1_12 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  reservedFreeList1_13 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  reservedFreeList1_14 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  reservedFreeList1_15 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  reservedFreeList1_16 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  reservedFreeList1_17 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  reservedFreeList1_18 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  reservedFreeList1_19 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  reservedFreeList1_20 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  reservedFreeList1_21 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  reservedFreeList1_22 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  reservedFreeList1_23 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  reservedFreeList1_24 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  reservedFreeList1_25 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  reservedFreeList1_26 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  reservedFreeList1_27 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  reservedFreeList1_28 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  reservedFreeList1_29 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  reservedFreeList1_30 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  reservedFreeList1_31 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  reservedFreeList1_32 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  reservedFreeList1_33 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  reservedFreeList1_34 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  reservedFreeList1_35 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  reservedFreeList1_36 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  reservedFreeList1_37 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  reservedFreeList1_38 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  reservedFreeList1_39 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  reservedFreeList1_40 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  reservedFreeList1_41 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  reservedFreeList1_42 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  reservedFreeList1_43 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  reservedFreeList1_44 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  reservedFreeList1_45 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  reservedFreeList1_46 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  reservedFreeList1_47 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  reservedFreeList1_48 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  reservedFreeList1_49 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  reservedFreeList1_50 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  reservedFreeList1_51 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  reservedFreeList1_52 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  reservedFreeList1_53 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  reservedFreeList1_54 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  reservedFreeList1_55 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  reservedFreeList1_56 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  reservedFreeList1_57 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  reservedFreeList1_58 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  reservedFreeList1_59 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  reservedFreeList1_60 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  reservedFreeList1_61 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  reservedFreeList1_62 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  reservedFreeList2_0 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  reservedFreeList2_1 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  reservedFreeList2_2 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  reservedFreeList2_3 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  reservedFreeList2_4 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  reservedFreeList2_5 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  reservedFreeList2_6 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  reservedFreeList2_7 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  reservedFreeList2_8 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  reservedFreeList2_9 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  reservedFreeList2_10 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  reservedFreeList2_11 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  reservedFreeList2_12 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  reservedFreeList2_13 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  reservedFreeList2_14 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  reservedFreeList2_15 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  reservedFreeList2_16 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  reservedFreeList2_17 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  reservedFreeList2_18 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  reservedFreeList2_19 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  reservedFreeList2_20 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  reservedFreeList2_21 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  reservedFreeList2_22 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  reservedFreeList2_23 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  reservedFreeList2_24 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  reservedFreeList2_25 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  reservedFreeList2_26 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  reservedFreeList2_27 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  reservedFreeList2_28 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  reservedFreeList2_29 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  reservedFreeList2_30 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  reservedFreeList2_31 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  reservedFreeList2_32 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  reservedFreeList2_33 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  reservedFreeList2_34 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  reservedFreeList2_35 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  reservedFreeList2_36 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  reservedFreeList2_37 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  reservedFreeList2_38 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  reservedFreeList2_39 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  reservedFreeList2_40 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  reservedFreeList2_41 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  reservedFreeList2_42 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  reservedFreeList2_43 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  reservedFreeList2_44 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  reservedFreeList2_45 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  reservedFreeList2_46 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  reservedFreeList2_47 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  reservedFreeList2_48 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  reservedFreeList2_49 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  reservedFreeList2_50 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  reservedFreeList2_51 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  reservedFreeList2_52 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  reservedFreeList2_53 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  reservedFreeList2_54 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  reservedFreeList2_55 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  reservedFreeList2_56 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  reservedFreeList2_57 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  reservedFreeList2_58 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  reservedFreeList2_59 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  reservedFreeList2_60 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  reservedFreeList2_61 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  reservedFreeList2_62 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  reservedFreeList3_0 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  reservedFreeList3_1 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  reservedFreeList3_2 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  reservedFreeList3_3 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  reservedFreeList3_4 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  reservedFreeList3_5 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  reservedFreeList3_6 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  reservedFreeList3_7 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  reservedFreeList3_8 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  reservedFreeList3_9 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  reservedFreeList3_10 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  reservedFreeList3_11 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  reservedFreeList3_12 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  reservedFreeList3_13 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  reservedFreeList3_14 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  reservedFreeList3_15 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  reservedFreeList3_16 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  reservedFreeList3_17 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  reservedFreeList3_18 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  reservedFreeList3_19 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  reservedFreeList3_20 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  reservedFreeList3_21 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  reservedFreeList3_22 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  reservedFreeList3_23 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  reservedFreeList3_24 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  reservedFreeList3_25 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  reservedFreeList3_26 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  reservedFreeList3_27 = _RAND_499[0:0];
  _RAND_500 = {1{`RANDOM}};
  reservedFreeList3_28 = _RAND_500[0:0];
  _RAND_501 = {1{`RANDOM}};
  reservedFreeList3_29 = _RAND_501[0:0];
  _RAND_502 = {1{`RANDOM}};
  reservedFreeList3_30 = _RAND_502[0:0];
  _RAND_503 = {1{`RANDOM}};
  reservedFreeList3_31 = _RAND_503[0:0];
  _RAND_504 = {1{`RANDOM}};
  reservedFreeList3_32 = _RAND_504[0:0];
  _RAND_505 = {1{`RANDOM}};
  reservedFreeList3_33 = _RAND_505[0:0];
  _RAND_506 = {1{`RANDOM}};
  reservedFreeList3_34 = _RAND_506[0:0];
  _RAND_507 = {1{`RANDOM}};
  reservedFreeList3_35 = _RAND_507[0:0];
  _RAND_508 = {1{`RANDOM}};
  reservedFreeList3_36 = _RAND_508[0:0];
  _RAND_509 = {1{`RANDOM}};
  reservedFreeList3_37 = _RAND_509[0:0];
  _RAND_510 = {1{`RANDOM}};
  reservedFreeList3_38 = _RAND_510[0:0];
  _RAND_511 = {1{`RANDOM}};
  reservedFreeList3_39 = _RAND_511[0:0];
  _RAND_512 = {1{`RANDOM}};
  reservedFreeList3_40 = _RAND_512[0:0];
  _RAND_513 = {1{`RANDOM}};
  reservedFreeList3_41 = _RAND_513[0:0];
  _RAND_514 = {1{`RANDOM}};
  reservedFreeList3_42 = _RAND_514[0:0];
  _RAND_515 = {1{`RANDOM}};
  reservedFreeList3_43 = _RAND_515[0:0];
  _RAND_516 = {1{`RANDOM}};
  reservedFreeList3_44 = _RAND_516[0:0];
  _RAND_517 = {1{`RANDOM}};
  reservedFreeList3_45 = _RAND_517[0:0];
  _RAND_518 = {1{`RANDOM}};
  reservedFreeList3_46 = _RAND_518[0:0];
  _RAND_519 = {1{`RANDOM}};
  reservedFreeList3_47 = _RAND_519[0:0];
  _RAND_520 = {1{`RANDOM}};
  reservedFreeList3_48 = _RAND_520[0:0];
  _RAND_521 = {1{`RANDOM}};
  reservedFreeList3_49 = _RAND_521[0:0];
  _RAND_522 = {1{`RANDOM}};
  reservedFreeList3_50 = _RAND_522[0:0];
  _RAND_523 = {1{`RANDOM}};
  reservedFreeList3_51 = _RAND_523[0:0];
  _RAND_524 = {1{`RANDOM}};
  reservedFreeList3_52 = _RAND_524[0:0];
  _RAND_525 = {1{`RANDOM}};
  reservedFreeList3_53 = _RAND_525[0:0];
  _RAND_526 = {1{`RANDOM}};
  reservedFreeList3_54 = _RAND_526[0:0];
  _RAND_527 = {1{`RANDOM}};
  reservedFreeList3_55 = _RAND_527[0:0];
  _RAND_528 = {1{`RANDOM}};
  reservedFreeList3_56 = _RAND_528[0:0];
  _RAND_529 = {1{`RANDOM}};
  reservedFreeList3_57 = _RAND_529[0:0];
  _RAND_530 = {1{`RANDOM}};
  reservedFreeList3_58 = _RAND_530[0:0];
  _RAND_531 = {1{`RANDOM}};
  reservedFreeList3_59 = _RAND_531[0:0];
  _RAND_532 = {1{`RANDOM}};
  reservedFreeList3_60 = _RAND_532[0:0];
  _RAND_533 = {1{`RANDOM}};
  reservedFreeList3_61 = _RAND_533[0:0];
  _RAND_534 = {1{`RANDOM}};
  reservedFreeList3_62 = _RAND_534[0:0];
  _RAND_535 = {1{`RANDOM}};
  reservedFreeList4_0 = _RAND_535[0:0];
  _RAND_536 = {1{`RANDOM}};
  reservedFreeList4_1 = _RAND_536[0:0];
  _RAND_537 = {1{`RANDOM}};
  reservedFreeList4_2 = _RAND_537[0:0];
  _RAND_538 = {1{`RANDOM}};
  reservedFreeList4_3 = _RAND_538[0:0];
  _RAND_539 = {1{`RANDOM}};
  reservedFreeList4_4 = _RAND_539[0:0];
  _RAND_540 = {1{`RANDOM}};
  reservedFreeList4_5 = _RAND_540[0:0];
  _RAND_541 = {1{`RANDOM}};
  reservedFreeList4_6 = _RAND_541[0:0];
  _RAND_542 = {1{`RANDOM}};
  reservedFreeList4_7 = _RAND_542[0:0];
  _RAND_543 = {1{`RANDOM}};
  reservedFreeList4_8 = _RAND_543[0:0];
  _RAND_544 = {1{`RANDOM}};
  reservedFreeList4_9 = _RAND_544[0:0];
  _RAND_545 = {1{`RANDOM}};
  reservedFreeList4_10 = _RAND_545[0:0];
  _RAND_546 = {1{`RANDOM}};
  reservedFreeList4_11 = _RAND_546[0:0];
  _RAND_547 = {1{`RANDOM}};
  reservedFreeList4_12 = _RAND_547[0:0];
  _RAND_548 = {1{`RANDOM}};
  reservedFreeList4_13 = _RAND_548[0:0];
  _RAND_549 = {1{`RANDOM}};
  reservedFreeList4_14 = _RAND_549[0:0];
  _RAND_550 = {1{`RANDOM}};
  reservedFreeList4_15 = _RAND_550[0:0];
  _RAND_551 = {1{`RANDOM}};
  reservedFreeList4_16 = _RAND_551[0:0];
  _RAND_552 = {1{`RANDOM}};
  reservedFreeList4_17 = _RAND_552[0:0];
  _RAND_553 = {1{`RANDOM}};
  reservedFreeList4_18 = _RAND_553[0:0];
  _RAND_554 = {1{`RANDOM}};
  reservedFreeList4_19 = _RAND_554[0:0];
  _RAND_555 = {1{`RANDOM}};
  reservedFreeList4_20 = _RAND_555[0:0];
  _RAND_556 = {1{`RANDOM}};
  reservedFreeList4_21 = _RAND_556[0:0];
  _RAND_557 = {1{`RANDOM}};
  reservedFreeList4_22 = _RAND_557[0:0];
  _RAND_558 = {1{`RANDOM}};
  reservedFreeList4_23 = _RAND_558[0:0];
  _RAND_559 = {1{`RANDOM}};
  reservedFreeList4_24 = _RAND_559[0:0];
  _RAND_560 = {1{`RANDOM}};
  reservedFreeList4_25 = _RAND_560[0:0];
  _RAND_561 = {1{`RANDOM}};
  reservedFreeList4_26 = _RAND_561[0:0];
  _RAND_562 = {1{`RANDOM}};
  reservedFreeList4_27 = _RAND_562[0:0];
  _RAND_563 = {1{`RANDOM}};
  reservedFreeList4_28 = _RAND_563[0:0];
  _RAND_564 = {1{`RANDOM}};
  reservedFreeList4_29 = _RAND_564[0:0];
  _RAND_565 = {1{`RANDOM}};
  reservedFreeList4_30 = _RAND_565[0:0];
  _RAND_566 = {1{`RANDOM}};
  reservedFreeList4_31 = _RAND_566[0:0];
  _RAND_567 = {1{`RANDOM}};
  reservedFreeList4_32 = _RAND_567[0:0];
  _RAND_568 = {1{`RANDOM}};
  reservedFreeList4_33 = _RAND_568[0:0];
  _RAND_569 = {1{`RANDOM}};
  reservedFreeList4_34 = _RAND_569[0:0];
  _RAND_570 = {1{`RANDOM}};
  reservedFreeList4_35 = _RAND_570[0:0];
  _RAND_571 = {1{`RANDOM}};
  reservedFreeList4_36 = _RAND_571[0:0];
  _RAND_572 = {1{`RANDOM}};
  reservedFreeList4_37 = _RAND_572[0:0];
  _RAND_573 = {1{`RANDOM}};
  reservedFreeList4_38 = _RAND_573[0:0];
  _RAND_574 = {1{`RANDOM}};
  reservedFreeList4_39 = _RAND_574[0:0];
  _RAND_575 = {1{`RANDOM}};
  reservedFreeList4_40 = _RAND_575[0:0];
  _RAND_576 = {1{`RANDOM}};
  reservedFreeList4_41 = _RAND_576[0:0];
  _RAND_577 = {1{`RANDOM}};
  reservedFreeList4_42 = _RAND_577[0:0];
  _RAND_578 = {1{`RANDOM}};
  reservedFreeList4_43 = _RAND_578[0:0];
  _RAND_579 = {1{`RANDOM}};
  reservedFreeList4_44 = _RAND_579[0:0];
  _RAND_580 = {1{`RANDOM}};
  reservedFreeList4_45 = _RAND_580[0:0];
  _RAND_581 = {1{`RANDOM}};
  reservedFreeList4_46 = _RAND_581[0:0];
  _RAND_582 = {1{`RANDOM}};
  reservedFreeList4_47 = _RAND_582[0:0];
  _RAND_583 = {1{`RANDOM}};
  reservedFreeList4_48 = _RAND_583[0:0];
  _RAND_584 = {1{`RANDOM}};
  reservedFreeList4_49 = _RAND_584[0:0];
  _RAND_585 = {1{`RANDOM}};
  reservedFreeList4_50 = _RAND_585[0:0];
  _RAND_586 = {1{`RANDOM}};
  reservedFreeList4_51 = _RAND_586[0:0];
  _RAND_587 = {1{`RANDOM}};
  reservedFreeList4_52 = _RAND_587[0:0];
  _RAND_588 = {1{`RANDOM}};
  reservedFreeList4_53 = _RAND_588[0:0];
  _RAND_589 = {1{`RANDOM}};
  reservedFreeList4_54 = _RAND_589[0:0];
  _RAND_590 = {1{`RANDOM}};
  reservedFreeList4_55 = _RAND_590[0:0];
  _RAND_591 = {1{`RANDOM}};
  reservedFreeList4_56 = _RAND_591[0:0];
  _RAND_592 = {1{`RANDOM}};
  reservedFreeList4_57 = _RAND_592[0:0];
  _RAND_593 = {1{`RANDOM}};
  reservedFreeList4_58 = _RAND_593[0:0];
  _RAND_594 = {1{`RANDOM}};
  reservedFreeList4_59 = _RAND_594[0:0];
  _RAND_595 = {1{`RANDOM}};
  reservedFreeList4_60 = _RAND_595[0:0];
  _RAND_596 = {1{`RANDOM}};
  reservedFreeList4_61 = _RAND_596[0:0];
  _RAND_597 = {1{`RANDOM}};
  reservedFreeList4_62 = _RAND_597[0:0];
  _RAND_598 = {1{`RANDOM}};
  reservedValidList1_0 = _RAND_598[0:0];
  _RAND_599 = {1{`RANDOM}};
  reservedValidList1_1 = _RAND_599[0:0];
  _RAND_600 = {1{`RANDOM}};
  reservedValidList1_2 = _RAND_600[0:0];
  _RAND_601 = {1{`RANDOM}};
  reservedValidList1_3 = _RAND_601[0:0];
  _RAND_602 = {1{`RANDOM}};
  reservedValidList1_4 = _RAND_602[0:0];
  _RAND_603 = {1{`RANDOM}};
  reservedValidList1_5 = _RAND_603[0:0];
  _RAND_604 = {1{`RANDOM}};
  reservedValidList1_6 = _RAND_604[0:0];
  _RAND_605 = {1{`RANDOM}};
  reservedValidList1_7 = _RAND_605[0:0];
  _RAND_606 = {1{`RANDOM}};
  reservedValidList1_8 = _RAND_606[0:0];
  _RAND_607 = {1{`RANDOM}};
  reservedValidList1_9 = _RAND_607[0:0];
  _RAND_608 = {1{`RANDOM}};
  reservedValidList1_10 = _RAND_608[0:0];
  _RAND_609 = {1{`RANDOM}};
  reservedValidList1_11 = _RAND_609[0:0];
  _RAND_610 = {1{`RANDOM}};
  reservedValidList1_12 = _RAND_610[0:0];
  _RAND_611 = {1{`RANDOM}};
  reservedValidList1_13 = _RAND_611[0:0];
  _RAND_612 = {1{`RANDOM}};
  reservedValidList1_14 = _RAND_612[0:0];
  _RAND_613 = {1{`RANDOM}};
  reservedValidList1_15 = _RAND_613[0:0];
  _RAND_614 = {1{`RANDOM}};
  reservedValidList1_16 = _RAND_614[0:0];
  _RAND_615 = {1{`RANDOM}};
  reservedValidList1_17 = _RAND_615[0:0];
  _RAND_616 = {1{`RANDOM}};
  reservedValidList1_18 = _RAND_616[0:0];
  _RAND_617 = {1{`RANDOM}};
  reservedValidList1_19 = _RAND_617[0:0];
  _RAND_618 = {1{`RANDOM}};
  reservedValidList1_20 = _RAND_618[0:0];
  _RAND_619 = {1{`RANDOM}};
  reservedValidList1_21 = _RAND_619[0:0];
  _RAND_620 = {1{`RANDOM}};
  reservedValidList1_22 = _RAND_620[0:0];
  _RAND_621 = {1{`RANDOM}};
  reservedValidList1_23 = _RAND_621[0:0];
  _RAND_622 = {1{`RANDOM}};
  reservedValidList1_24 = _RAND_622[0:0];
  _RAND_623 = {1{`RANDOM}};
  reservedValidList1_25 = _RAND_623[0:0];
  _RAND_624 = {1{`RANDOM}};
  reservedValidList1_26 = _RAND_624[0:0];
  _RAND_625 = {1{`RANDOM}};
  reservedValidList1_27 = _RAND_625[0:0];
  _RAND_626 = {1{`RANDOM}};
  reservedValidList1_28 = _RAND_626[0:0];
  _RAND_627 = {1{`RANDOM}};
  reservedValidList1_29 = _RAND_627[0:0];
  _RAND_628 = {1{`RANDOM}};
  reservedValidList1_30 = _RAND_628[0:0];
  _RAND_629 = {1{`RANDOM}};
  reservedValidList1_31 = _RAND_629[0:0];
  _RAND_630 = {1{`RANDOM}};
  reservedValidList1_32 = _RAND_630[0:0];
  _RAND_631 = {1{`RANDOM}};
  reservedValidList1_33 = _RAND_631[0:0];
  _RAND_632 = {1{`RANDOM}};
  reservedValidList1_34 = _RAND_632[0:0];
  _RAND_633 = {1{`RANDOM}};
  reservedValidList1_35 = _RAND_633[0:0];
  _RAND_634 = {1{`RANDOM}};
  reservedValidList1_36 = _RAND_634[0:0];
  _RAND_635 = {1{`RANDOM}};
  reservedValidList1_37 = _RAND_635[0:0];
  _RAND_636 = {1{`RANDOM}};
  reservedValidList1_38 = _RAND_636[0:0];
  _RAND_637 = {1{`RANDOM}};
  reservedValidList1_39 = _RAND_637[0:0];
  _RAND_638 = {1{`RANDOM}};
  reservedValidList1_40 = _RAND_638[0:0];
  _RAND_639 = {1{`RANDOM}};
  reservedValidList1_41 = _RAND_639[0:0];
  _RAND_640 = {1{`RANDOM}};
  reservedValidList1_42 = _RAND_640[0:0];
  _RAND_641 = {1{`RANDOM}};
  reservedValidList1_43 = _RAND_641[0:0];
  _RAND_642 = {1{`RANDOM}};
  reservedValidList1_44 = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  reservedValidList1_45 = _RAND_643[0:0];
  _RAND_644 = {1{`RANDOM}};
  reservedValidList1_46 = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  reservedValidList1_47 = _RAND_645[0:0];
  _RAND_646 = {1{`RANDOM}};
  reservedValidList1_48 = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  reservedValidList1_49 = _RAND_647[0:0];
  _RAND_648 = {1{`RANDOM}};
  reservedValidList1_50 = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  reservedValidList1_51 = _RAND_649[0:0];
  _RAND_650 = {1{`RANDOM}};
  reservedValidList1_52 = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  reservedValidList1_53 = _RAND_651[0:0];
  _RAND_652 = {1{`RANDOM}};
  reservedValidList1_54 = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  reservedValidList1_55 = _RAND_653[0:0];
  _RAND_654 = {1{`RANDOM}};
  reservedValidList1_56 = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  reservedValidList1_57 = _RAND_655[0:0];
  _RAND_656 = {1{`RANDOM}};
  reservedValidList1_58 = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  reservedValidList1_59 = _RAND_657[0:0];
  _RAND_658 = {1{`RANDOM}};
  reservedValidList1_60 = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  reservedValidList1_61 = _RAND_659[0:0];
  _RAND_660 = {1{`RANDOM}};
  reservedValidList1_62 = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  reservedValidList1_63 = _RAND_661[0:0];
  _RAND_662 = {1{`RANDOM}};
  reservedValidList2_0 = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  reservedValidList2_1 = _RAND_663[0:0];
  _RAND_664 = {1{`RANDOM}};
  reservedValidList2_2 = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  reservedValidList2_3 = _RAND_665[0:0];
  _RAND_666 = {1{`RANDOM}};
  reservedValidList2_4 = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  reservedValidList2_5 = _RAND_667[0:0];
  _RAND_668 = {1{`RANDOM}};
  reservedValidList2_6 = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  reservedValidList2_7 = _RAND_669[0:0];
  _RAND_670 = {1{`RANDOM}};
  reservedValidList2_8 = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  reservedValidList2_9 = _RAND_671[0:0];
  _RAND_672 = {1{`RANDOM}};
  reservedValidList2_10 = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  reservedValidList2_11 = _RAND_673[0:0];
  _RAND_674 = {1{`RANDOM}};
  reservedValidList2_12 = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  reservedValidList2_13 = _RAND_675[0:0];
  _RAND_676 = {1{`RANDOM}};
  reservedValidList2_14 = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  reservedValidList2_15 = _RAND_677[0:0];
  _RAND_678 = {1{`RANDOM}};
  reservedValidList2_16 = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  reservedValidList2_17 = _RAND_679[0:0];
  _RAND_680 = {1{`RANDOM}};
  reservedValidList2_18 = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  reservedValidList2_19 = _RAND_681[0:0];
  _RAND_682 = {1{`RANDOM}};
  reservedValidList2_20 = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  reservedValidList2_21 = _RAND_683[0:0];
  _RAND_684 = {1{`RANDOM}};
  reservedValidList2_22 = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  reservedValidList2_23 = _RAND_685[0:0];
  _RAND_686 = {1{`RANDOM}};
  reservedValidList2_24 = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  reservedValidList2_25 = _RAND_687[0:0];
  _RAND_688 = {1{`RANDOM}};
  reservedValidList2_26 = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  reservedValidList2_27 = _RAND_689[0:0];
  _RAND_690 = {1{`RANDOM}};
  reservedValidList2_28 = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  reservedValidList2_29 = _RAND_691[0:0];
  _RAND_692 = {1{`RANDOM}};
  reservedValidList2_30 = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  reservedValidList2_31 = _RAND_693[0:0];
  _RAND_694 = {1{`RANDOM}};
  reservedValidList2_32 = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  reservedValidList2_33 = _RAND_695[0:0];
  _RAND_696 = {1{`RANDOM}};
  reservedValidList2_34 = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  reservedValidList2_35 = _RAND_697[0:0];
  _RAND_698 = {1{`RANDOM}};
  reservedValidList2_36 = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  reservedValidList2_37 = _RAND_699[0:0];
  _RAND_700 = {1{`RANDOM}};
  reservedValidList2_38 = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  reservedValidList2_39 = _RAND_701[0:0];
  _RAND_702 = {1{`RANDOM}};
  reservedValidList2_40 = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  reservedValidList2_41 = _RAND_703[0:0];
  _RAND_704 = {1{`RANDOM}};
  reservedValidList2_42 = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  reservedValidList2_43 = _RAND_705[0:0];
  _RAND_706 = {1{`RANDOM}};
  reservedValidList2_44 = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  reservedValidList2_45 = _RAND_707[0:0];
  _RAND_708 = {1{`RANDOM}};
  reservedValidList2_46 = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  reservedValidList2_47 = _RAND_709[0:0];
  _RAND_710 = {1{`RANDOM}};
  reservedValidList2_48 = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  reservedValidList2_49 = _RAND_711[0:0];
  _RAND_712 = {1{`RANDOM}};
  reservedValidList2_50 = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  reservedValidList2_51 = _RAND_713[0:0];
  _RAND_714 = {1{`RANDOM}};
  reservedValidList2_52 = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  reservedValidList2_53 = _RAND_715[0:0];
  _RAND_716 = {1{`RANDOM}};
  reservedValidList2_54 = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  reservedValidList2_55 = _RAND_717[0:0];
  _RAND_718 = {1{`RANDOM}};
  reservedValidList2_56 = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  reservedValidList2_57 = _RAND_719[0:0];
  _RAND_720 = {1{`RANDOM}};
  reservedValidList2_58 = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  reservedValidList2_59 = _RAND_721[0:0];
  _RAND_722 = {1{`RANDOM}};
  reservedValidList2_60 = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  reservedValidList2_61 = _RAND_723[0:0];
  _RAND_724 = {1{`RANDOM}};
  reservedValidList2_62 = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  reservedValidList2_63 = _RAND_725[0:0];
  _RAND_726 = {1{`RANDOM}};
  reservedValidList3_0 = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  reservedValidList3_1 = _RAND_727[0:0];
  _RAND_728 = {1{`RANDOM}};
  reservedValidList3_2 = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  reservedValidList3_3 = _RAND_729[0:0];
  _RAND_730 = {1{`RANDOM}};
  reservedValidList3_4 = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  reservedValidList3_5 = _RAND_731[0:0];
  _RAND_732 = {1{`RANDOM}};
  reservedValidList3_6 = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  reservedValidList3_7 = _RAND_733[0:0];
  _RAND_734 = {1{`RANDOM}};
  reservedValidList3_8 = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  reservedValidList3_9 = _RAND_735[0:0];
  _RAND_736 = {1{`RANDOM}};
  reservedValidList3_10 = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  reservedValidList3_11 = _RAND_737[0:0];
  _RAND_738 = {1{`RANDOM}};
  reservedValidList3_12 = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  reservedValidList3_13 = _RAND_739[0:0];
  _RAND_740 = {1{`RANDOM}};
  reservedValidList3_14 = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  reservedValidList3_15 = _RAND_741[0:0];
  _RAND_742 = {1{`RANDOM}};
  reservedValidList3_16 = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  reservedValidList3_17 = _RAND_743[0:0];
  _RAND_744 = {1{`RANDOM}};
  reservedValidList3_18 = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  reservedValidList3_19 = _RAND_745[0:0];
  _RAND_746 = {1{`RANDOM}};
  reservedValidList3_20 = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  reservedValidList3_21 = _RAND_747[0:0];
  _RAND_748 = {1{`RANDOM}};
  reservedValidList3_22 = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  reservedValidList3_23 = _RAND_749[0:0];
  _RAND_750 = {1{`RANDOM}};
  reservedValidList3_24 = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  reservedValidList3_25 = _RAND_751[0:0];
  _RAND_752 = {1{`RANDOM}};
  reservedValidList3_26 = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  reservedValidList3_27 = _RAND_753[0:0];
  _RAND_754 = {1{`RANDOM}};
  reservedValidList3_28 = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  reservedValidList3_29 = _RAND_755[0:0];
  _RAND_756 = {1{`RANDOM}};
  reservedValidList3_30 = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  reservedValidList3_31 = _RAND_757[0:0];
  _RAND_758 = {1{`RANDOM}};
  reservedValidList3_32 = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  reservedValidList3_33 = _RAND_759[0:0];
  _RAND_760 = {1{`RANDOM}};
  reservedValidList3_34 = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  reservedValidList3_35 = _RAND_761[0:0];
  _RAND_762 = {1{`RANDOM}};
  reservedValidList3_36 = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  reservedValidList3_37 = _RAND_763[0:0];
  _RAND_764 = {1{`RANDOM}};
  reservedValidList3_38 = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  reservedValidList3_39 = _RAND_765[0:0];
  _RAND_766 = {1{`RANDOM}};
  reservedValidList3_40 = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  reservedValidList3_41 = _RAND_767[0:0];
  _RAND_768 = {1{`RANDOM}};
  reservedValidList3_42 = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  reservedValidList3_43 = _RAND_769[0:0];
  _RAND_770 = {1{`RANDOM}};
  reservedValidList3_44 = _RAND_770[0:0];
  _RAND_771 = {1{`RANDOM}};
  reservedValidList3_45 = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  reservedValidList3_46 = _RAND_772[0:0];
  _RAND_773 = {1{`RANDOM}};
  reservedValidList3_47 = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  reservedValidList3_48 = _RAND_774[0:0];
  _RAND_775 = {1{`RANDOM}};
  reservedValidList3_49 = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  reservedValidList3_50 = _RAND_776[0:0];
  _RAND_777 = {1{`RANDOM}};
  reservedValidList3_51 = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  reservedValidList3_52 = _RAND_778[0:0];
  _RAND_779 = {1{`RANDOM}};
  reservedValidList3_53 = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  reservedValidList3_54 = _RAND_780[0:0];
  _RAND_781 = {1{`RANDOM}};
  reservedValidList3_55 = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  reservedValidList3_56 = _RAND_782[0:0];
  _RAND_783 = {1{`RANDOM}};
  reservedValidList3_57 = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  reservedValidList3_58 = _RAND_784[0:0];
  _RAND_785 = {1{`RANDOM}};
  reservedValidList3_59 = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  reservedValidList3_60 = _RAND_786[0:0];
  _RAND_787 = {1{`RANDOM}};
  reservedValidList3_61 = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  reservedValidList3_62 = _RAND_788[0:0];
  _RAND_789 = {1{`RANDOM}};
  reservedValidList3_63 = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  reservedValidList4_0 = _RAND_790[0:0];
  _RAND_791 = {1{`RANDOM}};
  reservedValidList4_1 = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  reservedValidList4_2 = _RAND_792[0:0];
  _RAND_793 = {1{`RANDOM}};
  reservedValidList4_3 = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  reservedValidList4_4 = _RAND_794[0:0];
  _RAND_795 = {1{`RANDOM}};
  reservedValidList4_5 = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  reservedValidList4_6 = _RAND_796[0:0];
  _RAND_797 = {1{`RANDOM}};
  reservedValidList4_7 = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  reservedValidList4_8 = _RAND_798[0:0];
  _RAND_799 = {1{`RANDOM}};
  reservedValidList4_9 = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  reservedValidList4_10 = _RAND_800[0:0];
  _RAND_801 = {1{`RANDOM}};
  reservedValidList4_11 = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  reservedValidList4_12 = _RAND_802[0:0];
  _RAND_803 = {1{`RANDOM}};
  reservedValidList4_13 = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  reservedValidList4_14 = _RAND_804[0:0];
  _RAND_805 = {1{`RANDOM}};
  reservedValidList4_15 = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  reservedValidList4_16 = _RAND_806[0:0];
  _RAND_807 = {1{`RANDOM}};
  reservedValidList4_17 = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  reservedValidList4_18 = _RAND_808[0:0];
  _RAND_809 = {1{`RANDOM}};
  reservedValidList4_19 = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  reservedValidList4_20 = _RAND_810[0:0];
  _RAND_811 = {1{`RANDOM}};
  reservedValidList4_21 = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  reservedValidList4_22 = _RAND_812[0:0];
  _RAND_813 = {1{`RANDOM}};
  reservedValidList4_23 = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  reservedValidList4_24 = _RAND_814[0:0];
  _RAND_815 = {1{`RANDOM}};
  reservedValidList4_25 = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  reservedValidList4_26 = _RAND_816[0:0];
  _RAND_817 = {1{`RANDOM}};
  reservedValidList4_27 = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  reservedValidList4_28 = _RAND_818[0:0];
  _RAND_819 = {1{`RANDOM}};
  reservedValidList4_29 = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  reservedValidList4_30 = _RAND_820[0:0];
  _RAND_821 = {1{`RANDOM}};
  reservedValidList4_31 = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  reservedValidList4_32 = _RAND_822[0:0];
  _RAND_823 = {1{`RANDOM}};
  reservedValidList4_33 = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  reservedValidList4_34 = _RAND_824[0:0];
  _RAND_825 = {1{`RANDOM}};
  reservedValidList4_35 = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  reservedValidList4_36 = _RAND_826[0:0];
  _RAND_827 = {1{`RANDOM}};
  reservedValidList4_37 = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  reservedValidList4_38 = _RAND_828[0:0];
  _RAND_829 = {1{`RANDOM}};
  reservedValidList4_39 = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  reservedValidList4_40 = _RAND_830[0:0];
  _RAND_831 = {1{`RANDOM}};
  reservedValidList4_41 = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  reservedValidList4_42 = _RAND_832[0:0];
  _RAND_833 = {1{`RANDOM}};
  reservedValidList4_43 = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  reservedValidList4_44 = _RAND_834[0:0];
  _RAND_835 = {1{`RANDOM}};
  reservedValidList4_45 = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  reservedValidList4_46 = _RAND_836[0:0];
  _RAND_837 = {1{`RANDOM}};
  reservedValidList4_47 = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  reservedValidList4_48 = _RAND_838[0:0];
  _RAND_839 = {1{`RANDOM}};
  reservedValidList4_49 = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  reservedValidList4_50 = _RAND_840[0:0];
  _RAND_841 = {1{`RANDOM}};
  reservedValidList4_51 = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  reservedValidList4_52 = _RAND_842[0:0];
  _RAND_843 = {1{`RANDOM}};
  reservedValidList4_53 = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  reservedValidList4_54 = _RAND_844[0:0];
  _RAND_845 = {1{`RANDOM}};
  reservedValidList4_55 = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  reservedValidList4_56 = _RAND_846[0:0];
  _RAND_847 = {1{`RANDOM}};
  reservedValidList4_57 = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  reservedValidList4_58 = _RAND_848[0:0];
  _RAND_849 = {1{`RANDOM}};
  reservedValidList4_59 = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  reservedValidList4_60 = _RAND_850[0:0];
  _RAND_851 = {1{`RANDOM}};
  reservedValidList4_61 = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  reservedValidList4_62 = _RAND_852[0:0];
  _RAND_853 = {1{`RANDOM}};
  reservedValidList4_63 = _RAND_853[0:0];
  _RAND_854 = {2{`RANDOM}};
  ustatus = _RAND_854[63:0];
  _RAND_855 = {2{`RANDOM}};
  utvec = _RAND_855[63:0];
  _RAND_856 = {2{`RANDOM}};
  uepc = _RAND_856[63:0];
  _RAND_857 = {2{`RANDOM}};
  ucause = _RAND_857[63:0];
  _RAND_858 = {2{`RANDOM}};
  scounteren = _RAND_858[63:0];
  _RAND_859 = {2{`RANDOM}};
  satp = _RAND_859[63:0];
  _RAND_860 = {2{`RANDOM}};
  mstatus = _RAND_860[63:0];
  _RAND_861 = {2{`RANDOM}};
  misa = _RAND_861[63:0];
  _RAND_862 = {2{`RANDOM}};
  medeleg = _RAND_862[63:0];
  _RAND_863 = {2{`RANDOM}};
  mideleg = _RAND_863[63:0];
  _RAND_864 = {2{`RANDOM}};
  mie = _RAND_864[63:0];
  _RAND_865 = {2{`RANDOM}};
  mtvec = _RAND_865[63:0];
  _RAND_866 = {2{`RANDOM}};
  mcounteren = _RAND_866[63:0];
  _RAND_867 = {2{`RANDOM}};
  mscratch = _RAND_867[63:0];
  _RAND_868 = {2{`RANDOM}};
  mepc = _RAND_868[63:0];
  _RAND_869 = {2{`RANDOM}};
  mcause = _RAND_869[63:0];
  _RAND_870 = {2{`RANDOM}};
  mtval = _RAND_870[63:0];
  _RAND_871 = {2{`RANDOM}};
  mip = _RAND_871[63:0];
  _RAND_872 = {2{`RANDOM}};
  pmpcfg0 = _RAND_872[63:0];
  _RAND_873 = {2{`RANDOM}};
  pmpaddr0 = _RAND_873[63:0];
  _RAND_874 = {2{`RANDOM}};
  mvendorid = _RAND_874[63:0];
  _RAND_875 = {2{`RANDOM}};
  marchid = _RAND_875[63:0];
  _RAND_876 = {2{`RANDOM}};
  mimpid = _RAND_876[63:0];
  _RAND_877 = {2{`RANDOM}};
  mhartid = _RAND_877[63:0];
  _RAND_878 = {2{`RANDOM}};
  currentPrivilege = _RAND_878[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module storeDataIssue_Anon(
  input        clock,
  input        reset,
  output       io_enq_ready,
  input        io_enq_valid,
  input  [9:0] io_enq_bits,
  input        io_deq_ready,
  output       io_deq_valid,
  output [9:0] io_deq_bits,
  input  [3:0] modifyVal,
  input        modify,
  output [3:0] allocatedAddr
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [9:0] memReg [0:15]; // @[storeDataIssue.scala 31:19]
  wire  memReg_io_deq_bits_MPORT_en; // @[storeDataIssue.scala 31:19]
  wire [3:0] memReg_io_deq_bits_MPORT_addr; // @[storeDataIssue.scala 31:19]
  wire [9:0] memReg_io_deq_bits_MPORT_data; // @[storeDataIssue.scala 31:19]
  wire [9:0] memReg_MPORT_data; // @[storeDataIssue.scala 31:19]
  wire [3:0] memReg_MPORT_addr; // @[storeDataIssue.scala 31:19]
  wire  memReg_MPORT_mask; // @[storeDataIssue.scala 31:19]
  wire  memReg_MPORT_en; // @[storeDataIssue.scala 31:19]
  wire [9:0] memReg_MPORT_1_data; // @[storeDataIssue.scala 31:19]
  wire [3:0] memReg_MPORT_1_addr; // @[storeDataIssue.scala 31:19]
  wire  memReg_MPORT_1_mask; // @[storeDataIssue.scala 31:19]
  wire  memReg_MPORT_1_en; // @[storeDataIssue.scala 31:19]
  reg [3:0] readPtr; // @[storeDataIssue.scala 25:24]
  wire [3:0] _nextRead_T_2 = readPtr + 4'h1; // @[storeDataIssue.scala 26:62]
  wire [3:0] nextRead = readPtr == 4'hf ? 4'h0 : _nextRead_T_2; // @[storeDataIssue.scala 26:21]
  reg [3:0] writePtr; // @[storeDataIssue.scala 27:25]
  wire [3:0] _nextWrite_T_2 = writePtr + 4'h1; // @[storeDataIssue.scala 28:65]
  wire [3:0] nextWrite = writePtr == 4'hf ? 4'h0 : _nextWrite_T_2; // @[storeDataIssue.scala 28:22]
  reg  emptyReg; // @[storeDataIssue.scala 34:25]
  reg  fullReg; // @[storeDataIssue.scala 35:24]
  wire  _T_2 = io_deq_ready & io_deq_valid; // @[storeDataIssue.scala 64:21]
  wire  _T_3 = io_deq_ready & io_deq_valid & io_enq_valid; // @[storeDataIssue.scala 64:37]
  wire  _T_4 = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready; // @[storeDataIssue.scala 64:53]
  wire  _T_5 = io_enq_valid & io_enq_ready; // @[storeDataIssue.scala 70:27]
  wire  _GEN_110 = io_enq_valid & io_enq_ready ? 1'h0 : _T_2; // @[storeDataIssue.scala 70:44]
  wire  incrRead = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready | _GEN_110; // @[storeDataIssue.scala 64:70 69:14]
  wire  _T = ~emptyReg; // @[storeDataIssue.scala 53:19]
  wire  incrWrite = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready | _T_5; // @[storeDataIssue.scala 64:70 68:15]
  wire  _GEN_3 = modify & ~emptyReg ? modifyVal == readPtr : emptyReg; // @[storeDataIssue.scala 53:29 58:14 34:25]
  wire  _GEN_69 = _T_2 ? nextRead == writePtr : _GEN_3; // @[storeDataIssue.scala 76:44 78:14]
  wire  _GEN_108 = io_enq_valid & io_enq_ready ? 1'h0 : _GEN_69; // @[storeDataIssue.scala 70:44 73:14]
  wire  _GEN_139 = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready ? _GEN_3 : _GEN_108; // @[storeDataIssue.scala 64:70]
  wire  _io_enq_ready_T_3 = ~modify; // @[storeDataIssue.scala 84:64]
  assign memReg_io_deq_bits_MPORT_en = 1'h1;
  assign memReg_io_deq_bits_MPORT_addr = readPtr;
  assign memReg_io_deq_bits_MPORT_data = memReg[memReg_io_deq_bits_MPORT_addr]; // @[storeDataIssue.scala 31:19]
  assign memReg_MPORT_data = io_enq_bits;
  assign memReg_MPORT_addr = writePtr;
  assign memReg_MPORT_mask = 1'h1;
  assign memReg_MPORT_en = _T_3 & io_enq_ready;
  assign memReg_MPORT_1_data = io_enq_bits;
  assign memReg_MPORT_1_addr = writePtr;
  assign memReg_MPORT_1_mask = 1'h1;
  assign memReg_MPORT_1_en = _T_4 ? 1'h0 : _T_5;
  assign io_enq_ready = (~fullReg | io_deq_valid & io_deq_ready) & ~modify; // @[storeDataIssue.scala 84:62]
  assign io_deq_valid = _T & _io_enq_ready_T_3; // @[storeDataIssue.scala 85:29]
  assign io_deq_bits = memReg_io_deq_bits_MPORT_data; // @[storeDataIssue.scala 83:15]
  assign allocatedAddr = writePtr; // @[storeDataIssue.scala 92:17]
  always @(posedge clock) begin
    if (memReg_MPORT_en & memReg_MPORT_mask) begin
      memReg[memReg_MPORT_addr] <= memReg_MPORT_data; // @[storeDataIssue.scala 31:19]
    end
    if (memReg_MPORT_1_en & memReg_MPORT_1_mask) begin
      memReg[memReg_MPORT_1_addr] <= memReg_MPORT_1_data; // @[storeDataIssue.scala 31:19]
    end
    if (reset) begin // @[storeDataIssue.scala 25:24]
      readPtr <= 4'h0; // @[storeDataIssue.scala 25:24]
    end else if (incrRead) begin // @[storeDataIssue.scala 48:19]
      if (readPtr == 4'hf) begin // @[storeDataIssue.scala 26:21]
        readPtr <= 4'h0;
      end else begin
        readPtr <= _nextRead_T_2;
      end
    end
    if (reset) begin // @[storeDataIssue.scala 27:25]
      writePtr <= 4'h0; // @[storeDataIssue.scala 27:25]
    end else if (modify & ~emptyReg) begin // @[storeDataIssue.scala 53:29]
      writePtr <= modifyVal; // @[storeDataIssue.scala 56:14]
    end else if (incrWrite) begin // @[storeDataIssue.scala 59:24]
      if (writePtr == 4'hf) begin // @[storeDataIssue.scala 28:22]
        writePtr <= 4'h0;
      end else begin
        writePtr <= _nextWrite_T_2;
      end
    end
    emptyReg <= reset | _GEN_139; // @[storeDataIssue.scala 34:{25,25}]
    if (reset) begin // @[storeDataIssue.scala 35:24]
      fullReg <= 1'h0; // @[storeDataIssue.scala 35:24]
    end else if (!(io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready)) begin // @[storeDataIssue.scala 64:70]
      if (io_enq_valid & io_enq_ready) begin // @[storeDataIssue.scala 70:44]
        fullReg <= nextWrite == readPtr; // @[storeDataIssue.scala 74:13]
      end else if (_T_2) begin // @[storeDataIssue.scala 76:44]
        fullReg <= 1'h0; // @[storeDataIssue.scala 77:13]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    memReg[initvar] = _RAND_0[9:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  readPtr = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  writePtr = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  emptyReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  fullReg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module storeDataIssue(
  input        clock,
  input        reset,
  input        fromROB_readyNow,
  input        fromBranch_passOrFail,
  input  [3:0] fromBranch_robAddr,
  input        fromBranch_valid,
  output       fromDecode_ready,
  input        fromDecode_valid,
  input  [5:0] fromDecode_rs2Addr,
  input  [3:0] fromDecode_branchMask,
  output       toPRF_valid,
  output [5:0] toPRF_rs2Addr,
  input        robMapUpdate_valid,
  input  [3:0] robMapUpdate_robAddr
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  wire  sdiFifo_clock; // @[storeDataIssue.scala 146:27]
  wire  sdiFifo_reset; // @[storeDataIssue.scala 146:27]
  wire  sdiFifo_io_enq_ready; // @[storeDataIssue.scala 146:27]
  wire  sdiFifo_io_enq_valid; // @[storeDataIssue.scala 146:27]
  wire [9:0] sdiFifo_io_enq_bits; // @[storeDataIssue.scala 146:27]
  wire  sdiFifo_io_deq_ready; // @[storeDataIssue.scala 146:27]
  wire  sdiFifo_io_deq_valid; // @[storeDataIssue.scala 146:27]
  wire [9:0] sdiFifo_io_deq_bits; // @[storeDataIssue.scala 146:27]
  wire [3:0] sdiFifo_modifyVal; // @[storeDataIssue.scala 146:27]
  wire  sdiFifo_modify; // @[storeDataIssue.scala 146:27]
  wire [3:0] sdiFifo_allocatedAddr; // @[storeDataIssue.scala 146:27]
  reg [3:0] map [0:15]; // @[storeDataIssue.scala 152:16]
  wire  map_sdiFifo_modifyVal_MPORT_en; // @[storeDataIssue.scala 152:16]
  wire [3:0] map_sdiFifo_modifyVal_MPORT_addr; // @[storeDataIssue.scala 152:16]
  wire [3:0] map_sdiFifo_modifyVal_MPORT_data; // @[storeDataIssue.scala 152:16]
  wire [3:0] map_MPORT_data; // @[storeDataIssue.scala 152:16]
  wire [3:0] map_MPORT_addr; // @[storeDataIssue.scala 152:16]
  wire  map_MPORT_mask; // @[storeDataIssue.scala 152:16]
  wire  map_MPORT_en; // @[storeDataIssue.scala 152:16]
  storeDataIssue_Anon sdiFifo ( // @[storeDataIssue.scala 146:27]
    .clock(sdiFifo_clock),
    .reset(sdiFifo_reset),
    .io_enq_ready(sdiFifo_io_enq_ready),
    .io_enq_valid(sdiFifo_io_enq_valid),
    .io_enq_bits(sdiFifo_io_enq_bits),
    .io_deq_ready(sdiFifo_io_deq_ready),
    .io_deq_valid(sdiFifo_io_deq_valid),
    .io_deq_bits(sdiFifo_io_deq_bits),
    .modifyVal(sdiFifo_modifyVal),
    .modify(sdiFifo_modify),
    .allocatedAddr(sdiFifo_allocatedAddr)
  );
  assign map_sdiFifo_modifyVal_MPORT_en = 1'h1;
  assign map_sdiFifo_modifyVal_MPORT_addr = fromBranch_robAddr;
  assign map_sdiFifo_modifyVal_MPORT_data = map[map_sdiFifo_modifyVal_MPORT_addr]; // @[storeDataIssue.scala 152:16]
  assign map_MPORT_data = sdiFifo_allocatedAddr;
  assign map_MPORT_addr = robMapUpdate_robAddr;
  assign map_MPORT_mask = 1'h1;
  assign map_MPORT_en = robMapUpdate_valid;
  assign fromDecode_ready = sdiFifo_io_enq_ready; // @[storeDataIssue.scala 167:29]
  assign toPRF_valid = sdiFifo_io_deq_valid; // @[storeDataIssue.scala 179:21]
  assign toPRF_rs2Addr = sdiFifo_io_deq_bits[5:0]; // @[storeDataIssue.scala 176:43]
  assign sdiFifo_clock = clock;
  assign sdiFifo_reset = reset;
  assign sdiFifo_io_enq_valid = fromDecode_valid; // @[storeDataIssue.scala 166:29]
  assign sdiFifo_io_enq_bits = {fromDecode_branchMask,fromDecode_rs2Addr}; // @[Cat.scala 33:92]
  assign sdiFifo_io_deq_ready = fromROB_readyNow; // @[storeDataIssue.scala 172:29]
  assign sdiFifo_modifyVal = map_sdiFifo_modifyVal_MPORT_data; // @[storeDataIssue.scala 169:21]
  assign sdiFifo_modify = fromBranch_valid & ~fromBranch_passOrFail; // @[storeDataIssue.scala 170:41]
  always @(posedge clock) begin
    if (map_MPORT_en & map_MPORT_mask) begin
      map[map_MPORT_addr] <= map_MPORT_data; // @[storeDataIssue.scala 152:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    map[initvar] = _RAND_0[3:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module rob_Anon(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [101:0] io_enq_bits,
  input          io_deq_ready,
  output         io_deq_valid,
  output [101:0] io_deq_bits,
  input          modify,
  input  [3:0]   modifyVal
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [101:0] memReg [0:15]; // @[Fifo.scala 86:19]
  wire  memReg_io_deq_bits_MPORT_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_io_deq_bits_MPORT_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_io_deq_bits_MPORT_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_2_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_2_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_2_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_3_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_3_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_3_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_4_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_4_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_4_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_5_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_5_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_5_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_6_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_6_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_6_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_7_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_7_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_7_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_8_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_8_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_8_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_9_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_9_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_9_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_10_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_10_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_10_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_11_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_11_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_11_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_12_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_12_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_12_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_13_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_13_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_13_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_14_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_14_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_14_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_15_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_15_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_15_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_16_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_16_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_16_data; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_17_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_17_addr; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_17_data; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_data; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_addr; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_mask; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_en; // @[Fifo.scala 86:19]
  wire [101:0] memReg_MPORT_1_data; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_1_addr; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_1_mask; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_1_en; // @[Fifo.scala 86:19]
  reg [3:0] readPtr; // @[Fifo.scala 75:25]
  wire [3:0] _nextRead_T_2 = readPtr + 4'h1; // @[Fifo.scala 76:61]
  wire [3:0] nextRead = readPtr == 4'hf ? 4'h0 : _nextRead_T_2; // @[Fifo.scala 76:21]
  wire  _T = io_deq_ready & io_deq_valid; // @[Fifo.scala 105:21]
  wire  _T_1 = io_deq_ready & io_deq_valid & io_enq_valid; // @[Fifo.scala 105:37]
  wire  _T_2 = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready; // @[Fifo.scala 105:53]
  wire  _T_3 = io_enq_valid & io_enq_ready; // @[Fifo.scala 109:27]
  wire  _GEN_14 = io_enq_valid & io_enq_ready ? 1'h0 : _T; // @[Fifo.scala 109:44]
  wire  incrRead = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready | _GEN_14; // @[Fifo.scala 105:70 108:14]
  reg [3:0] writePtr; // @[Fifo.scala 81:25]
  wire [3:0] _nextWrite_T_2 = writePtr + 4'h1; // @[Fifo.scala 82:65]
  wire [3:0] nextWrite = writePtr == 4'hf ? 4'h0 : _nextWrite_T_2; // @[Fifo.scala 82:22]
  reg  fullReg; // @[Fifo.scala 84:24]
  reg  emptyReg; // @[Fifo.scala 89:25]
  wire [3:0] _nextval_T_2 = modifyVal + 4'h1; // @[Fifo.scala 91:65]
  wire [3:0] nextval = modifyVal == 4'hf ? 4'h0 : _nextval_T_2; // @[Fifo.scala 91:20]
  wire  incrWrite = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready | _T_3; // @[Fifo.scala 105:70 107:15]
  wire  _GEN_3 = modify ? nextval == readPtr : fullReg; // @[Fifo.scala 93:16 96:13 84:24]
  wire  _GEN_5 = _T ? nextRead == writePtr : emptyReg; // @[Fifo.scala 114:44 116:14 89:25]
  wire  _GEN_12 = io_enq_valid & io_enq_ready ? 1'h0 : _GEN_5; // @[Fifo.scala 109:44 111:14]
  wire  _GEN_27 = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready ? emptyReg : _GEN_12; // @[Fifo.scala 105:70 89:25]
  wire  _io_enq_ready_T_3 = ~modify; // @[Fifo.scala 121:64]
  assign memReg_io_deq_bits_MPORT_en = 1'h1;
  assign memReg_io_deq_bits_MPORT_addr = readPtr;
  assign memReg_io_deq_bits_MPORT_data = memReg[memReg_io_deq_bits_MPORT_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_2_en = 1'h1;
  assign memReg_MPORT_2_addr = 4'h0;
  assign memReg_MPORT_2_data = memReg[memReg_MPORT_2_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_3_en = 1'h1;
  assign memReg_MPORT_3_addr = 4'h1;
  assign memReg_MPORT_3_data = memReg[memReg_MPORT_3_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_4_en = 1'h1;
  assign memReg_MPORT_4_addr = 4'h2;
  assign memReg_MPORT_4_data = memReg[memReg_MPORT_4_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_5_en = 1'h1;
  assign memReg_MPORT_5_addr = 4'h3;
  assign memReg_MPORT_5_data = memReg[memReg_MPORT_5_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_6_en = 1'h1;
  assign memReg_MPORT_6_addr = 4'h4;
  assign memReg_MPORT_6_data = memReg[memReg_MPORT_6_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_7_en = 1'h1;
  assign memReg_MPORT_7_addr = 4'h5;
  assign memReg_MPORT_7_data = memReg[memReg_MPORT_7_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_8_en = 1'h1;
  assign memReg_MPORT_8_addr = 4'h6;
  assign memReg_MPORT_8_data = memReg[memReg_MPORT_8_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_9_en = 1'h1;
  assign memReg_MPORT_9_addr = 4'h7;
  assign memReg_MPORT_9_data = memReg[memReg_MPORT_9_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_10_en = 1'h1;
  assign memReg_MPORT_10_addr = 4'h8;
  assign memReg_MPORT_10_data = memReg[memReg_MPORT_10_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_11_en = 1'h1;
  assign memReg_MPORT_11_addr = 4'h9;
  assign memReg_MPORT_11_data = memReg[memReg_MPORT_11_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_12_en = 1'h1;
  assign memReg_MPORT_12_addr = 4'ha;
  assign memReg_MPORT_12_data = memReg[memReg_MPORT_12_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_13_en = 1'h1;
  assign memReg_MPORT_13_addr = 4'hb;
  assign memReg_MPORT_13_data = memReg[memReg_MPORT_13_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_14_en = 1'h1;
  assign memReg_MPORT_14_addr = 4'hc;
  assign memReg_MPORT_14_data = memReg[memReg_MPORT_14_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_15_en = 1'h1;
  assign memReg_MPORT_15_addr = 4'hd;
  assign memReg_MPORT_15_data = memReg[memReg_MPORT_15_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_16_en = 1'h1;
  assign memReg_MPORT_16_addr = 4'he;
  assign memReg_MPORT_16_data = memReg[memReg_MPORT_16_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_17_en = 1'h1;
  assign memReg_MPORT_17_addr = 4'hf;
  assign memReg_MPORT_17_data = memReg[memReg_MPORT_17_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_data = io_enq_bits;
  assign memReg_MPORT_addr = writePtr;
  assign memReg_MPORT_mask = 1'h1;
  assign memReg_MPORT_en = _T_1 & io_enq_ready;
  assign memReg_MPORT_1_data = io_enq_bits;
  assign memReg_MPORT_1_addr = writePtr;
  assign memReg_MPORT_1_mask = 1'h1;
  assign memReg_MPORT_1_en = _T_2 ? 1'h0 : _T_3;
  assign io_enq_ready = (~fullReg | io_deq_valid & io_deq_ready) & ~modify; // @[Fifo.scala 121:62]
  assign io_deq_valid = ~emptyReg & _io_enq_ready_T_3; // @[Fifo.scala 122:29]
  assign io_deq_bits = memReg_io_deq_bits_MPORT_data; // @[Fifo.scala 120:15]
  always @(posedge clock) begin
    if (memReg_MPORT_en & memReg_MPORT_mask) begin
      memReg[memReg_MPORT_addr] <= memReg_MPORT_data; // @[Fifo.scala 86:19]
    end
    if (memReg_MPORT_1_en & memReg_MPORT_1_mask) begin
      memReg[memReg_MPORT_1_addr] <= memReg_MPORT_1_data; // @[Fifo.scala 86:19]
    end
    if (reset) begin // @[Fifo.scala 75:25]
      readPtr <= 4'h0; // @[Fifo.scala 75:25]
    end else if (incrRead) begin // @[Fifo.scala 77:19]
      if (readPtr == 4'hf) begin // @[Fifo.scala 76:21]
        readPtr <= 4'h0;
      end else begin
        readPtr <= _nextRead_T_2;
      end
    end
    if (reset) begin // @[Fifo.scala 81:25]
      writePtr <= 4'h0; // @[Fifo.scala 81:25]
    end else if (modify) begin // @[Fifo.scala 93:16]
      if (modifyVal == 4'hf) begin // @[Fifo.scala 91:20]
        writePtr <= 4'h0;
      end else begin
        writePtr <= _nextval_T_2;
      end
    end else if (incrWrite) begin // @[Fifo.scala 98:24]
      if (writePtr == 4'hf) begin // @[Fifo.scala 82:22]
        writePtr <= 4'h0;
      end else begin
        writePtr <= _nextWrite_T_2;
      end
    end
    if (reset) begin // @[Fifo.scala 84:24]
      fullReg <= 1'h0; // @[Fifo.scala 84:24]
    end else if (io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready) begin // @[Fifo.scala 105:70]
      fullReg <= _GEN_3;
    end else if (io_enq_valid & io_enq_ready) begin // @[Fifo.scala 109:44]
      fullReg <= nextWrite == readPtr; // @[Fifo.scala 112:13]
    end else if (_T) begin // @[Fifo.scala 114:44]
      fullReg <= 1'h0; // @[Fifo.scala 115:13]
    end else begin
      fullReg <= _GEN_3;
    end
    emptyReg <= reset | _GEN_27; // @[Fifo.scala 89:{25,25}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    memReg[initvar] = _RAND_0[101:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  readPtr = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  writePtr = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  fullReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  emptyReg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module rob_Anon_1(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [129:0] io_enq_bits,
  input          io_deq_ready,
  output         io_deq_valid,
  output [129:0] io_deq_bits,
  input          modify,
  input  [3:0]   modifyVal,
  input          writeports_0_valid,
  input  [129:0] writeports_0_data,
  input  [3:0]   writeports_0_addr,
  input          writeports_1_valid,
  input  [3:0]   writeports_1_addr,
  input          writeports_2_valid,
  input  [3:0]   writeports_2_addr,
  input          writeports_3_valid,
  input  [3:0]   writeports_3_addr,
  input          writeports_4_valid,
  input  [3:0]   writeports_4_addr,
  output [3:0]   allocatedAddr,
  output [3:0]   robAddrRelease
);
`ifdef RANDOMIZE_MEM_INIT
  reg [159:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [129:0] memReg [0:15]; // @[Fifo.scala 86:19]
  wire  memReg_io_deq_bits_MPORT_en; // @[Fifo.scala 86:19]
  wire [3:0] memReg_io_deq_bits_MPORT_addr; // @[Fifo.scala 86:19]
  wire [129:0] memReg_io_deq_bits_MPORT_data; // @[Fifo.scala 86:19]
  wire [129:0] memReg_MPORT_data; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_addr; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_mask; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_en; // @[Fifo.scala 86:19]
  wire [129:0] memReg_MPORT_1_data; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_1_addr; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_1_mask; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_1_en; // @[Fifo.scala 86:19]
  wire [129:0] memReg_MPORT_2_data; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_2_addr; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_2_mask; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_2_en; // @[Fifo.scala 86:19]
  wire [129:0] memReg_MPORT_3_data; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_3_addr; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_3_mask; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_3_en; // @[Fifo.scala 86:19]
  wire [129:0] memReg_MPORT_4_data; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_4_addr; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_4_mask; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_4_en; // @[Fifo.scala 86:19]
  wire [129:0] memReg_MPORT_5_data; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_5_addr; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_5_mask; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_5_en; // @[Fifo.scala 86:19]
  wire [129:0] memReg_MPORT_6_data; // @[Fifo.scala 86:19]
  wire [3:0] memReg_MPORT_6_addr; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_6_mask; // @[Fifo.scala 86:19]
  wire  memReg_MPORT_6_en; // @[Fifo.scala 86:19]
  reg [3:0] readPtr; // @[Fifo.scala 75:25]
  wire [3:0] _nextRead_T_2 = readPtr + 4'h1; // @[Fifo.scala 76:61]
  wire [3:0] nextRead = readPtr == 4'hf ? 4'h0 : _nextRead_T_2; // @[Fifo.scala 76:21]
  wire  _T = io_deq_ready & io_deq_valid; // @[Fifo.scala 105:21]
  wire  _T_1 = io_deq_ready & io_deq_valid & io_enq_valid; // @[Fifo.scala 105:37]
  wire  _T_2 = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready; // @[Fifo.scala 105:53]
  wire  _T_3 = io_enq_valid & io_enq_ready; // @[Fifo.scala 109:27]
  wire  _GEN_14 = io_enq_valid & io_enq_ready ? 1'h0 : _T; // @[Fifo.scala 109:44]
  wire  incrRead = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready | _GEN_14; // @[Fifo.scala 105:70 108:14]
  reg [3:0] writePtr; // @[Fifo.scala 81:25]
  wire [3:0] _nextWrite_T_2 = writePtr + 4'h1; // @[Fifo.scala 82:65]
  wire [3:0] nextWrite = writePtr == 4'hf ? 4'h0 : _nextWrite_T_2; // @[Fifo.scala 82:22]
  reg  fullReg; // @[Fifo.scala 84:24]
  reg  emptyReg; // @[Fifo.scala 89:25]
  wire [3:0] _nextval_T_2 = modifyVal + 4'h1; // @[Fifo.scala 91:65]
  wire [3:0] nextval = modifyVal == 4'hf ? 4'h0 : _nextval_T_2; // @[Fifo.scala 91:20]
  wire  incrWrite = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready | _T_3; // @[Fifo.scala 105:70 107:15]
  wire  _GEN_3 = modify ? nextval == readPtr : fullReg; // @[Fifo.scala 93:16 96:13 84:24]
  wire  _GEN_5 = _T ? nextRead == writePtr : emptyReg; // @[Fifo.scala 114:44 116:14 89:25]
  wire  _GEN_12 = io_enq_valid & io_enq_ready ? 1'h0 : _GEN_5; // @[Fifo.scala 109:44 111:14]
  wire  _GEN_27 = io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready ? emptyReg : _GEN_12; // @[Fifo.scala 105:70 89:25]
  wire  _io_enq_ready_T_3 = ~modify; // @[Fifo.scala 121:64]
  assign memReg_io_deq_bits_MPORT_en = 1'h1;
  assign memReg_io_deq_bits_MPORT_addr = readPtr;
  assign memReg_io_deq_bits_MPORT_data = memReg[memReg_io_deq_bits_MPORT_addr]; // @[Fifo.scala 86:19]
  assign memReg_MPORT_data = io_enq_bits;
  assign memReg_MPORT_addr = writePtr;
  assign memReg_MPORT_mask = 1'h1;
  assign memReg_MPORT_en = _T_1 & io_enq_ready;
  assign memReg_MPORT_1_data = io_enq_bits;
  assign memReg_MPORT_1_addr = writePtr;
  assign memReg_MPORT_1_mask = 1'h1;
  assign memReg_MPORT_1_en = _T_2 ? 1'h0 : _T_3;
  assign memReg_MPORT_2_data = writeports_0_data;
  assign memReg_MPORT_2_addr = writeports_0_addr;
  assign memReg_MPORT_2_mask = 1'h1;
  assign memReg_MPORT_2_en = writeports_0_valid;
  assign memReg_MPORT_3_data = 130'h1;
  assign memReg_MPORT_3_addr = writeports_1_addr;
  assign memReg_MPORT_3_mask = 1'h1;
  assign memReg_MPORT_3_en = writeports_1_valid;
  assign memReg_MPORT_4_data = 130'h1;
  assign memReg_MPORT_4_addr = writeports_2_addr;
  assign memReg_MPORT_4_mask = 1'h1;
  assign memReg_MPORT_4_en = writeports_2_valid;
  assign memReg_MPORT_5_data = 130'h1;
  assign memReg_MPORT_5_addr = writeports_3_addr;
  assign memReg_MPORT_5_mask = 1'h1;
  assign memReg_MPORT_5_en = writeports_3_valid;
  assign memReg_MPORT_6_data = 130'h1;
  assign memReg_MPORT_6_addr = writeports_4_addr;
  assign memReg_MPORT_6_mask = 1'h1;
  assign memReg_MPORT_6_en = writeports_4_valid;
  assign io_enq_ready = (~fullReg | io_deq_valid & io_deq_ready) & ~modify; // @[Fifo.scala 121:62]
  assign io_deq_valid = ~emptyReg & _io_enq_ready_T_3; // @[Fifo.scala 122:29]
  assign io_deq_bits = memReg_io_deq_bits_MPORT_data; // @[Fifo.scala 120:15]
  assign allocatedAddr = writePtr; // @[Fifo.scala 145:17]
  assign robAddrRelease = readPtr; // @[rob.scala 63:20]
  always @(posedge clock) begin
    if (memReg_MPORT_en & memReg_MPORT_mask) begin
      memReg[memReg_MPORT_addr] <= memReg_MPORT_data; // @[Fifo.scala 86:19]
    end
    if (memReg_MPORT_1_en & memReg_MPORT_1_mask) begin
      memReg[memReg_MPORT_1_addr] <= memReg_MPORT_1_data; // @[Fifo.scala 86:19]
    end
    if (memReg_MPORT_2_en & memReg_MPORT_2_mask) begin
      memReg[memReg_MPORT_2_addr] <= memReg_MPORT_2_data; // @[Fifo.scala 86:19]
    end
    if (memReg_MPORT_3_en & memReg_MPORT_3_mask) begin
      memReg[memReg_MPORT_3_addr] <= memReg_MPORT_3_data; // @[Fifo.scala 86:19]
    end
    if (memReg_MPORT_4_en & memReg_MPORT_4_mask) begin
      memReg[memReg_MPORT_4_addr] <= memReg_MPORT_4_data; // @[Fifo.scala 86:19]
    end
    if (memReg_MPORT_5_en & memReg_MPORT_5_mask) begin
      memReg[memReg_MPORT_5_addr] <= memReg_MPORT_5_data; // @[Fifo.scala 86:19]
    end
    if (memReg_MPORT_6_en & memReg_MPORT_6_mask) begin
      memReg[memReg_MPORT_6_addr] <= memReg_MPORT_6_data; // @[Fifo.scala 86:19]
    end
    if (reset) begin // @[Fifo.scala 75:25]
      readPtr <= 4'h0; // @[Fifo.scala 75:25]
    end else if (incrRead) begin // @[Fifo.scala 77:19]
      if (readPtr == 4'hf) begin // @[Fifo.scala 76:21]
        readPtr <= 4'h0;
      end else begin
        readPtr <= _nextRead_T_2;
      end
    end
    if (reset) begin // @[Fifo.scala 81:25]
      writePtr <= 4'h0; // @[Fifo.scala 81:25]
    end else if (modify) begin // @[Fifo.scala 93:16]
      if (modifyVal == 4'hf) begin // @[Fifo.scala 91:20]
        writePtr <= 4'h0;
      end else begin
        writePtr <= _nextval_T_2;
      end
    end else if (incrWrite) begin // @[Fifo.scala 98:24]
      if (writePtr == 4'hf) begin // @[Fifo.scala 82:22]
        writePtr <= 4'h0;
      end else begin
        writePtr <= _nextWrite_T_2;
      end
    end
    if (reset) begin // @[Fifo.scala 84:24]
      fullReg <= 1'h0; // @[Fifo.scala 84:24]
    end else if (io_deq_ready & io_deq_valid & io_enq_valid & io_enq_ready) begin // @[Fifo.scala 105:70]
      fullReg <= _GEN_3;
    end else if (io_enq_valid & io_enq_ready) begin // @[Fifo.scala 109:44]
      fullReg <= nextWrite == readPtr; // @[Fifo.scala 112:13]
    end else if (_T) begin // @[Fifo.scala 114:44]
      fullReg <= 1'h0; // @[Fifo.scala 115:13]
    end else begin
      fullReg <= _GEN_3;
    end
    emptyReg <= reset | _GEN_27; // @[Fifo.scala 89:{25,25}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {5{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    memReg[initvar] = _RAND_0[129:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  readPtr = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  writePtr = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  fullReg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  emptyReg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module rob(
  input         clock,
  input         reset,
  output        allocate_ready,
  input         allocate_fired,
  input  [63:0] allocate_pc,
  input  [31:0] allocate_instruction,
  input  [5:0]  allocate_prfDest,
  output [3:0]  allocate_robAddr,
  input         allocate_isReady,
  output        commit_ready,
  input         commit_fired,
  output [5:0]  commit_prfDest,
  output [31:0] commit_instruction,
  output        commit_exceptionOccurred,
  output [63:0] commit_mtval,
  output        commit_isStore,
  output        commit_is_fence,
  output [3:0]  commit_robAddr,
  input         branch_valid,
  input         branch_pass,
  input  [3:0]  branch_robAddr,
  input  [3:0]  execPorts_0_robAddr,
  input  [63:0] execPorts_0_mtval,
  input         execPorts_0_valid,
  input  [3:0]  execPorts_1_robAddr,
  input         execPorts_1_valid,
  input  [3:0]  execPorts_2_robAddr,
  input         execPorts_2_valid,
  input  [3:0]  execPorts_3_robAddr,
  input         execPorts_3_valid
);
  wire  fifo_clock; // @[rob.scala 24:20]
  wire  fifo_reset; // @[rob.scala 24:20]
  wire  fifo_io_enq_ready; // @[rob.scala 24:20]
  wire  fifo_io_enq_valid; // @[rob.scala 24:20]
  wire [101:0] fifo_io_enq_bits; // @[rob.scala 24:20]
  wire  fifo_io_deq_ready; // @[rob.scala 24:20]
  wire  fifo_io_deq_valid; // @[rob.scala 24:20]
  wire [101:0] fifo_io_deq_bits; // @[rob.scala 24:20]
  wire  fifo_modify; // @[rob.scala 24:20]
  wire [3:0] fifo_modifyVal; // @[rob.scala 24:20]
  wire  results_clock; // @[rob.scala 61:23]
  wire  results_reset; // @[rob.scala 61:23]
  wire  results_io_enq_ready; // @[rob.scala 61:23]
  wire  results_io_enq_valid; // @[rob.scala 61:23]
  wire [129:0] results_io_enq_bits; // @[rob.scala 61:23]
  wire  results_io_deq_ready; // @[rob.scala 61:23]
  wire  results_io_deq_valid; // @[rob.scala 61:23]
  wire [129:0] results_io_deq_bits; // @[rob.scala 61:23]
  wire  results_modify; // @[rob.scala 61:23]
  wire [3:0] results_modifyVal; // @[rob.scala 61:23]
  wire  results_writeports_0_valid; // @[rob.scala 61:23]
  wire [129:0] results_writeports_0_data; // @[rob.scala 61:23]
  wire [3:0] results_writeports_0_addr; // @[rob.scala 61:23]
  wire  results_writeports_1_valid; // @[rob.scala 61:23]
  wire [3:0] results_writeports_1_addr; // @[rob.scala 61:23]
  wire  results_writeports_2_valid; // @[rob.scala 61:23]
  wire [3:0] results_writeports_2_addr; // @[rob.scala 61:23]
  wire  results_writeports_3_valid; // @[rob.scala 61:23]
  wire [3:0] results_writeports_3_addr; // @[rob.scala 61:23]
  wire  results_writeports_4_valid; // @[rob.scala 61:23]
  wire [3:0] results_writeports_4_addr; // @[rob.scala 61:23]
  wire [3:0] results_allocatedAddr; // @[rob.scala 61:23]
  wire [3:0] results_robAddrRelease; // @[rob.scala 61:23]
  wire [37:0] _fifo_data_T = {allocate_instruction,allocate_prfDest}; // @[Cat.scala 33:92]
  wire  is_fence = commit_instruction[6:0] == 7'hf; // @[rob.scala 81:42]
  wire  _fifo_modify_T = ~branch_pass; // @[rob.scala 105:33]
  wire [128:0] _writeval_T_1 = {execPorts_0_mtval,65'h1}; // @[Cat.scala 33:92]
  rob_Anon fifo ( // @[rob.scala 24:20]
    .clock(fifo_clock),
    .reset(fifo_reset),
    .io_enq_ready(fifo_io_enq_ready),
    .io_enq_valid(fifo_io_enq_valid),
    .io_enq_bits(fifo_io_enq_bits),
    .io_deq_ready(fifo_io_deq_ready),
    .io_deq_valid(fifo_io_deq_valid),
    .io_deq_bits(fifo_io_deq_bits),
    .modify(fifo_modify),
    .modifyVal(fifo_modifyVal)
  );
  rob_Anon_1 results ( // @[rob.scala 61:23]
    .clock(results_clock),
    .reset(results_reset),
    .io_enq_ready(results_io_enq_ready),
    .io_enq_valid(results_io_enq_valid),
    .io_enq_bits(results_io_enq_bits),
    .io_deq_ready(results_io_deq_ready),
    .io_deq_valid(results_io_deq_valid),
    .io_deq_bits(results_io_deq_bits),
    .modify(results_modify),
    .modifyVal(results_modifyVal),
    .writeports_0_valid(results_writeports_0_valid),
    .writeports_0_data(results_writeports_0_data),
    .writeports_0_addr(results_writeports_0_addr),
    .writeports_1_valid(results_writeports_1_valid),
    .writeports_1_addr(results_writeports_1_addr),
    .writeports_2_valid(results_writeports_2_valid),
    .writeports_2_addr(results_writeports_2_addr),
    .writeports_3_valid(results_writeports_3_valid),
    .writeports_3_addr(results_writeports_3_addr),
    .writeports_4_valid(results_writeports_4_valid),
    .writeports_4_addr(results_writeports_4_addr),
    .allocatedAddr(results_allocatedAddr),
    .robAddrRelease(results_robAddrRelease)
  );
  assign allocate_ready = commit_ready & ~commit_fired ? 1'h0 : fifo_io_enq_ready & results_io_enq_ready; // @[rob.scala 142:{39,56} 67:18]
  assign allocate_robAddr = results_allocatedAddr; // @[rob.scala 72:20]
  assign commit_ready = (results_io_deq_bits[0] | is_fence | commit_isStore) & fifo_io_deq_valid & results_io_deq_valid; // @[rob.scala 84:92]
  assign commit_prfDest = fifo_io_deq_bits[5:0]; // @[rob.scala 88:37]
  assign commit_instruction = fifo_io_deq_bits[37:6]; // @[rob.scala 89:41]
  assign commit_exceptionOccurred = results_io_deq_bits[129]; // @[rob.scala 87:50]
  assign commit_mtval = results_io_deq_bits[128:65]; // @[rob.scala 86:38]
  assign commit_isStore = fifo_io_deq_bits[12:6] == 7'h23; // @[rob.scala 102:44]
  assign commit_is_fence = commit_instruction[6:0] == 7'hf; // @[rob.scala 81:42]
  assign commit_robAddr = results_robAddrRelease; // @[rob.scala 92:18]
  assign fifo_clock = clock;
  assign fifo_reset = commit_exceptionOccurred & commit_fired | reset; // @[rob.scala 123:49 124:19]
  assign fifo_io_enq_valid = allocate_fired; // @[rob.scala 73:23 74:23 77:23]
  assign fifo_io_enq_bits = {allocate_pc,_fifo_data_T}; // @[Cat.scala 33:92]
  assign fifo_io_deq_ready = commit_fired; // @[rob.scala 94:22 95:23 98:23]
  assign fifo_modify = branch_valid & ~branch_pass; // @[rob.scala 105:31]
  assign fifo_modifyVal = branch_robAddr; // @[rob.scala 106:18]
  assign results_clock = clock;
  assign results_reset = commit_exceptionOccurred & commit_fired | reset; // @[rob.scala 123:49 124:19]
  assign results_io_enq_valid = allocate_fired; // @[rob.scala 73:23 74:23 77:23]
  assign results_io_enq_bits = {129'h0,allocate_isReady}; // @[Cat.scala 33:92]
  assign results_io_deq_ready = commit_fired; // @[rob.scala 94:22 95:23 98:23]
  assign results_modify = branch_valid & _fifo_modify_T; // @[rob.scala 107:34]
  assign results_modifyVal = branch_robAddr; // @[rob.scala 108:21]
  assign results_writeports_0_valid = execPorts_0_valid; // @[rob.scala 117:33]
  assign results_writeports_0_data = {1'h0,_writeval_T_1}; // @[Cat.scala 33:92]
  assign results_writeports_0_addr = execPorts_0_robAddr; // @[rob.scala 119:32]
  assign results_writeports_1_valid = execPorts_1_valid; // @[rob.scala 117:33]
  assign results_writeports_1_addr = execPorts_1_robAddr; // @[rob.scala 119:32]
  assign results_writeports_2_valid = execPorts_2_valid; // @[rob.scala 117:33]
  assign results_writeports_2_addr = execPorts_2_robAddr; // @[rob.scala 119:32]
  assign results_writeports_3_valid = execPorts_3_valid; // @[rob.scala 117:33]
  assign results_writeports_3_addr = execPorts_3_robAddr; // @[rob.scala 119:32]
  assign results_writeports_4_valid = branch_valid; // @[rob.scala 109:43]
  assign results_writeports_4_addr = branch_robAddr; // @[rob.scala 110:42]
endmodule
module scheduler(
  input         clock,
  input         reset,
  output        allocate_ready,
  input         allocate_fired,
  input  [31:0] allocate_instruction,
  input  [3:0]  allocate_branchMask,
  input         allocate_rs1_ready,
  input  [5:0]  allocate_rs1_prfAddr,
  input         allocate_rs2_ready,
  input  [5:0]  allocate_rs2_prfAddr,
  input  [5:0]  allocate_prfDest,
  input  [3:0]  allocate_robAddr,
  output        release_ready,
  input         release_fired,
  output [31:0] release_instruction,
  output [3:0]  release_branchMask,
  output [5:0]  release_rs1prfAddr,
  output [5:0]  release_rs2prfAddr,
  output [5:0]  release_prfDest,
  output [3:0]  release_robAddr,
  input         wakeUpExt_0_valid,
  input  [5:0]  wakeUpExt_0_prfAddr,
  input         wakeUpExt_1_valid,
  input  [5:0]  wakeUpExt_1_prfAddr,
  input         branchOps_valid,
  input  [3:0]  branchOps_branchMask,
  input         branchOps_passed,
  input         memoryReady,
  input         multuplyAndDivideReady,
  output        instrRetired_valid,
  output [5:0]  instrRetired_prfAddr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
`endif // RANDOMIZE_REG_INIT
  reg  queue_0_opcodeMeta_isBranch; // @[scheduler.scala 26:22]
  reg  queue_0_opcodeMeta_isMemAccess; // @[scheduler.scala 26:22]
  reg  queue_0_opcodeMeta_isM; // @[scheduler.scala 26:22]
  reg  queue_0_valid; // @[scheduler.scala 26:22]
  reg [31:0] queue_0_instruction; // @[scheduler.scala 26:22]
  reg [3:0] queue_0_branchMask; // @[scheduler.scala 26:22]
  reg  queue_0_rs1_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_0_rs1_prfAddr; // @[scheduler.scala 26:22]
  reg  queue_0_rs2_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_0_rs2_prfAddr; // @[scheduler.scala 26:22]
  reg [5:0] queue_0_prfDest; // @[scheduler.scala 26:22]
  reg [3:0] queue_0_robAddr; // @[scheduler.scala 26:22]
  reg  queue_1_opcodeMeta_isBranch; // @[scheduler.scala 26:22]
  reg  queue_1_opcodeMeta_isMemAccess; // @[scheduler.scala 26:22]
  reg  queue_1_opcodeMeta_isM; // @[scheduler.scala 26:22]
  reg  queue_1_valid; // @[scheduler.scala 26:22]
  reg [31:0] queue_1_instruction; // @[scheduler.scala 26:22]
  reg [3:0] queue_1_branchMask; // @[scheduler.scala 26:22]
  reg  queue_1_rs1_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_1_rs1_prfAddr; // @[scheduler.scala 26:22]
  reg  queue_1_rs2_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_1_rs2_prfAddr; // @[scheduler.scala 26:22]
  reg [5:0] queue_1_prfDest; // @[scheduler.scala 26:22]
  reg [3:0] queue_1_robAddr; // @[scheduler.scala 26:22]
  reg  queue_2_opcodeMeta_isBranch; // @[scheduler.scala 26:22]
  reg  queue_2_opcodeMeta_isMemAccess; // @[scheduler.scala 26:22]
  reg  queue_2_opcodeMeta_isM; // @[scheduler.scala 26:22]
  reg  queue_2_valid; // @[scheduler.scala 26:22]
  reg [31:0] queue_2_instruction; // @[scheduler.scala 26:22]
  reg [3:0] queue_2_branchMask; // @[scheduler.scala 26:22]
  reg  queue_2_rs1_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_2_rs1_prfAddr; // @[scheduler.scala 26:22]
  reg  queue_2_rs2_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_2_rs2_prfAddr; // @[scheduler.scala 26:22]
  reg [5:0] queue_2_prfDest; // @[scheduler.scala 26:22]
  reg [3:0] queue_2_robAddr; // @[scheduler.scala 26:22]
  reg  queue_3_opcodeMeta_isBranch; // @[scheduler.scala 26:22]
  reg  queue_3_opcodeMeta_isMemAccess; // @[scheduler.scala 26:22]
  reg  queue_3_opcodeMeta_isM; // @[scheduler.scala 26:22]
  reg  queue_3_valid; // @[scheduler.scala 26:22]
  reg [31:0] queue_3_instruction; // @[scheduler.scala 26:22]
  reg [3:0] queue_3_branchMask; // @[scheduler.scala 26:22]
  reg  queue_3_rs1_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_3_rs1_prfAddr; // @[scheduler.scala 26:22]
  reg  queue_3_rs2_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_3_rs2_prfAddr; // @[scheduler.scala 26:22]
  reg [5:0] queue_3_prfDest; // @[scheduler.scala 26:22]
  reg [3:0] queue_3_robAddr; // @[scheduler.scala 26:22]
  reg  queue_4_opcodeMeta_isBranch; // @[scheduler.scala 26:22]
  reg  queue_4_opcodeMeta_isMemAccess; // @[scheduler.scala 26:22]
  reg  queue_4_opcodeMeta_isM; // @[scheduler.scala 26:22]
  reg  queue_4_valid; // @[scheduler.scala 26:22]
  reg [31:0] queue_4_instruction; // @[scheduler.scala 26:22]
  reg [3:0] queue_4_branchMask; // @[scheduler.scala 26:22]
  reg  queue_4_rs1_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_4_rs1_prfAddr; // @[scheduler.scala 26:22]
  reg  queue_4_rs2_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_4_rs2_prfAddr; // @[scheduler.scala 26:22]
  reg [5:0] queue_4_prfDest; // @[scheduler.scala 26:22]
  reg [3:0] queue_4_robAddr; // @[scheduler.scala 26:22]
  reg  queue_5_opcodeMeta_isBranch; // @[scheduler.scala 26:22]
  reg  queue_5_opcodeMeta_isMemAccess; // @[scheduler.scala 26:22]
  reg  queue_5_opcodeMeta_isM; // @[scheduler.scala 26:22]
  reg  queue_5_valid; // @[scheduler.scala 26:22]
  reg [31:0] queue_5_instruction; // @[scheduler.scala 26:22]
  reg [3:0] queue_5_branchMask; // @[scheduler.scala 26:22]
  reg  queue_5_rs1_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_5_rs1_prfAddr; // @[scheduler.scala 26:22]
  reg  queue_5_rs2_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_5_rs2_prfAddr; // @[scheduler.scala 26:22]
  reg [5:0] queue_5_prfDest; // @[scheduler.scala 26:22]
  reg [3:0] queue_5_robAddr; // @[scheduler.scala 26:22]
  reg  queue_6_opcodeMeta_isBranch; // @[scheduler.scala 26:22]
  reg  queue_6_opcodeMeta_isMemAccess; // @[scheduler.scala 26:22]
  reg  queue_6_opcodeMeta_isM; // @[scheduler.scala 26:22]
  reg  queue_6_valid; // @[scheduler.scala 26:22]
  reg [31:0] queue_6_instruction; // @[scheduler.scala 26:22]
  reg [3:0] queue_6_branchMask; // @[scheduler.scala 26:22]
  reg  queue_6_rs1_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_6_rs1_prfAddr; // @[scheduler.scala 26:22]
  reg  queue_6_rs2_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_6_rs2_prfAddr; // @[scheduler.scala 26:22]
  reg [5:0] queue_6_prfDest; // @[scheduler.scala 26:22]
  reg [3:0] queue_6_robAddr; // @[scheduler.scala 26:22]
  reg  queue_7_opcodeMeta_isBranch; // @[scheduler.scala 26:22]
  reg  queue_7_opcodeMeta_isMemAccess; // @[scheduler.scala 26:22]
  reg  queue_7_opcodeMeta_isM; // @[scheduler.scala 26:22]
  reg  queue_7_valid; // @[scheduler.scala 26:22]
  reg [31:0] queue_7_instruction; // @[scheduler.scala 26:22]
  reg [3:0] queue_7_branchMask; // @[scheduler.scala 26:22]
  reg  queue_7_rs1_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_7_rs1_prfAddr; // @[scheduler.scala 26:22]
  reg  queue_7_rs2_ready; // @[scheduler.scala 26:22]
  reg [5:0] queue_7_rs2_prfAddr; // @[scheduler.scala 26:22]
  reg [5:0] queue_7_prfDest; // @[scheduler.scala 26:22]
  reg [3:0] queue_7_robAddr; // @[scheduler.scala 26:22]
  wire  _readyVector_T_1 = queue_0_valid & queue_0_rs1_ready & queue_0_rs2_ready; // @[scheduler.scala 51:42]
  wire  _readyVector_T_7 = ~queue_0_opcodeMeta_isMemAccess | memoryReady; // @[scheduler.scala 53:39]
  wire  _readyVector_T_8 = _readyVector_T_1 & _readyVector_T_7; // @[scheduler.scala 52:151]
  wire  _readyVector_T_10 = ~queue_0_opcodeMeta_isM | multuplyAndDivideReady; // @[scheduler.scala 54:31]
  wire  _readyVector_T_11 = _readyVector_T_8 & _readyVector_T_10; // @[scheduler.scala 53:174]
  wire  _readyVector_T_17 = ~queue_1_opcodeMeta_isBranch | ~(queue_0_valid & queue_0_opcodeMeta_isBranch); // @[scheduler.scala 52:36]
  wire  _readyVector_T_18 = queue_1_valid & queue_1_rs1_ready & queue_1_rs2_ready & _readyVector_T_17; // @[scheduler.scala 51:64]
  wire  _readyVector_T_23 = ~queue_1_opcodeMeta_isMemAccess | ~(queue_0_valid & queue_0_opcodeMeta_isMemAccess) &
    memoryReady; // @[scheduler.scala 53:39]
  wire  _readyVector_T_24 = _readyVector_T_18 & _readyVector_T_23; // @[scheduler.scala 52:151]
  wire  _readyVector_T_26 = ~queue_1_opcodeMeta_isM | multuplyAndDivideReady; // @[scheduler.scala 54:31]
  wire  _readyVector_T_27 = _readyVector_T_24 & _readyVector_T_26; // @[scheduler.scala 53:174]
  wire  _readyVector_T_35 = ~queue_2_opcodeMeta_isBranch | ~(queue_0_valid & queue_0_opcodeMeta_isBranch | queue_1_valid
     & queue_1_opcodeMeta_isBranch); // @[scheduler.scala 52:36]
  wire  _readyVector_T_36 = queue_2_valid & queue_2_rs1_ready & queue_2_rs2_ready & _readyVector_T_35; // @[scheduler.scala 51:64]
  wire  _readyVector_T_43 = ~queue_2_opcodeMeta_isMemAccess | ~(queue_0_valid & queue_0_opcodeMeta_isMemAccess |
    queue_1_valid & queue_1_opcodeMeta_isMemAccess) & memoryReady; // @[scheduler.scala 53:39]
  wire  _readyVector_T_44 = _readyVector_T_36 & _readyVector_T_43; // @[scheduler.scala 52:151]
  wire  _readyVector_T_46 = ~queue_2_opcodeMeta_isM | multuplyAndDivideReady; // @[scheduler.scala 54:31]
  wire  _readyVector_T_47 = _readyVector_T_44 & _readyVector_T_46; // @[scheduler.scala 53:174]
  wire  _readyVector_T_57 = ~queue_3_opcodeMeta_isBranch | ~(queue_0_valid & queue_0_opcodeMeta_isBranch | queue_1_valid
     & queue_1_opcodeMeta_isBranch | queue_2_valid & queue_2_opcodeMeta_isBranch); // @[scheduler.scala 52:36]
  wire  _readyVector_T_58 = queue_3_valid & queue_3_rs1_ready & queue_3_rs2_ready & _readyVector_T_57; // @[scheduler.scala 51:64]
  wire  _readyVector_T_67 = ~queue_3_opcodeMeta_isMemAccess | ~(queue_0_valid & queue_0_opcodeMeta_isMemAccess |
    queue_1_valid & queue_1_opcodeMeta_isMemAccess | queue_2_valid & queue_2_opcodeMeta_isMemAccess) & memoryReady; // @[scheduler.scala 53:39]
  wire  _readyVector_T_68 = _readyVector_T_58 & _readyVector_T_67; // @[scheduler.scala 52:151]
  wire  _readyVector_T_70 = ~queue_3_opcodeMeta_isM | multuplyAndDivideReady; // @[scheduler.scala 54:31]
  wire  _readyVector_T_71 = _readyVector_T_68 & _readyVector_T_70; // @[scheduler.scala 53:174]
  wire  _readyVector_T_83 = ~queue_4_opcodeMeta_isBranch | ~(queue_0_valid & queue_0_opcodeMeta_isBranch | queue_1_valid
     & queue_1_opcodeMeta_isBranch | queue_2_valid & queue_2_opcodeMeta_isBranch | queue_3_valid &
    queue_3_opcodeMeta_isBranch); // @[scheduler.scala 52:36]
  wire  _readyVector_T_84 = queue_4_valid & queue_4_rs1_ready & queue_4_rs2_ready & _readyVector_T_83; // @[scheduler.scala 51:64]
  wire  _readyVector_T_95 = ~queue_4_opcodeMeta_isMemAccess | ~(queue_0_valid & queue_0_opcodeMeta_isMemAccess |
    queue_1_valid & queue_1_opcodeMeta_isMemAccess | queue_2_valid & queue_2_opcodeMeta_isMemAccess | queue_3_valid &
    queue_3_opcodeMeta_isMemAccess) & memoryReady; // @[scheduler.scala 53:39]
  wire  _readyVector_T_96 = _readyVector_T_84 & _readyVector_T_95; // @[scheduler.scala 52:151]
  wire  _readyVector_T_98 = ~queue_4_opcodeMeta_isM | multuplyAndDivideReady; // @[scheduler.scala 54:31]
  wire  _readyVector_T_99 = _readyVector_T_96 & _readyVector_T_98; // @[scheduler.scala 53:174]
  wire  _readyVector_T_113 = ~queue_5_opcodeMeta_isBranch | ~(queue_0_valid & queue_0_opcodeMeta_isBranch |
    queue_1_valid & queue_1_opcodeMeta_isBranch | queue_2_valid & queue_2_opcodeMeta_isBranch | queue_3_valid &
    queue_3_opcodeMeta_isBranch | queue_4_valid & queue_4_opcodeMeta_isBranch); // @[scheduler.scala 52:36]
  wire  _readyVector_T_114 = queue_5_valid & queue_5_rs1_ready & queue_5_rs2_ready & _readyVector_T_113; // @[scheduler.scala 51:64]
  wire  _readyVector_T_127 = ~queue_5_opcodeMeta_isMemAccess | ~(queue_0_valid & queue_0_opcodeMeta_isMemAccess |
    queue_1_valid & queue_1_opcodeMeta_isMemAccess | queue_2_valid & queue_2_opcodeMeta_isMemAccess | queue_3_valid &
    queue_3_opcodeMeta_isMemAccess | queue_4_valid & queue_4_opcodeMeta_isMemAccess) & memoryReady; // @[scheduler.scala 53:39]
  wire  _readyVector_T_128 = _readyVector_T_114 & _readyVector_T_127; // @[scheduler.scala 52:151]
  wire  _readyVector_T_130 = ~queue_5_opcodeMeta_isM | multuplyAndDivideReady; // @[scheduler.scala 54:31]
  wire  _readyVector_T_131 = _readyVector_T_128 & _readyVector_T_130; // @[scheduler.scala 53:174]
  wire  _readyVector_T_147 = ~queue_6_opcodeMeta_isBranch | ~(queue_0_valid & queue_0_opcodeMeta_isBranch |
    queue_1_valid & queue_1_opcodeMeta_isBranch | queue_2_valid & queue_2_opcodeMeta_isBranch | queue_3_valid &
    queue_3_opcodeMeta_isBranch | queue_4_valid & queue_4_opcodeMeta_isBranch | queue_5_valid &
    queue_5_opcodeMeta_isBranch); // @[scheduler.scala 52:36]
  wire  _readyVector_T_148 = queue_6_valid & queue_6_rs1_ready & queue_6_rs2_ready & _readyVector_T_147; // @[scheduler.scala 51:64]
  wire  _readyVector_T_163 = ~queue_6_opcodeMeta_isMemAccess | ~(queue_0_valid & queue_0_opcodeMeta_isMemAccess |
    queue_1_valid & queue_1_opcodeMeta_isMemAccess | queue_2_valid & queue_2_opcodeMeta_isMemAccess | queue_3_valid &
    queue_3_opcodeMeta_isMemAccess | queue_4_valid & queue_4_opcodeMeta_isMemAccess | queue_5_valid &
    queue_5_opcodeMeta_isMemAccess) & memoryReady; // @[scheduler.scala 53:39]
  wire  _readyVector_T_164 = _readyVector_T_148 & _readyVector_T_163; // @[scheduler.scala 52:151]
  wire  _readyVector_T_166 = ~queue_6_opcodeMeta_isM | multuplyAndDivideReady; // @[scheduler.scala 54:31]
  wire  _readyVector_T_167 = _readyVector_T_164 & _readyVector_T_166; // @[scheduler.scala 53:174]
  wire  _readyVector_T_185 = ~queue_7_opcodeMeta_isBranch | ~(queue_0_valid & queue_0_opcodeMeta_isBranch |
    queue_1_valid & queue_1_opcodeMeta_isBranch | queue_2_valid & queue_2_opcodeMeta_isBranch | queue_3_valid &
    queue_3_opcodeMeta_isBranch | queue_4_valid & queue_4_opcodeMeta_isBranch | queue_5_valid &
    queue_5_opcodeMeta_isBranch | queue_6_valid & queue_6_opcodeMeta_isBranch); // @[scheduler.scala 52:36]
  wire  _readyVector_T_186 = queue_7_valid & queue_7_rs1_ready & queue_7_rs2_ready & _readyVector_T_185; // @[scheduler.scala 51:64]
  wire  _readyVector_T_203 = ~queue_7_opcodeMeta_isMemAccess | ~(queue_0_valid & queue_0_opcodeMeta_isMemAccess |
    queue_1_valid & queue_1_opcodeMeta_isMemAccess | queue_2_valid & queue_2_opcodeMeta_isMemAccess | queue_3_valid &
    queue_3_opcodeMeta_isMemAccess | queue_4_valid & queue_4_opcodeMeta_isMemAccess | queue_5_valid &
    queue_5_opcodeMeta_isMemAccess | queue_6_valid & queue_6_opcodeMeta_isMemAccess) & memoryReady; // @[scheduler.scala 53:39]
  wire  _readyVector_T_204 = _readyVector_T_186 & _readyVector_T_203; // @[scheduler.scala 52:151]
  wire  _readyVector_T_206 = ~queue_7_opcodeMeta_isM | multuplyAndDivideReady; // @[scheduler.scala 54:31]
  wire  _readyVector_T_207 = _readyVector_T_204 & _readyVector_T_206; // @[scheduler.scala 53:174]
  wire [7:0] readyVector = {_readyVector_T_207,_readyVector_T_167,_readyVector_T_131,_readyVector_T_99,_readyVector_T_71
    ,_readyVector_T_47,_readyVector_T_27,_readyVector_T_11}; // @[Cat.scala 33:92]
  wire [2:0] _dequeuedIndex_T_16 = readyVector[7] ? 3'h7 : 3'h0; // @[Mux.scala 101:16]
  wire [2:0] _dequeuedIndex_T_17 = readyVector[6] ? 3'h6 : _dequeuedIndex_T_16; // @[Mux.scala 101:16]
  wire [2:0] _dequeuedIndex_T_18 = readyVector[5] ? 3'h5 : _dequeuedIndex_T_17; // @[Mux.scala 101:16]
  wire [2:0] _dequeuedIndex_T_19 = readyVector[4] ? 3'h4 : _dequeuedIndex_T_18; // @[Mux.scala 101:16]
  wire [2:0] _dequeuedIndex_T_20 = readyVector[3] ? 3'h3 : _dequeuedIndex_T_19; // @[Mux.scala 101:16]
  wire [2:0] _dequeuedIndex_T_21 = readyVector[2] ? 3'h2 : _dequeuedIndex_T_20; // @[Mux.scala 101:16]
  wire [2:0] _dequeuedIndex_T_22 = readyVector[1] ? 3'h1 : _dequeuedIndex_T_21; // @[Mux.scala 101:16]
  wire [2:0] dequeuedIndex = readyVector[0] ? 3'h0 : _dequeuedIndex_T_22; // @[Mux.scala 101:16]
  wire  _dequeued_T_14_opcodeMeta_isM = readyVector[6] ? queue_6_opcodeMeta_isM : queue_7_opcodeMeta_isM; // @[Mux.scala 101:16]
  wire  _dequeued_T_14_valid = readyVector[6] ? queue_6_valid : queue_7_valid; // @[Mux.scala 101:16]
  wire [31:0] _dequeued_T_14_instruction = readyVector[6] ? queue_6_instruction : queue_7_instruction; // @[Mux.scala 101:16]
  wire [3:0] _dequeued_T_14_branchMask = readyVector[6] ? queue_6_branchMask : queue_7_branchMask; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_14_rs1_prfAddr = readyVector[6] ? queue_6_rs1_prfAddr : queue_7_rs1_prfAddr; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_14_rs2_prfAddr = readyVector[6] ? queue_6_rs2_prfAddr : queue_7_rs2_prfAddr; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_14_prfDest = readyVector[6] ? queue_6_prfDest : queue_7_prfDest; // @[Mux.scala 101:16]
  wire [3:0] _dequeued_T_14_robAddr = readyVector[6] ? queue_6_robAddr : queue_7_robAddr; // @[Mux.scala 101:16]
  wire  _dequeued_T_15_opcodeMeta_isM = readyVector[5] ? queue_5_opcodeMeta_isM : _dequeued_T_14_opcodeMeta_isM; // @[Mux.scala 101:16]
  wire  _dequeued_T_15_valid = readyVector[5] ? queue_5_valid : _dequeued_T_14_valid; // @[Mux.scala 101:16]
  wire [31:0] _dequeued_T_15_instruction = readyVector[5] ? queue_5_instruction : _dequeued_T_14_instruction; // @[Mux.scala 101:16]
  wire [3:0] _dequeued_T_15_branchMask = readyVector[5] ? queue_5_branchMask : _dequeued_T_14_branchMask; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_15_rs1_prfAddr = readyVector[5] ? queue_5_rs1_prfAddr : _dequeued_T_14_rs1_prfAddr; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_15_rs2_prfAddr = readyVector[5] ? queue_5_rs2_prfAddr : _dequeued_T_14_rs2_prfAddr; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_15_prfDest = readyVector[5] ? queue_5_prfDest : _dequeued_T_14_prfDest; // @[Mux.scala 101:16]
  wire [3:0] _dequeued_T_15_robAddr = readyVector[5] ? queue_5_robAddr : _dequeued_T_14_robAddr; // @[Mux.scala 101:16]
  wire  _dequeued_T_16_opcodeMeta_isM = readyVector[4] ? queue_4_opcodeMeta_isM : _dequeued_T_15_opcodeMeta_isM; // @[Mux.scala 101:16]
  wire  _dequeued_T_16_valid = readyVector[4] ? queue_4_valid : _dequeued_T_15_valid; // @[Mux.scala 101:16]
  wire [31:0] _dequeued_T_16_instruction = readyVector[4] ? queue_4_instruction : _dequeued_T_15_instruction; // @[Mux.scala 101:16]
  wire [3:0] _dequeued_T_16_branchMask = readyVector[4] ? queue_4_branchMask : _dequeued_T_15_branchMask; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_16_rs1_prfAddr = readyVector[4] ? queue_4_rs1_prfAddr : _dequeued_T_15_rs1_prfAddr; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_16_rs2_prfAddr = readyVector[4] ? queue_4_rs2_prfAddr : _dequeued_T_15_rs2_prfAddr; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_16_prfDest = readyVector[4] ? queue_4_prfDest : _dequeued_T_15_prfDest; // @[Mux.scala 101:16]
  wire [3:0] _dequeued_T_16_robAddr = readyVector[4] ? queue_4_robAddr : _dequeued_T_15_robAddr; // @[Mux.scala 101:16]
  wire  _dequeued_T_17_opcodeMeta_isM = readyVector[3] ? queue_3_opcodeMeta_isM : _dequeued_T_16_opcodeMeta_isM; // @[Mux.scala 101:16]
  wire  _dequeued_T_17_valid = readyVector[3] ? queue_3_valid : _dequeued_T_16_valid; // @[Mux.scala 101:16]
  wire [31:0] _dequeued_T_17_instruction = readyVector[3] ? queue_3_instruction : _dequeued_T_16_instruction; // @[Mux.scala 101:16]
  wire [3:0] _dequeued_T_17_branchMask = readyVector[3] ? queue_3_branchMask : _dequeued_T_16_branchMask; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_17_rs1_prfAddr = readyVector[3] ? queue_3_rs1_prfAddr : _dequeued_T_16_rs1_prfAddr; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_17_rs2_prfAddr = readyVector[3] ? queue_3_rs2_prfAddr : _dequeued_T_16_rs2_prfAddr; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_17_prfDest = readyVector[3] ? queue_3_prfDest : _dequeued_T_16_prfDest; // @[Mux.scala 101:16]
  wire [3:0] _dequeued_T_17_robAddr = readyVector[3] ? queue_3_robAddr : _dequeued_T_16_robAddr; // @[Mux.scala 101:16]
  wire  _dequeued_T_18_opcodeMeta_isM = readyVector[2] ? queue_2_opcodeMeta_isM : _dequeued_T_17_opcodeMeta_isM; // @[Mux.scala 101:16]
  wire  _dequeued_T_18_valid = readyVector[2] ? queue_2_valid : _dequeued_T_17_valid; // @[Mux.scala 101:16]
  wire [31:0] _dequeued_T_18_instruction = readyVector[2] ? queue_2_instruction : _dequeued_T_17_instruction; // @[Mux.scala 101:16]
  wire [3:0] _dequeued_T_18_branchMask = readyVector[2] ? queue_2_branchMask : _dequeued_T_17_branchMask; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_18_prfDest = readyVector[2] ? queue_2_prfDest : _dequeued_T_17_prfDest; // @[Mux.scala 101:16]
  wire  _dequeued_T_19_opcodeMeta_isM = readyVector[1] ? queue_1_opcodeMeta_isM : _dequeued_T_18_opcodeMeta_isM; // @[Mux.scala 101:16]
  wire  _dequeued_T_19_valid = readyVector[1] ? queue_1_valid : _dequeued_T_18_valid; // @[Mux.scala 101:16]
  wire [31:0] _dequeued_T_19_instruction = readyVector[1] ? queue_1_instruction : _dequeued_T_18_instruction; // @[Mux.scala 101:16]
  wire [3:0] _dequeued_T_19_branchMask = readyVector[1] ? queue_1_branchMask : _dequeued_T_18_branchMask; // @[Mux.scala 101:16]
  wire [5:0] _dequeued_T_19_prfDest = readyVector[1] ? queue_1_prfDest : _dequeued_T_18_prfDest; // @[Mux.scala 101:16]
  wire  dequeued_opcodeMeta_isM = readyVector[0] ? queue_0_opcodeMeta_isM : _dequeued_T_19_opcodeMeta_isM; // @[Mux.scala 101:16]
  wire  dequeued_valid = readyVector[0] ? queue_0_valid : _dequeued_T_19_valid; // @[Mux.scala 101:16]
  wire [31:0] dequeued_instruction = readyVector[0] ? queue_0_instruction : _dequeued_T_19_instruction; // @[Mux.scala 101:16]
  wire [3:0] dequeued_branchMask = readyVector[0] ? queue_0_branchMask : _dequeued_T_19_branchMask; // @[Mux.scala 101:16]
  wire [5:0] dequeued_prfDest = readyVector[0] ? queue_0_prfDest : _dequeued_T_19_prfDest; // @[Mux.scala 101:16]
  reg  releasedBuffer_valid; // @[scheduler.scala 59:31]
  reg [31:0] releasedBuffer_instruction; // @[scheduler.scala 59:31]
  reg [3:0] releasedBuffer_branchMask; // @[scheduler.scala 59:31]
  reg [5:0] releasedBuffer_rs1prfAddr; // @[scheduler.scala 59:31]
  reg [5:0] releasedBuffer_rs2prfAddr; // @[scheduler.scala 59:31]
  reg [5:0] releasedBuffer_prfDest; // @[scheduler.scala 59:31]
  reg [3:0] releasedBuffer_robAddr; // @[scheduler.scala 59:31]
  wire  dequeue = ~releasedBuffer_valid | release_fired; // @[scheduler.scala 70:39]
  wire [4:0] _tempQueue_8_opcodeMeta_meta_isM_T_1 = allocate_instruction[6:2] & 5'h1d; // @[scheduler.scala 78:44]
  wire  tempQueue_8_opcodeMeta_meta_isM = 5'hc == _tempQueue_8_opcodeMeta_meta_isM_T_1 & allocate_instruction[25]; // @[scheduler.scala 78:66]
  wire  tempQueue_8_opcodeMeta_meta_isMemAccess = ~allocate_instruction[6] & ~allocate_instruction[4] & ~(5'h3 ==
    allocate_instruction[6:2]); // @[scheduler.scala 79:92]
  wire  tempQueue_8_opcodeMeta_meta_isBranch = allocate_instruction[6:5] == 2'h3; // @[scheduler.scala 80:48]
  wire  tempQueue_8_rs2_ready = allocate_fired & tempQueue_8_opcodeMeta_meta_isMemAccess | allocate_rs2_ready; // @[scheduler.scala 89:116 86:34 89:77]
  wire [4:0] _wakeUpInt_valid_T_1 = dequeued_instruction[6:2] & 5'h15; // @[scheduler.scala 95:49]
  wire  _wakeUpInt_valid_T_6 = |readyVector; // @[scheduler.scala 95:125]
  wire  wakeUpInt_valid = 5'h4 == _wakeUpInt_valid_T_1 & ~dequeued_opcodeMeta_isM & dequeue & |readyVector & |
    dequeued_instruction[11:7]; // @[scheduler.scala 95:129]
  wire  updatedEntries_0_rs1_ready = queue_0_valid & (queue_0_rs1_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_0_rs1_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_0_rs1_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_0_rs1_prfAddr)); // @[scheduler.scala 98:109]
  wire  updatedEntries_1_rs1_ready = queue_1_valid & (queue_1_rs1_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_1_rs1_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_1_rs1_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_1_rs1_prfAddr)); // @[scheduler.scala 98:109]
  wire  updatedEntries_2_rs1_ready = queue_2_valid & (queue_2_rs1_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_2_rs1_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_2_rs1_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_2_rs1_prfAddr)); // @[scheduler.scala 98:109]
  wire  updatedEntries_3_rs1_ready = queue_3_valid & (queue_3_rs1_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_3_rs1_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_3_rs1_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_3_rs1_prfAddr)); // @[scheduler.scala 98:109]
  wire  updatedEntries_4_rs1_ready = queue_4_valid & (queue_4_rs1_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_4_rs1_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_4_rs1_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_4_rs1_prfAddr)); // @[scheduler.scala 98:109]
  wire  updatedEntries_5_rs1_ready = queue_5_valid & (queue_5_rs1_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_5_rs1_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_5_rs1_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_5_rs1_prfAddr)); // @[scheduler.scala 98:109]
  wire  updatedEntries_6_rs1_ready = queue_6_valid & (queue_6_rs1_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_6_rs1_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_6_rs1_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_6_rs1_prfAddr)); // @[scheduler.scala 98:109]
  wire  updatedEntries_7_rs1_ready = queue_7_valid & (queue_7_rs1_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_7_rs1_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_7_rs1_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_7_rs1_prfAddr)); // @[scheduler.scala 98:109]
  wire  updatedEntries_8_rs1_ready = allocate_fired & (allocate_rs1_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    allocate_rs1_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == allocate_rs1_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == allocate_rs1_prfAddr)); // @[scheduler.scala 98:109]
  reg  instrRetired_REG_valid; // @[scheduler.scala 101:26]
  reg [5:0] instrRetired_REG_prfAddr; // @[scheduler.scala 101:26]
  wire  updatedEntries_0_rs2_ready = queue_0_valid & (queue_0_rs2_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_0_rs2_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_0_rs2_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_0_rs2_prfAddr)); // @[scheduler.scala 104:42]
  wire  updatedEntries_1_rs2_ready = queue_1_valid & (queue_1_rs2_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_1_rs2_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_1_rs2_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_1_rs2_prfAddr)); // @[scheduler.scala 104:42]
  wire  updatedEntries_2_rs2_ready = queue_2_valid & (queue_2_rs2_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_2_rs2_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_2_rs2_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_2_rs2_prfAddr)); // @[scheduler.scala 104:42]
  wire  updatedEntries_3_rs2_ready = queue_3_valid & (queue_3_rs2_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_3_rs2_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_3_rs2_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_3_rs2_prfAddr)); // @[scheduler.scala 104:42]
  wire  updatedEntries_4_rs2_ready = queue_4_valid & (queue_4_rs2_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_4_rs2_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_4_rs2_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_4_rs2_prfAddr)); // @[scheduler.scala 104:42]
  wire  updatedEntries_5_rs2_ready = queue_5_valid & (queue_5_rs2_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_5_rs2_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_5_rs2_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_5_rs2_prfAddr)); // @[scheduler.scala 104:42]
  wire  updatedEntries_6_rs2_ready = queue_6_valid & (queue_6_rs2_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_6_rs2_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_6_rs2_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_6_rs2_prfAddr)); // @[scheduler.scala 104:42]
  wire  updatedEntries_7_rs2_ready = queue_7_valid & (queue_7_rs2_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr ==
    queue_7_rs2_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == queue_7_rs2_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == queue_7_rs2_prfAddr)); // @[scheduler.scala 104:42]
  wire  updatedEntries_8_rs2_ready = allocate_fired & (tempQueue_8_rs2_ready | (wakeUpExt_0_valid & wakeUpExt_0_prfAddr
     == allocate_rs2_prfAddr | wakeUpExt_1_valid & wakeUpExt_1_prfAddr == allocate_rs2_prfAddr | wakeUpInt_valid &
    dequeued_prfDest == allocate_rs2_prfAddr)); // @[scheduler.scala 104:42]
  wire [3:0] _T_1 = queue_0_branchMask & branchOps_branchMask; // @[scheduler.scala 109:53]
  wire  _T_2 = |_T_1; // @[scheduler.scala 109:77]
  wire [3:0] _updatedEntries_0_branchMask_T = queue_0_branchMask ^ branchOps_branchMask; // @[scheduler.scala 109:127]
  wire  _GEN_2 = branchOps_passed & |_T_1 ? queue_0_valid : queue_0_valid & ~_T_2; // @[scheduler.scala 109:82 110:35 92:81]
  wire  _GEN_4 = branchOps_valid ? _GEN_2 : queue_0_valid; // @[scheduler.scala 108:27 92:81]
  wire [3:0] _T_4 = queue_1_branchMask & branchOps_branchMask; // @[scheduler.scala 109:53]
  wire  _T_5 = |_T_4; // @[scheduler.scala 109:77]
  wire [3:0] _updatedEntries_1_branchMask_T = queue_1_branchMask ^ branchOps_branchMask; // @[scheduler.scala 109:127]
  wire  _GEN_6 = branchOps_passed & |_T_4 ? queue_1_valid : queue_1_valid & ~_T_5; // @[scheduler.scala 109:82 110:35 92:81]
  wire  _GEN_8 = branchOps_valid ? _GEN_6 : queue_1_valid; // @[scheduler.scala 108:27 92:81]
  wire [3:0] _T_7 = queue_2_branchMask & branchOps_branchMask; // @[scheduler.scala 109:53]
  wire  _T_8 = |_T_7; // @[scheduler.scala 109:77]
  wire [3:0] _updatedEntries_2_branchMask_T = queue_2_branchMask ^ branchOps_branchMask; // @[scheduler.scala 109:127]
  wire  _GEN_10 = branchOps_passed & |_T_7 ? queue_2_valid : queue_2_valid & ~_T_8; // @[scheduler.scala 109:82 110:35 92:81]
  wire  _GEN_12 = branchOps_valid ? _GEN_10 : queue_2_valid; // @[scheduler.scala 108:27 92:81]
  wire [3:0] _T_10 = queue_3_branchMask & branchOps_branchMask; // @[scheduler.scala 109:53]
  wire  _T_11 = |_T_10; // @[scheduler.scala 109:77]
  wire [3:0] _updatedEntries_3_branchMask_T = queue_3_branchMask ^ branchOps_branchMask; // @[scheduler.scala 109:127]
  wire  _GEN_14 = branchOps_passed & |_T_10 ? queue_3_valid : queue_3_valid & ~_T_11; // @[scheduler.scala 109:82 110:35 92:81]
  wire  _GEN_16 = branchOps_valid ? _GEN_14 : queue_3_valid; // @[scheduler.scala 108:27 92:81]
  wire [3:0] _T_13 = queue_4_branchMask & branchOps_branchMask; // @[scheduler.scala 109:53]
  wire  _T_14 = |_T_13; // @[scheduler.scala 109:77]
  wire [3:0] _updatedEntries_4_branchMask_T = queue_4_branchMask ^ branchOps_branchMask; // @[scheduler.scala 109:127]
  wire  _GEN_18 = branchOps_passed & |_T_13 ? queue_4_valid : queue_4_valid & ~_T_14; // @[scheduler.scala 109:82 110:35 92:81]
  wire  _GEN_20 = branchOps_valid ? _GEN_18 : queue_4_valid; // @[scheduler.scala 108:27 92:81]
  wire [3:0] _T_16 = queue_5_branchMask & branchOps_branchMask; // @[scheduler.scala 109:53]
  wire  _T_17 = |_T_16; // @[scheduler.scala 109:77]
  wire [3:0] _updatedEntries_5_branchMask_T = queue_5_branchMask ^ branchOps_branchMask; // @[scheduler.scala 109:127]
  wire  _GEN_22 = branchOps_passed & |_T_16 ? queue_5_valid : queue_5_valid & ~_T_17; // @[scheduler.scala 109:82 110:35 92:81]
  wire  _GEN_24 = branchOps_valid ? _GEN_22 : queue_5_valid; // @[scheduler.scala 108:27 92:81]
  wire [3:0] _T_19 = queue_6_branchMask & branchOps_branchMask; // @[scheduler.scala 109:53]
  wire  _T_20 = |_T_19; // @[scheduler.scala 109:77]
  wire [3:0] _updatedEntries_6_branchMask_T = queue_6_branchMask ^ branchOps_branchMask; // @[scheduler.scala 109:127]
  wire  _GEN_26 = branchOps_passed & |_T_19 ? queue_6_valid : queue_6_valid & ~_T_20; // @[scheduler.scala 109:82 110:35 92:81]
  wire  _GEN_28 = branchOps_valid ? _GEN_26 : queue_6_valid; // @[scheduler.scala 108:27 92:81]
  wire [3:0] _T_22 = queue_7_branchMask & branchOps_branchMask; // @[scheduler.scala 109:53]
  wire  _T_23 = |_T_22; // @[scheduler.scala 109:77]
  wire [3:0] _updatedEntries_7_branchMask_T = queue_7_branchMask ^ branchOps_branchMask; // @[scheduler.scala 109:127]
  wire  _GEN_30 = branchOps_passed & |_T_22 ? queue_7_valid : queue_7_valid & ~_T_23; // @[scheduler.scala 109:82 110:35 92:81]
  wire  _GEN_32 = branchOps_valid ? _GEN_30 : queue_7_valid; // @[scheduler.scala 108:27 92:81]
  wire [3:0] _T_25 = allocate_branchMask & branchOps_branchMask; // @[scheduler.scala 109:53]
  wire  _T_26 = |_T_25; // @[scheduler.scala 109:77]
  wire [3:0] _updatedEntries_8_branchMask_T = allocate_branchMask ^ branchOps_branchMask; // @[scheduler.scala 109:127]
  wire  _T_29 = dequeue & _wakeUpInt_valid_T_6; // @[scheduler.scala 114:16]
  wire  _newQueue_T_69 = queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid
     & queue_6_valid & queue_7_valid; // @[scheduler.scala 116:110]
  wire [3:0] _releasedBuffer_branchMask_T = branchOps_branchMask & dequeued_branchMask; // @[scheduler.scala 137:79]
  wire [3:0] _releasedBuffer_branchMask_T_4 = dequeued_branchMask ^ branchOps_branchMask; // @[scheduler.scala 137:147]
  wire  _releasedBuffer_valid_T = ~branchOps_valid; // @[scheduler.scala 143:48]
  wire [3:0] _releasedBuffer_valid_T_1 = dequeued_branchMask & branchOps_branchMask; // @[scheduler.scala 143:90]
  wire [3:0] _releasedBuffer_branchMask_T_6 = releasedBuffer_branchMask ^ branchOps_branchMask; // @[scheduler.scala 145:60]
  wire [3:0] _releasedBuffer_valid_T_10 = releasedBuffer_branchMask & branchOps_branchMask; // @[scheduler.scala 146:102]
  assign allocate_ready = ~_newQueue_T_69; // @[scheduler.scala 134:21]
  assign release_ready = releasedBuffer_valid; // @[scheduler.scala 133:17]
  assign release_instruction = releasedBuffer_instruction; // @[scheduler.scala 128:23]
  assign release_branchMask = releasedBuffer_branchMask; // @[scheduler.scala 127:22]
  assign release_rs1prfAddr = releasedBuffer_rs1prfAddr; // @[scheduler.scala 131:22]
  assign release_rs2prfAddr = releasedBuffer_rs2prfAddr; // @[scheduler.scala 132:22]
  assign release_prfDest = releasedBuffer_prfDest; // @[scheduler.scala 129:19]
  assign release_robAddr = releasedBuffer_robAddr; // @[scheduler.scala 130:19]
  assign instrRetired_valid = instrRetired_REG_valid; // @[scheduler.scala 101:16]
  assign instrRetired_prfAddr = instrRetired_REG_prfAddr; // @[scheduler.scala 101:16]
  always @(posedge clock) begin
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_opcodeMeta_isBranch <= queue_1_opcodeMeta_isBranch;
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_opcodeMeta_isMemAccess <= queue_1_opcodeMeta_isMemAccess;
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_opcodeMeta_isM <= queue_1_opcodeMeta_isM;
    end
    if (reset) begin // @[scheduler.scala 26:22]
      queue_0_valid <= 1'h0; // @[scheduler.scala 26:22]
    end else if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
        if (3'h1 == dequeuedIndex) begin // @[scheduler.scala 114:106]
          queue_0_valid <= 1'h0; // @[scheduler.scala 114:132]
        end else begin
          queue_0_valid <= _GEN_8;
        end
      end else begin
        queue_0_valid <= _GEN_8;
      end
    end else if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
      if (3'h0 == dequeuedIndex) begin // @[scheduler.scala 114:106]
        queue_0_valid <= 1'h0; // @[scheduler.scala 114:132]
      end else begin
        queue_0_valid <= _GEN_4;
      end
    end else begin
      queue_0_valid <= _GEN_4;
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_instruction <= queue_1_instruction;
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      if (branchOps_valid) begin // @[scheduler.scala 108:27]
        if (branchOps_passed & |_T_4) begin // @[scheduler.scala 109:82]
          queue_0_branchMask <= _updatedEntries_1_branchMask_T; // @[scheduler.scala 109:104]
        end else begin
          queue_0_branchMask <= queue_1_branchMask; // @[scheduler.scala 92:81]
        end
      end else begin
        queue_0_branchMask <= queue_1_branchMask; // @[scheduler.scala 92:81]
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 108:27]
      if (branchOps_passed & |_T_1) begin // @[scheduler.scala 109:82]
        queue_0_branchMask <= _updatedEntries_0_branchMask_T; // @[scheduler.scala 109:104]
      end
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_rs1_ready <= updatedEntries_1_rs1_ready;
    end else begin
      queue_0_rs1_ready <= updatedEntries_0_rs1_ready;
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_rs1_prfAddr <= queue_1_rs1_prfAddr;
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_rs2_ready <= updatedEntries_1_rs2_ready;
    end else begin
      queue_0_rs2_ready <= updatedEntries_0_rs2_ready;
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_rs2_prfAddr <= queue_1_rs2_prfAddr;
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_prfDest <= queue_1_prfDest;
    end
    if (~queue_0_valid | dequeue & |readyVector[0]) begin // @[scheduler.scala 116:60]
      queue_0_robAddr <= queue_1_robAddr;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_opcodeMeta_isBranch <= queue_2_opcodeMeta_isBranch;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_opcodeMeta_isMemAccess <= queue_2_opcodeMeta_isMemAccess;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_opcodeMeta_isM <= queue_2_opcodeMeta_isM;
    end
    if (reset) begin // @[scheduler.scala 26:22]
      queue_1_valid <= 1'h0; // @[scheduler.scala 26:22]
    end else if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
        if (3'h2 == dequeuedIndex) begin // @[scheduler.scala 114:106]
          queue_1_valid <= 1'h0; // @[scheduler.scala 114:132]
        end else begin
          queue_1_valid <= _GEN_12;
        end
      end else begin
        queue_1_valid <= _GEN_12;
      end
    end else if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
      if (3'h1 == dequeuedIndex) begin // @[scheduler.scala 114:106]
        queue_1_valid <= 1'h0; // @[scheduler.scala 114:132]
      end else begin
        queue_1_valid <= _GEN_8;
      end
    end else begin
      queue_1_valid <= _GEN_8;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_instruction <= queue_2_instruction;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      if (branchOps_valid) begin // @[scheduler.scala 108:27]
        if (branchOps_passed & |_T_7) begin // @[scheduler.scala 109:82]
          queue_1_branchMask <= _updatedEntries_2_branchMask_T; // @[scheduler.scala 109:104]
        end else begin
          queue_1_branchMask <= queue_2_branchMask; // @[scheduler.scala 92:81]
        end
      end else begin
        queue_1_branchMask <= queue_2_branchMask; // @[scheduler.scala 92:81]
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 108:27]
      if (branchOps_passed & |_T_4) begin // @[scheduler.scala 109:82]
        queue_1_branchMask <= _updatedEntries_1_branchMask_T; // @[scheduler.scala 109:104]
      end
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_rs1_ready <= updatedEntries_2_rs1_ready;
    end else begin
      queue_1_rs1_ready <= updatedEntries_1_rs1_ready;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_rs1_prfAddr <= queue_2_rs1_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_rs2_ready <= updatedEntries_2_rs2_ready;
    end else begin
      queue_1_rs2_ready <= updatedEntries_1_rs2_ready;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_rs2_prfAddr <= queue_2_rs2_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_prfDest <= queue_2_prfDest;
    end
    if (~(queue_0_valid & queue_1_valid) | dequeue & |readyVector[1:0]) begin // @[scheduler.scala 116:60]
      queue_1_robAddr <= queue_2_robAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_opcodeMeta_isBranch <= queue_3_opcodeMeta_isBranch;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_opcodeMeta_isMemAccess <= queue_3_opcodeMeta_isMemAccess;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_opcodeMeta_isM <= queue_3_opcodeMeta_isM;
    end
    if (reset) begin // @[scheduler.scala 26:22]
      queue_2_valid <= 1'h0; // @[scheduler.scala 26:22]
    end else if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
        if (3'h3 == dequeuedIndex) begin // @[scheduler.scala 114:106]
          queue_2_valid <= 1'h0; // @[scheduler.scala 114:132]
        end else begin
          queue_2_valid <= _GEN_16;
        end
      end else begin
        queue_2_valid <= _GEN_16;
      end
    end else if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
      if (3'h2 == dequeuedIndex) begin // @[scheduler.scala 114:106]
        queue_2_valid <= 1'h0; // @[scheduler.scala 114:132]
      end else begin
        queue_2_valid <= _GEN_12;
      end
    end else begin
      queue_2_valid <= _GEN_12;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_instruction <= queue_3_instruction;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      if (branchOps_valid) begin // @[scheduler.scala 108:27]
        if (branchOps_passed & |_T_10) begin // @[scheduler.scala 109:82]
          queue_2_branchMask <= _updatedEntries_3_branchMask_T; // @[scheduler.scala 109:104]
        end else begin
          queue_2_branchMask <= queue_3_branchMask; // @[scheduler.scala 92:81]
        end
      end else begin
        queue_2_branchMask <= queue_3_branchMask; // @[scheduler.scala 92:81]
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 108:27]
      if (branchOps_passed & |_T_7) begin // @[scheduler.scala 109:82]
        queue_2_branchMask <= _updatedEntries_2_branchMask_T; // @[scheduler.scala 109:104]
      end
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_rs1_ready <= updatedEntries_3_rs1_ready;
    end else begin
      queue_2_rs1_ready <= updatedEntries_2_rs1_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_rs1_prfAddr <= queue_3_rs1_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_rs2_ready <= updatedEntries_3_rs2_ready;
    end else begin
      queue_2_rs2_ready <= updatedEntries_2_rs2_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_rs2_prfAddr <= queue_3_rs2_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_prfDest <= queue_3_prfDest;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid) | dequeue & |readyVector[2:0]) begin // @[scheduler.scala 116:60]
      queue_2_robAddr <= queue_3_robAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_opcodeMeta_isBranch <= queue_4_opcodeMeta_isBranch;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_opcodeMeta_isMemAccess <= queue_4_opcodeMeta_isMemAccess;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_opcodeMeta_isM <= queue_4_opcodeMeta_isM;
    end
    if (reset) begin // @[scheduler.scala 26:22]
      queue_3_valid <= 1'h0; // @[scheduler.scala 26:22]
    end else if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
        if (3'h4 == dequeuedIndex) begin // @[scheduler.scala 114:106]
          queue_3_valid <= 1'h0; // @[scheduler.scala 114:132]
        end else begin
          queue_3_valid <= _GEN_20;
        end
      end else begin
        queue_3_valid <= _GEN_20;
      end
    end else if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
      if (3'h3 == dequeuedIndex) begin // @[scheduler.scala 114:106]
        queue_3_valid <= 1'h0; // @[scheduler.scala 114:132]
      end else begin
        queue_3_valid <= _GEN_16;
      end
    end else begin
      queue_3_valid <= _GEN_16;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_instruction <= queue_4_instruction;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      if (branchOps_valid) begin // @[scheduler.scala 108:27]
        if (branchOps_passed & |_T_13) begin // @[scheduler.scala 109:82]
          queue_3_branchMask <= _updatedEntries_4_branchMask_T; // @[scheduler.scala 109:104]
        end else begin
          queue_3_branchMask <= queue_4_branchMask; // @[scheduler.scala 92:81]
        end
      end else begin
        queue_3_branchMask <= queue_4_branchMask; // @[scheduler.scala 92:81]
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 108:27]
      if (branchOps_passed & |_T_10) begin // @[scheduler.scala 109:82]
        queue_3_branchMask <= _updatedEntries_3_branchMask_T; // @[scheduler.scala 109:104]
      end
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_rs1_ready <= updatedEntries_4_rs1_ready;
    end else begin
      queue_3_rs1_ready <= updatedEntries_3_rs1_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_rs1_prfAddr <= queue_4_rs1_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_rs2_ready <= updatedEntries_4_rs2_ready;
    end else begin
      queue_3_rs2_ready <= updatedEntries_3_rs2_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_rs2_prfAddr <= queue_4_rs2_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_prfDest <= queue_4_prfDest;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid) | dequeue & |readyVector[3:0]) begin // @[scheduler.scala 116:60]
      queue_3_robAddr <= queue_4_robAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_opcodeMeta_isBranch <= queue_5_opcodeMeta_isBranch;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_opcodeMeta_isMemAccess <= queue_5_opcodeMeta_isMemAccess;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_opcodeMeta_isM <= queue_5_opcodeMeta_isM;
    end
    if (reset) begin // @[scheduler.scala 26:22]
      queue_4_valid <= 1'h0; // @[scheduler.scala 26:22]
    end else if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |
      readyVector[4:0]) begin // @[scheduler.scala 116:60]
      if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
        if (3'h5 == dequeuedIndex) begin // @[scheduler.scala 114:106]
          queue_4_valid <= 1'h0; // @[scheduler.scala 114:132]
        end else begin
          queue_4_valid <= _GEN_24;
        end
      end else begin
        queue_4_valid <= _GEN_24;
      end
    end else if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
      if (3'h4 == dequeuedIndex) begin // @[scheduler.scala 114:106]
        queue_4_valid <= 1'h0; // @[scheduler.scala 114:132]
      end else begin
        queue_4_valid <= _GEN_20;
      end
    end else begin
      queue_4_valid <= _GEN_20;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_instruction <= queue_5_instruction;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      if (branchOps_valid) begin // @[scheduler.scala 108:27]
        if (branchOps_passed & |_T_16) begin // @[scheduler.scala 109:82]
          queue_4_branchMask <= _updatedEntries_5_branchMask_T; // @[scheduler.scala 109:104]
        end else begin
          queue_4_branchMask <= queue_5_branchMask; // @[scheduler.scala 92:81]
        end
      end else begin
        queue_4_branchMask <= queue_5_branchMask; // @[scheduler.scala 92:81]
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 108:27]
      if (branchOps_passed & |_T_13) begin // @[scheduler.scala 109:82]
        queue_4_branchMask <= _updatedEntries_4_branchMask_T; // @[scheduler.scala 109:104]
      end
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_rs1_ready <= updatedEntries_5_rs1_ready;
    end else begin
      queue_4_rs1_ready <= updatedEntries_4_rs1_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_rs1_prfAddr <= queue_5_rs1_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_rs2_ready <= updatedEntries_5_rs2_ready;
    end else begin
      queue_4_rs2_ready <= updatedEntries_4_rs2_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_rs2_prfAddr <= queue_5_rs2_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_prfDest <= queue_5_prfDest;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid) | dequeue & |readyVector[4:0]
      ) begin // @[scheduler.scala 116:60]
      queue_4_robAddr <= queue_5_robAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_opcodeMeta_isBranch <= queue_6_opcodeMeta_isBranch;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_opcodeMeta_isMemAccess <= queue_6_opcodeMeta_isMemAccess;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_opcodeMeta_isM <= queue_6_opcodeMeta_isM;
    end
    if (reset) begin // @[scheduler.scala 26:22]
      queue_5_valid <= 1'h0; // @[scheduler.scala 26:22]
    end else if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) |
      dequeue & |readyVector[5:0]) begin // @[scheduler.scala 116:60]
      if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
        if (3'h6 == dequeuedIndex) begin // @[scheduler.scala 114:106]
          queue_5_valid <= 1'h0; // @[scheduler.scala 114:132]
        end else begin
          queue_5_valid <= _GEN_28;
        end
      end else begin
        queue_5_valid <= _GEN_28;
      end
    end else if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
      if (3'h5 == dequeuedIndex) begin // @[scheduler.scala 114:106]
        queue_5_valid <= 1'h0; // @[scheduler.scala 114:132]
      end else begin
        queue_5_valid <= _GEN_24;
      end
    end else begin
      queue_5_valid <= _GEN_24;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_instruction <= queue_6_instruction;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      if (branchOps_valid) begin // @[scheduler.scala 108:27]
        if (branchOps_passed & |_T_19) begin // @[scheduler.scala 109:82]
          queue_5_branchMask <= _updatedEntries_6_branchMask_T; // @[scheduler.scala 109:104]
        end else begin
          queue_5_branchMask <= queue_6_branchMask; // @[scheduler.scala 92:81]
        end
      end else begin
        queue_5_branchMask <= queue_6_branchMask; // @[scheduler.scala 92:81]
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 108:27]
      if (branchOps_passed & |_T_16) begin // @[scheduler.scala 109:82]
        queue_5_branchMask <= _updatedEntries_5_branchMask_T; // @[scheduler.scala 109:104]
      end
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_rs1_ready <= updatedEntries_6_rs1_ready;
    end else begin
      queue_5_rs1_ready <= updatedEntries_5_rs1_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_rs1_prfAddr <= queue_6_rs1_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_rs2_ready <= updatedEntries_6_rs2_ready;
    end else begin
      queue_5_rs2_ready <= updatedEntries_5_rs2_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_rs2_prfAddr <= queue_6_rs2_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_prfDest <= queue_6_prfDest;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid) | dequeue & |
      readyVector[5:0]) begin // @[scheduler.scala 116:60]
      queue_5_robAddr <= queue_6_robAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_opcodeMeta_isBranch <= queue_7_opcodeMeta_isBranch;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_opcodeMeta_isMemAccess <= queue_7_opcodeMeta_isMemAccess;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_opcodeMeta_isM <= queue_7_opcodeMeta_isM;
    end
    if (reset) begin // @[scheduler.scala 26:22]
      queue_6_valid <= 1'h0; // @[scheduler.scala 26:22]
    end else if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid &
      queue_6_valid) | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
        if (3'h7 == dequeuedIndex) begin // @[scheduler.scala 114:106]
          queue_6_valid <= 1'h0; // @[scheduler.scala 114:132]
        end else begin
          queue_6_valid <= _GEN_32;
        end
      end else begin
        queue_6_valid <= _GEN_32;
      end
    end else if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
      if (3'h6 == dequeuedIndex) begin // @[scheduler.scala 114:106]
        queue_6_valid <= 1'h0; // @[scheduler.scala 114:132]
      end else begin
        queue_6_valid <= _GEN_28;
      end
    end else begin
      queue_6_valid <= _GEN_28;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_instruction <= queue_7_instruction;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      if (branchOps_valid) begin // @[scheduler.scala 108:27]
        if (branchOps_passed & |_T_22) begin // @[scheduler.scala 109:82]
          queue_6_branchMask <= _updatedEntries_7_branchMask_T; // @[scheduler.scala 109:104]
        end else begin
          queue_6_branchMask <= queue_7_branchMask; // @[scheduler.scala 92:81]
        end
      end else begin
        queue_6_branchMask <= queue_7_branchMask; // @[scheduler.scala 92:81]
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 108:27]
      if (branchOps_passed & |_T_19) begin // @[scheduler.scala 109:82]
        queue_6_branchMask <= _updatedEntries_6_branchMask_T; // @[scheduler.scala 109:104]
      end
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_rs1_ready <= updatedEntries_7_rs1_ready;
    end else begin
      queue_6_rs1_ready <= updatedEntries_6_rs1_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_rs1_prfAddr <= queue_7_rs1_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_rs2_ready <= updatedEntries_7_rs2_ready;
    end else begin
      queue_6_rs2_ready <= updatedEntries_6_rs2_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_rs2_prfAddr <= queue_7_rs2_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_prfDest <= queue_7_prfDest;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid)
       | dequeue & |readyVector[6:0]) begin // @[scheduler.scala 116:60]
      queue_6_robAddr <= queue_7_robAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_opcodeMeta_isBranch <= tempQueue_8_opcodeMeta_meta_isBranch;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_opcodeMeta_isMemAccess <= tempQueue_8_opcodeMeta_meta_isMemAccess;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_opcodeMeta_isM <= tempQueue_8_opcodeMeta_meta_isM;
    end
    if (reset) begin // @[scheduler.scala 26:22]
      queue_7_valid <= 1'h0; // @[scheduler.scala 26:22]
    end else if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid &
      queue_6_valid & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      if (branchOps_valid) begin // @[scheduler.scala 108:27]
        if (branchOps_passed & |_T_25) begin // @[scheduler.scala 109:82]
          queue_7_valid <= allocate_fired; // @[scheduler.scala 92:81]
        end else begin
          queue_7_valid <= allocate_fired & ~_T_26; // @[scheduler.scala 110:35]
        end
      end else begin
        queue_7_valid <= allocate_fired; // @[scheduler.scala 92:81]
      end
    end else if (dequeue & _wakeUpInt_valid_T_6) begin // @[scheduler.scala 114:36]
      if (3'h7 == dequeuedIndex) begin // @[scheduler.scala 114:106]
        queue_7_valid <= 1'h0; // @[scheduler.scala 114:132]
      end else begin
        queue_7_valid <= _GEN_32;
      end
    end else begin
      queue_7_valid <= _GEN_32;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_instruction <= allocate_instruction;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      if (branchOps_valid) begin // @[scheduler.scala 108:27]
        if (branchOps_passed & |_T_25) begin // @[scheduler.scala 109:82]
          queue_7_branchMask <= _updatedEntries_8_branchMask_T; // @[scheduler.scala 109:104]
        end else begin
          queue_7_branchMask <= allocate_branchMask; // @[scheduler.scala 92:81]
        end
      end else begin
        queue_7_branchMask <= allocate_branchMask; // @[scheduler.scala 92:81]
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 108:27]
      if (branchOps_passed & |_T_22) begin // @[scheduler.scala 109:82]
        queue_7_branchMask <= _updatedEntries_7_branchMask_T; // @[scheduler.scala 109:104]
      end
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_rs1_ready <= updatedEntries_8_rs1_ready;
    end else begin
      queue_7_rs1_ready <= updatedEntries_7_rs1_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_rs1_prfAddr <= allocate_rs1_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_rs2_ready <= updatedEntries_8_rs2_ready;
    end else begin
      queue_7_rs2_ready <= updatedEntries_7_rs2_ready;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_rs2_prfAddr <= allocate_rs2_prfAddr;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_prfDest <= allocate_prfDest;
    end
    if (~(queue_0_valid & queue_1_valid & queue_2_valid & queue_3_valid & queue_4_valid & queue_5_valid & queue_6_valid
       & queue_7_valid) | _T_29) begin // @[scheduler.scala 116:60]
      queue_7_robAddr <= allocate_robAddr;
    end
    if (reset) begin // @[scheduler.scala 59:31]
      releasedBuffer_valid <= 1'h0; // @[scheduler.scala 59:31]
    end else if (dequeue) begin // @[scheduler.scala 136:17]
      releasedBuffer_valid <= dequeued_valid & (~branchOps_valid | ~(|_releasedBuffer_valid_T_1) | branchOps_passed) &
        _wakeUpInt_valid_T_6; // @[scheduler.scala 143:26]
    end else if (branchOps_valid) begin // @[scheduler.scala 144:31]
      releasedBuffer_valid <= releasedBuffer_valid & (_releasedBuffer_valid_T | ~(|_releasedBuffer_valid_T_10) |
        branchOps_passed); // @[scheduler.scala 146:26]
    end
    if (dequeue) begin // @[scheduler.scala 136:17]
      if (readyVector[0]) begin // @[Mux.scala 101:16]
        releasedBuffer_instruction <= queue_0_instruction;
      end else if (readyVector[1]) begin // @[Mux.scala 101:16]
        releasedBuffer_instruction <= queue_1_instruction;
      end else if (readyVector[2]) begin // @[Mux.scala 101:16]
        releasedBuffer_instruction <= queue_2_instruction;
      end else begin
        releasedBuffer_instruction <= _dequeued_T_17_instruction;
      end
    end
    if (dequeue) begin // @[scheduler.scala 136:17]
      if (branchOps_valid & |_releasedBuffer_branchMask_T & branchOps_passed) begin // @[scheduler.scala 137:37]
        releasedBuffer_branchMask <= _releasedBuffer_branchMask_T_4;
      end else if (readyVector[0]) begin // @[Mux.scala 101:16]
        releasedBuffer_branchMask <= queue_0_branchMask;
      end else if (readyVector[1]) begin // @[Mux.scala 101:16]
        releasedBuffer_branchMask <= queue_1_branchMask;
      end else begin
        releasedBuffer_branchMask <= _dequeued_T_18_branchMask;
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 144:31]
      releasedBuffer_branchMask <= _releasedBuffer_branchMask_T_6; // @[scheduler.scala 145:31]
    end
    if (dequeue) begin // @[scheduler.scala 136:17]
      if (readyVector[0]) begin // @[Mux.scala 101:16]
        releasedBuffer_rs1prfAddr <= queue_0_rs1_prfAddr;
      end else if (readyVector[1]) begin // @[Mux.scala 101:16]
        releasedBuffer_rs1prfAddr <= queue_1_rs1_prfAddr;
      end else if (readyVector[2]) begin // @[Mux.scala 101:16]
        releasedBuffer_rs1prfAddr <= queue_2_rs1_prfAddr;
      end else begin
        releasedBuffer_rs1prfAddr <= _dequeued_T_17_rs1_prfAddr;
      end
    end
    if (dequeue) begin // @[scheduler.scala 136:17]
      if (readyVector[0]) begin // @[Mux.scala 101:16]
        releasedBuffer_rs2prfAddr <= queue_0_rs2_prfAddr;
      end else if (readyVector[1]) begin // @[Mux.scala 101:16]
        releasedBuffer_rs2prfAddr <= queue_1_rs2_prfAddr;
      end else if (readyVector[2]) begin // @[Mux.scala 101:16]
        releasedBuffer_rs2prfAddr <= queue_2_rs2_prfAddr;
      end else begin
        releasedBuffer_rs2prfAddr <= _dequeued_T_17_rs2_prfAddr;
      end
    end
    if (dequeue) begin // @[scheduler.scala 136:17]
      if (readyVector[0]) begin // @[Mux.scala 101:16]
        releasedBuffer_prfDest <= queue_0_prfDest;
      end else if (readyVector[1]) begin // @[Mux.scala 101:16]
        releasedBuffer_prfDest <= queue_1_prfDest;
      end else if (readyVector[2]) begin // @[Mux.scala 101:16]
        releasedBuffer_prfDest <= queue_2_prfDest;
      end else begin
        releasedBuffer_prfDest <= _dequeued_T_17_prfDest;
      end
    end
    if (dequeue) begin // @[scheduler.scala 136:17]
      if (readyVector[0]) begin // @[Mux.scala 101:16]
        releasedBuffer_robAddr <= queue_0_robAddr;
      end else if (readyVector[1]) begin // @[Mux.scala 101:16]
        releasedBuffer_robAddr <= queue_1_robAddr;
      end else if (readyVector[2]) begin // @[Mux.scala 101:16]
        releasedBuffer_robAddr <= queue_2_robAddr;
      end else begin
        releasedBuffer_robAddr <= _dequeued_T_17_robAddr;
      end
    end
    instrRetired_REG_valid <= 5'h4 == _wakeUpInt_valid_T_1 & ~dequeued_opcodeMeta_isM & dequeue & |readyVector & |
      dequeued_instruction[11:7]; // @[scheduler.scala 95:129]
    if (readyVector[0]) begin // @[Mux.scala 101:16]
      instrRetired_REG_prfAddr <= queue_0_prfDest;
    end else if (readyVector[1]) begin // @[Mux.scala 101:16]
      instrRetired_REG_prfAddr <= queue_1_prfDest;
    end else if (readyVector[2]) begin // @[Mux.scala 101:16]
      instrRetired_REG_prfAddr <= queue_2_prfDest;
    end else if (readyVector[3]) begin // @[Mux.scala 101:16]
      instrRetired_REG_prfAddr <= queue_3_prfDest;
    end else begin
      instrRetired_REG_prfAddr <= _dequeued_T_16_prfDest;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  queue_0_opcodeMeta_isBranch = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  queue_0_opcodeMeta_isMemAccess = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  queue_0_opcodeMeta_isM = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  queue_0_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  queue_0_instruction = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  queue_0_branchMask = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  queue_0_rs1_ready = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  queue_0_rs1_prfAddr = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  queue_0_rs2_ready = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  queue_0_rs2_prfAddr = _RAND_9[5:0];
  _RAND_10 = {1{`RANDOM}};
  queue_0_prfDest = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  queue_0_robAddr = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  queue_1_opcodeMeta_isBranch = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  queue_1_opcodeMeta_isMemAccess = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  queue_1_opcodeMeta_isM = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  queue_1_valid = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  queue_1_instruction = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  queue_1_branchMask = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  queue_1_rs1_ready = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  queue_1_rs1_prfAddr = _RAND_19[5:0];
  _RAND_20 = {1{`RANDOM}};
  queue_1_rs2_ready = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  queue_1_rs2_prfAddr = _RAND_21[5:0];
  _RAND_22 = {1{`RANDOM}};
  queue_1_prfDest = _RAND_22[5:0];
  _RAND_23 = {1{`RANDOM}};
  queue_1_robAddr = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  queue_2_opcodeMeta_isBranch = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  queue_2_opcodeMeta_isMemAccess = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  queue_2_opcodeMeta_isM = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  queue_2_valid = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  queue_2_instruction = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  queue_2_branchMask = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  queue_2_rs1_ready = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  queue_2_rs1_prfAddr = _RAND_31[5:0];
  _RAND_32 = {1{`RANDOM}};
  queue_2_rs2_ready = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  queue_2_rs2_prfAddr = _RAND_33[5:0];
  _RAND_34 = {1{`RANDOM}};
  queue_2_prfDest = _RAND_34[5:0];
  _RAND_35 = {1{`RANDOM}};
  queue_2_robAddr = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  queue_3_opcodeMeta_isBranch = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  queue_3_opcodeMeta_isMemAccess = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  queue_3_opcodeMeta_isM = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  queue_3_valid = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  queue_3_instruction = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  queue_3_branchMask = _RAND_41[3:0];
  _RAND_42 = {1{`RANDOM}};
  queue_3_rs1_ready = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  queue_3_rs1_prfAddr = _RAND_43[5:0];
  _RAND_44 = {1{`RANDOM}};
  queue_3_rs2_ready = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  queue_3_rs2_prfAddr = _RAND_45[5:0];
  _RAND_46 = {1{`RANDOM}};
  queue_3_prfDest = _RAND_46[5:0];
  _RAND_47 = {1{`RANDOM}};
  queue_3_robAddr = _RAND_47[3:0];
  _RAND_48 = {1{`RANDOM}};
  queue_4_opcodeMeta_isBranch = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  queue_4_opcodeMeta_isMemAccess = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  queue_4_opcodeMeta_isM = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  queue_4_valid = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  queue_4_instruction = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  queue_4_branchMask = _RAND_53[3:0];
  _RAND_54 = {1{`RANDOM}};
  queue_4_rs1_ready = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  queue_4_rs1_prfAddr = _RAND_55[5:0];
  _RAND_56 = {1{`RANDOM}};
  queue_4_rs2_ready = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  queue_4_rs2_prfAddr = _RAND_57[5:0];
  _RAND_58 = {1{`RANDOM}};
  queue_4_prfDest = _RAND_58[5:0];
  _RAND_59 = {1{`RANDOM}};
  queue_4_robAddr = _RAND_59[3:0];
  _RAND_60 = {1{`RANDOM}};
  queue_5_opcodeMeta_isBranch = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  queue_5_opcodeMeta_isMemAccess = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  queue_5_opcodeMeta_isM = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  queue_5_valid = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  queue_5_instruction = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  queue_5_branchMask = _RAND_65[3:0];
  _RAND_66 = {1{`RANDOM}};
  queue_5_rs1_ready = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  queue_5_rs1_prfAddr = _RAND_67[5:0];
  _RAND_68 = {1{`RANDOM}};
  queue_5_rs2_ready = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  queue_5_rs2_prfAddr = _RAND_69[5:0];
  _RAND_70 = {1{`RANDOM}};
  queue_5_prfDest = _RAND_70[5:0];
  _RAND_71 = {1{`RANDOM}};
  queue_5_robAddr = _RAND_71[3:0];
  _RAND_72 = {1{`RANDOM}};
  queue_6_opcodeMeta_isBranch = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  queue_6_opcodeMeta_isMemAccess = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  queue_6_opcodeMeta_isM = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  queue_6_valid = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  queue_6_instruction = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  queue_6_branchMask = _RAND_77[3:0];
  _RAND_78 = {1{`RANDOM}};
  queue_6_rs1_ready = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  queue_6_rs1_prfAddr = _RAND_79[5:0];
  _RAND_80 = {1{`RANDOM}};
  queue_6_rs2_ready = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  queue_6_rs2_prfAddr = _RAND_81[5:0];
  _RAND_82 = {1{`RANDOM}};
  queue_6_prfDest = _RAND_82[5:0];
  _RAND_83 = {1{`RANDOM}};
  queue_6_robAddr = _RAND_83[3:0];
  _RAND_84 = {1{`RANDOM}};
  queue_7_opcodeMeta_isBranch = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  queue_7_opcodeMeta_isMemAccess = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  queue_7_opcodeMeta_isM = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  queue_7_valid = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  queue_7_instruction = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  queue_7_branchMask = _RAND_89[3:0];
  _RAND_90 = {1{`RANDOM}};
  queue_7_rs1_ready = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  queue_7_rs1_prfAddr = _RAND_91[5:0];
  _RAND_92 = {1{`RANDOM}};
  queue_7_rs2_ready = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  queue_7_rs2_prfAddr = _RAND_93[5:0];
  _RAND_94 = {1{`RANDOM}};
  queue_7_prfDest = _RAND_94[5:0];
  _RAND_95 = {1{`RANDOM}};
  queue_7_robAddr = _RAND_95[3:0];
  _RAND_96 = {1{`RANDOM}};
  releasedBuffer_valid = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  releasedBuffer_instruction = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  releasedBuffer_branchMask = _RAND_98[3:0];
  _RAND_99 = {1{`RANDOM}};
  releasedBuffer_rs1prfAddr = _RAND_99[5:0];
  _RAND_100 = {1{`RANDOM}};
  releasedBuffer_rs2prfAddr = _RAND_100[5:0];
  _RAND_101 = {1{`RANDOM}};
  releasedBuffer_prfDest = _RAND_101[5:0];
  _RAND_102 = {1{`RANDOM}};
  releasedBuffer_robAddr = _RAND_102[3:0];
  _RAND_103 = {1{`RANDOM}};
  instrRetired_REG_valid = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  instrRetired_REG_prfAddr = _RAND_104[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module queryScheduler(
  input         clock,
  input         reset,
  output        toCache_queryWithData_query_valid,
  output [31:0] toCache_queryWithData_query_address,
  output [31:0] toCache_queryWithData_query_instruction,
  output [3:0]  toCache_queryWithData_query_branchMask,
  output [3:0]  toCache_queryWithData_query_robAddr,
  output [5:0]  toCache_queryWithData_query_prfDest,
  output [63:0] toCache_queryWithData_data,
  output        toCache_replaying,
  output        storeCommit_ready,
  input         storeCommit_fired,
  input         replaying,
  input         cacheStalled,
  input         replayQueue_query_valid,
  input  [31:0] replayQueue_query_address,
  input  [31:0] replayQueue_query_instruction,
  input  [3:0]  replayQueue_query_branchMask,
  input  [3:0]  replayQueue_query_robAddr,
  input  [5:0]  replayQueue_query_prfDest,
  input  [63:0] replayQueue_data,
  input         branchOps_valid,
  input  [3:0]  branchOps_branchMask,
  input         branchOps_passed,
  input         peripheral_ready,
  output        peripheral_bits_valid,
  output [31:0] peripheral_bits_address,
  output [31:0] peripheral_bits_instruction,
  output [3:0]  peripheral_bits_branchMask,
  output [3:0]  peripheral_bits_robAddr,
  output [5:0]  peripheral_bits_prfDest,
  input         newInstruction_valid,
  input  [31:0] newInstruction_address,
  input  [31:0] newInstruction_instruction,
  input  [3:0]  newInstruction_branchMask,
  input  [3:0]  newInstruction_robAddr,
  input  [5:0]  newInstruction_prfDest,
  output        canAllocate,
  output        clean
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
`endif // RANDOMIZE_REG_INIT
  reg  scheduledInstruction_query_valid; // @[scheduler.scala 52:37]
  reg [31:0] scheduledInstruction_query_address; // @[scheduler.scala 52:37]
  reg [31:0] scheduledInstruction_query_instruction; // @[scheduler.scala 52:37]
  reg [3:0] scheduledInstruction_query_branchMask; // @[scheduler.scala 52:37]
  reg [3:0] scheduledInstruction_query_robAddr; // @[scheduler.scala 52:37]
  reg [5:0] scheduledInstruction_query_prfDest; // @[scheduler.scala 52:37]
  reg [63:0] scheduledInstruction_data; // @[scheduler.scala 52:37]
  reg  dependentReads_0_valid; // @[scheduler.scala 65:31]
  reg [31:0] dependentReads_0_address; // @[scheduler.scala 65:31]
  reg [31:0] dependentReads_0_instruction; // @[scheduler.scala 65:31]
  reg [3:0] dependentReads_0_branchMask; // @[scheduler.scala 65:31]
  reg [3:0] dependentReads_0_robAddr; // @[scheduler.scala 65:31]
  reg [5:0] dependentReads_0_prfDest; // @[scheduler.scala 65:31]
  reg  dependentReads_0_dependency_free; // @[scheduler.scala 65:31]
  reg [3:0] dependentReads_0_dependency_robAddr; // @[scheduler.scala 65:31]
  reg  dependentReads_1_valid; // @[scheduler.scala 65:31]
  reg [31:0] dependentReads_1_address; // @[scheduler.scala 65:31]
  reg [31:0] dependentReads_1_instruction; // @[scheduler.scala 65:31]
  reg [3:0] dependentReads_1_branchMask; // @[scheduler.scala 65:31]
  reg [3:0] dependentReads_1_robAddr; // @[scheduler.scala 65:31]
  reg [5:0] dependentReads_1_prfDest; // @[scheduler.scala 65:31]
  reg  dependentReads_1_dependency_free; // @[scheduler.scala 65:31]
  reg [3:0] dependentReads_1_dependency_robAddr; // @[scheduler.scala 65:31]
  reg  dependentReads_2_valid; // @[scheduler.scala 65:31]
  reg [31:0] dependentReads_2_address; // @[scheduler.scala 65:31]
  reg [31:0] dependentReads_2_instruction; // @[scheduler.scala 65:31]
  reg [3:0] dependentReads_2_branchMask; // @[scheduler.scala 65:31]
  reg [3:0] dependentReads_2_robAddr; // @[scheduler.scala 65:31]
  reg [5:0] dependentReads_2_prfDest; // @[scheduler.scala 65:31]
  reg  dependentReads_2_dependency_free; // @[scheduler.scala 65:31]
  reg [3:0] dependentReads_2_dependency_robAddr; // @[scheduler.scala 65:31]
  reg  dependentReads_3_valid; // @[scheduler.scala 65:31]
  reg [31:0] dependentReads_3_address; // @[scheduler.scala 65:31]
  reg [31:0] dependentReads_3_instruction; // @[scheduler.scala 65:31]
  reg [3:0] dependentReads_3_branchMask; // @[scheduler.scala 65:31]
  reg [3:0] dependentReads_3_robAddr; // @[scheduler.scala 65:31]
  reg [5:0] dependentReads_3_prfDest; // @[scheduler.scala 65:31]
  reg  dependentReads_3_dependency_free; // @[scheduler.scala 65:31]
  reg [3:0] dependentReads_3_dependency_robAddr; // @[scheduler.scala 65:31]
  wire  _dependentRead_T_valid = dependentReads_2_valid ? dependentReads_2_valid : dependentReads_3_valid; // @[Mux.scala 101:16]
  wire [31:0] _dependentRead_T_address = dependentReads_2_valid ? dependentReads_2_address : dependentReads_3_address; // @[Mux.scala 101:16]
  wire [31:0] _dependentRead_T_instruction = dependentReads_2_valid ? dependentReads_2_instruction :
    dependentReads_3_instruction; // @[Mux.scala 101:16]
  wire [3:0] _dependentRead_T_branchMask = dependentReads_2_valid ? dependentReads_2_branchMask :
    dependentReads_3_branchMask; // @[Mux.scala 101:16]
  wire [3:0] _dependentRead_T_robAddr = dependentReads_2_valid ? dependentReads_2_robAddr : dependentReads_3_robAddr; // @[Mux.scala 101:16]
  wire [5:0] _dependentRead_T_prfDest = dependentReads_2_valid ? dependentReads_2_prfDest : dependentReads_3_prfDest; // @[Mux.scala 101:16]
  wire  _dependentRead_T_dependency_free = dependentReads_2_valid ? dependentReads_2_dependency_free :
    dependentReads_3_dependency_free; // @[Mux.scala 101:16]
  wire  _dependentRead_T_1_valid = dependentReads_1_valid ? dependentReads_1_valid : _dependentRead_T_valid; // @[Mux.scala 101:16]
  wire [31:0] _dependentRead_T_1_address = dependentReads_1_valid ? dependentReads_1_address : _dependentRead_T_address; // @[Mux.scala 101:16]
  wire [31:0] _dependentRead_T_1_instruction = dependentReads_1_valid ? dependentReads_1_instruction :
    _dependentRead_T_instruction; // @[Mux.scala 101:16]
  wire [3:0] _dependentRead_T_1_branchMask = dependentReads_1_valid ? dependentReads_1_branchMask :
    _dependentRead_T_branchMask; // @[Mux.scala 101:16]
  wire [3:0] _dependentRead_T_1_robAddr = dependentReads_1_valid ? dependentReads_1_robAddr : _dependentRead_T_robAddr; // @[Mux.scala 101:16]
  wire [5:0] _dependentRead_T_1_prfDest = dependentReads_1_valid ? dependentReads_1_prfDest : _dependentRead_T_prfDest; // @[Mux.scala 101:16]
  wire  _dependentRead_T_1_dependency_free = dependentReads_1_valid ? dependentReads_1_dependency_free :
    _dependentRead_T_dependency_free; // @[Mux.scala 101:16]
  wire  dependentRead_valid = dependentReads_0_valid ? dependentReads_0_valid : _dependentRead_T_1_valid; // @[Mux.scala 101:16]
  wire [31:0] dependentRead_address = dependentReads_0_valid ? dependentReads_0_address : _dependentRead_T_1_address; // @[Mux.scala 101:16]
  wire [31:0] dependentRead_instruction = dependentReads_0_valid ? dependentReads_0_instruction :
    _dependentRead_T_1_instruction; // @[Mux.scala 101:16]
  wire [3:0] dependentRead_branchMask = dependentReads_0_valid ? dependentReads_0_branchMask :
    _dependentRead_T_1_branchMask; // @[Mux.scala 101:16]
  wire [3:0] dependentRead_robAddr = dependentReads_0_valid ? dependentReads_0_robAddr : _dependentRead_T_1_robAddr; // @[Mux.scala 101:16]
  wire [5:0] dependentRead_prfDest = dependentReads_0_valid ? dependentReads_0_prfDest : _dependentRead_T_1_prfDest; // @[Mux.scala 101:16]
  wire  dependentRead_dependency_free = dependentReads_0_valid ? dependentReads_0_dependency_free :
    _dependentRead_T_1_dependency_free; // @[Mux.scala 101:16]
  reg  storeInstructions_0_valid; // @[scheduler.scala 76:34]
  reg [31:0] storeInstructions_0_address; // @[scheduler.scala 76:34]
  reg [31:0] storeInstructions_0_instruction; // @[scheduler.scala 76:34]
  reg [3:0] storeInstructions_0_branchMask; // @[scheduler.scala 76:34]
  reg [3:0] storeInstructions_0_robAddr; // @[scheduler.scala 76:34]
  reg [5:0] storeInstructions_0_prfDest; // @[scheduler.scala 76:34]
  reg  storeInstructions_1_valid; // @[scheduler.scala 76:34]
  reg [31:0] storeInstructions_1_address; // @[scheduler.scala 76:34]
  reg [31:0] storeInstructions_1_instruction; // @[scheduler.scala 76:34]
  reg [3:0] storeInstructions_1_branchMask; // @[scheduler.scala 76:34]
  reg [3:0] storeInstructions_1_robAddr; // @[scheduler.scala 76:34]
  reg [5:0] storeInstructions_1_prfDest; // @[scheduler.scala 76:34]
  reg  storeInstructions_2_valid; // @[scheduler.scala 76:34]
  reg [31:0] storeInstructions_2_address; // @[scheduler.scala 76:34]
  reg [31:0] storeInstructions_2_instruction; // @[scheduler.scala 76:34]
  reg [3:0] storeInstructions_2_branchMask; // @[scheduler.scala 76:34]
  reg [3:0] storeInstructions_2_robAddr; // @[scheduler.scala 76:34]
  reg [5:0] storeInstructions_2_prfDest; // @[scheduler.scala 76:34]
  reg  storeInstructions_3_valid; // @[scheduler.scala 76:34]
  reg [31:0] storeInstructions_3_address; // @[scheduler.scala 76:34]
  reg [31:0] storeInstructions_3_instruction; // @[scheduler.scala 76:34]
  reg [3:0] storeInstructions_3_branchMask; // @[scheduler.scala 76:34]
  reg [3:0] storeInstructions_3_robAddr; // @[scheduler.scala 76:34]
  reg [5:0] storeInstructions_3_prfDest; // @[scheduler.scala 76:34]
  wire  _storeInstruction_T_1_valid = storeInstructions_2_valid ? storeInstructions_2_valid : storeInstructions_3_valid; // @[Mux.scala 101:16]
  wire [31:0] _storeInstruction_T_1_address = storeInstructions_2_valid ? storeInstructions_2_address :
    storeInstructions_3_address; // @[Mux.scala 101:16]
  wire [31:0] _storeInstruction_T_1_instruction = storeInstructions_2_valid ? storeInstructions_2_instruction :
    storeInstructions_3_instruction; // @[Mux.scala 101:16]
  wire [3:0] _storeInstruction_T_1_branchMask = storeInstructions_2_valid ? storeInstructions_2_branchMask :
    storeInstructions_3_branchMask; // @[Mux.scala 101:16]
  wire [3:0] _storeInstruction_T_1_robAddr = storeInstructions_2_valid ? storeInstructions_2_robAddr :
    storeInstructions_3_robAddr; // @[Mux.scala 101:16]
  wire [5:0] _storeInstruction_T_1_prfDest = storeInstructions_2_valid ? storeInstructions_2_prfDest :
    storeInstructions_3_prfDest; // @[Mux.scala 101:16]
  wire  _storeInstruction_T_2_valid = storeInstructions_1_valid ? storeInstructions_1_valid :
    _storeInstruction_T_1_valid; // @[Mux.scala 101:16]
  wire [31:0] _storeInstruction_T_2_address = storeInstructions_1_valid ? storeInstructions_1_address :
    _storeInstruction_T_1_address; // @[Mux.scala 101:16]
  wire [31:0] _storeInstruction_T_2_instruction = storeInstructions_1_valid ? storeInstructions_1_instruction :
    _storeInstruction_T_1_instruction; // @[Mux.scala 101:16]
  wire [3:0] _storeInstruction_T_2_branchMask = storeInstructions_1_valid ? storeInstructions_1_branchMask :
    _storeInstruction_T_1_branchMask; // @[Mux.scala 101:16]
  wire [3:0] _storeInstruction_T_2_robAddr = storeInstructions_1_valid ? storeInstructions_1_robAddr :
    _storeInstruction_T_1_robAddr; // @[Mux.scala 101:16]
  wire [5:0] _storeInstruction_T_2_prfDest = storeInstructions_1_valid ? storeInstructions_1_prfDest :
    _storeInstruction_T_1_prfDest; // @[Mux.scala 101:16]
  wire  storeInstruction_valid = storeInstructions_0_valid ? storeInstructions_0_valid : _storeInstruction_T_2_valid; // @[Mux.scala 101:16]
  wire [3:0] storeInstruction_branchMask = storeInstructions_0_valid ? storeInstructions_0_branchMask :
    _storeInstruction_T_2_branchMask; // @[Mux.scala 101:16]
  reg  fromBuffer_valid; // @[scheduler.scala 86:27]
  reg [31:0] fromBuffer_address; // @[scheduler.scala 86:27]
  reg [31:0] fromBuffer_instruction; // @[scheduler.scala 86:27]
  reg [3:0] fromBuffer_branchMask; // @[scheduler.scala 86:27]
  reg [3:0] fromBuffer_robAddr; // @[scheduler.scala 86:27]
  reg [5:0] fromBuffer_prfDest; // @[scheduler.scala 86:27]
  reg  toCache_replaying_REG; // @[scheduler.scala 92:31]
  reg  toPeripheral; // @[scheduler.scala 117:25]
  wire  _storeInstructionsFree_T = storeInstructions_0_valid & storeInstructions_1_valid; // @[scheduler.scala 141:98]
  wire  _storeInstructionsFree_T_1 = storeInstructions_0_valid & storeInstructions_1_valid & storeInstructions_2_valid; // @[scheduler.scala 141:98]
  wire  _storeInstructionsFree_T_2 = storeInstructions_0_valid & storeInstructions_1_valid & storeInstructions_2_valid
     & storeInstructions_3_valid; // @[scheduler.scala 141:98]
  wire  storeInstructionsFree = storeCommit_fired | ~(storeInstructions_0_valid & storeInstructions_1_valid &
    storeInstructions_2_valid & storeInstructions_3_valid); // @[scheduler.scala 141:54]
  wire  _readCanDequeue_T = dependentReads_0_valid & dependentReads_1_valid; // @[scheduler.scala 145:48]
  wire  _readCanDequeue_T_1 = dependentReads_0_valid & dependentReads_1_valid & dependentReads_2_valid; // @[scheduler.scala 145:48]
  wire  _readCanDequeue_T_4 = dependentRead_valid & dependentRead_dependency_free; // @[scheduler.scala 145:78]
  wire  _readCanDequeue_T_5 = ~(dependentReads_0_valid & dependentReads_1_valid & dependentReads_2_valid &
    dependentReads_3_valid) | dependentRead_valid & dependentRead_dependency_free; // @[scheduler.scala 145:54]
  wire  _readCanDequeue_T_10 = ~(replaying | cacheStalled | _readCanDequeue_T_4 | storeCommit_fired); // @[scheduler.scala 147:9]
  wire  _T_80 = ~branchOps_passed; // @[scheduler.scala 243:12]
  wire [3:0] _T_81 = fromBuffer_branchMask & branchOps_branchMask; // @[scheduler.scala 243:50]
  wire  _T_82 = |_T_81; // @[scheduler.scala 243:74]
  wire  _T_83 = ~branchOps_passed & |_T_81; // @[scheduler.scala 243:30]
  wire  _currDependentReads_newEntry_valid_T_25 = storeInstructions_0_valid & storeInstructions_0_address[31:3] ==
    fromBuffer_address[31:3]; // @[scheduler.scala 221:51]
  wire  _currDependentReads_newEntry_valid_T_29 = storeInstructions_1_valid & storeInstructions_1_address[31:3] ==
    fromBuffer_address[31:3]; // @[scheduler.scala 221:51]
  wire  _currDependentReads_newEntry_valid_T_33 = storeInstructions_2_valid & storeInstructions_2_address[31:3] ==
    fromBuffer_address[31:3]; // @[scheduler.scala 221:51]
  wire  _currDependentReads_newEntry_valid_T_37 = storeInstructions_3_valid & storeInstructions_3_address[31:3] ==
    fromBuffer_address[31:3]; // @[scheduler.scala 221:51]
  wire  _currDependentReads_newEntry_valid_T_40 = storeInstructions_0_valid & storeInstructions_0_address[31:3] ==
    fromBuffer_address[31:3] | storeInstructions_1_valid & storeInstructions_1_address[31:3] == fromBuffer_address[31:3]
     | storeInstructions_2_valid & storeInstructions_2_address[31:3] == fromBuffer_address[31:3] |
    storeInstructions_3_valid & storeInstructions_3_address[31:3] == fromBuffer_address[31:3]; // @[scheduler.scala 221:118]
  wire  _currDependentReads_newEntry_valid_T_41 = scheduledInstruction_query_instruction[5] &
    scheduledInstruction_query_address[31:3] == fromBuffer_address[31:3] & scheduledInstruction_query_valid & ~
    toCache_replaying | _currDependentReads_newEntry_valid_T_40; // @[scheduler.scala 220:192]
  wire  currDependentReads_4_valid = fromBuffer_valid & (~fromBuffer_instruction[5] | fromBuffer_instruction[3] &
    storeInstructionsFree) & _currDependentReads_newEntry_valid_T_41; // @[scheduler.scala 219:174]
  wire  _GEN_112 = ~branchOps_passed & |_T_81 ? 1'h0 : currDependentReads_4_valid; // @[scheduler.scala 238:10 243:{79,92}]
  wire  dependentReadsUpdate_4_valid = branchOps_valid ? _GEN_112 : currDependentReads_4_valid; // @[scheduler.scala 238:10 239:27]
  wire  readCanDequeue = dependentReadsUpdate_4_valid ? _readCanDequeue_T_5 : _readCanDequeue_T_10; // @[scheduler.scala 142:31]
  wire  _dequeuedFromBuffer_T_1 = ~toPeripheral | peripheral_ready; // @[scheduler.scala 154:73]
  wire  _GEN_0 = 5'hb == fromBuffer_instruction[6:2] & (readCanDequeue & storeInstructionsFree); // @[scheduler.scala 149:44 157:30]
  wire  _GEN_1 = 5'h8 == fromBuffer_instruction[6:2] ? storeInstructionsFree & (~toPeripheral | peripheral_ready) :
    _GEN_0; // @[scheduler.scala 149:44 154:30]
  wire  _GEN_2 = 5'h0 == fromBuffer_instruction[6:2] ? readCanDequeue : _GEN_1; // @[scheduler.scala 149:44 151:30]
  wire  dequeuedFromBuffer = fromBuffer_valid & _GEN_2; // @[scheduler.scala 135:26]
  wire  _T_4 = ~cacheStalled; // @[scheduler.scala 163:22]
  wire  _GEN_5 = cacheStalled ? 1'h0 : scheduledInstruction_query_valid; // @[scheduler.scala 164:{27,62} 52:37]
  wire  _storeInstructionsUpdate_4_valid_T_6 = fromBuffer_valid & fromBuffer_instruction[5] & _dequeuedFromBuffer_T_1 &
    dequeuedFromBuffer; // @[scheduler.scala 187:97]
  wire [3:0] _storeInstructionsUpdate_4_valid_T_7 = branchOps_branchMask & fromBuffer_branchMask; // @[scheduler.scala 188:51]
  wire  storeInstructionsUpdate_4_valid = _storeInstructionsUpdate_4_valid_T_6 & ~(branchOps_valid & |
    _storeInstructionsUpdate_4_valid_T_7 & _T_80); // @[scheduler.scala 188:5]
  wire  _GEN_189 = toPeripheral | dependentReadsUpdate_4_valid | storeInstructionsUpdate_4_valid & ~
    fromBuffer_instruction[3] ? 1'h0 : fromBuffer_valid; // @[scheduler.scala 283:175 281:25 284:33]
  wire  _GEN_191 = ~dequeuedFromBuffer | toPeripheral ? 1'h0 : _GEN_189; // @[scheduler.scala 289:47 290:33]
  wire  _GEN_197 = _readCanDequeue_T_4 ? dependentRead_valid : _GEN_191; // @[scheduler.scala 272:67 278:31]
  wire  _GEN_198 = storeCommit_fired ? storeInstruction_valid : _GEN_197; // @[scheduler.scala 271:{32,54}]
  wire  nextScheduled_query_valid = replaying ? replayQueue_query_valid : _GEN_198; // @[scheduler.scala 270:{19,35}]
  wire  _GEN_6 = replaying | ~cacheStalled ? nextScheduled_query_valid : _GEN_5; // @[scheduler.scala 163:{38,61}]
  wire [2:0] _T_182 = {fromBuffer_instruction[28],fromBuffer_instruction[27],fromBuffer_instruction[3]}; // @[Cat.scala 33:92]
  wire [31:0] _nextScheduled_query_instruction_T_3 = {fromBuffer_instruction[31:7],7'hf}; // @[Cat.scala 33:92]
  wire [31:0] _nextScheduled_query_instruction_T_1 = {fromBuffer_instruction[31:7],7'h3}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_190 = _T_182 == 3'h7 ? _nextScheduled_query_instruction_T_3 : _nextScheduled_query_instruction_T_1; // @[scheduler.scala 282:37 286:80 287:39]
  wire [3:0] _GEN_193 = _readCanDequeue_T_4 ? dependentRead_branchMask : fromBuffer_branchMask; // @[scheduler.scala 272:67 274:36 281:25]
  wire [3:0] _GEN_201 = storeCommit_fired ? storeInstruction_branchMask : _GEN_193; // @[scheduler.scala 271:{32,54}]
  wire [3:0] nextScheduled_query_branchMask = replaying ? replayQueue_query_branchMask : _GEN_201; // @[scheduler.scala 270:{19,35}]
  wire [3:0] _GEN_9 = replaying | ~cacheStalled ? nextScheduled_query_branchMask : scheduledInstruction_query_branchMask
    ; // @[scheduler.scala 163:{38,61} 52:37]
  wire [3:0] _T_6 = nextScheduled_query_branchMask & branchOps_branchMask; // @[scheduler.scala 166:42]
  wire  _T_7 = |_T_6; // @[scheduler.scala 166:66]
  wire [3:0] _scheduledInstruction_query_branchMask_T = nextScheduled_query_branchMask ^ branchOps_branchMask; // @[scheduler.scala 167:79]
  wire [3:0] _T_12 = storeInstructions_0_branchMask & branchOps_branchMask; // @[scheduler.scala 178:29]
  wire  _T_13 = |_T_12; // @[scheduler.scala 178:53]
  wire [3:0] _storeInstructionsUpdate_0_branchMask_T = storeInstructions_0_branchMask ^ branchOps_branchMask; // @[scheduler.scala 178:96]
  wire  _GEN_18 = _T_80 & _T_13 ? 1'h0 : storeInstructions_0_valid; // @[scheduler.scala 176:10 179:{79,92}]
  wire  _GEN_20 = branchOps_valid ? _GEN_18 : storeInstructions_0_valid; // @[scheduler.scala 176:10 177:27]
  wire [3:0] _T_18 = storeInstructions_1_branchMask & branchOps_branchMask; // @[scheduler.scala 178:29]
  wire  _T_19 = |_T_18; // @[scheduler.scala 178:53]
  wire [3:0] _storeInstructionsUpdate_1_branchMask_T = storeInstructions_1_branchMask ^ branchOps_branchMask; // @[scheduler.scala 178:96]
  wire [3:0] _GEN_21 = |_T_18 ? _storeInstructionsUpdate_1_branchMask_T : storeInstructions_1_branchMask; // @[scheduler.scala 176:10 178:{59,77}]
  wire  _GEN_22 = _T_80 & _T_19 ? 1'h0 : storeInstructions_1_valid; // @[scheduler.scala 176:10 179:{79,92}]
  wire [3:0] storeInstructionsUpdate_1_branchMask = branchOps_valid ? _GEN_21 : storeInstructions_1_branchMask; // @[scheduler.scala 176:10 177:27]
  wire  storeInstructionsUpdate_1_valid = branchOps_valid ? _GEN_22 : storeInstructions_1_valid; // @[scheduler.scala 176:10 177:27]
  wire [3:0] _T_24 = storeInstructions_2_branchMask & branchOps_branchMask; // @[scheduler.scala 178:29]
  wire  _T_25 = |_T_24; // @[scheduler.scala 178:53]
  wire [3:0] _storeInstructionsUpdate_2_branchMask_T = storeInstructions_2_branchMask ^ branchOps_branchMask; // @[scheduler.scala 178:96]
  wire [3:0] _GEN_25 = |_T_24 ? _storeInstructionsUpdate_2_branchMask_T : storeInstructions_2_branchMask; // @[scheduler.scala 176:10 178:{59,77}]
  wire  _GEN_26 = _T_80 & _T_25 ? 1'h0 : storeInstructions_2_valid; // @[scheduler.scala 176:10 179:{79,92}]
  wire [3:0] storeInstructionsUpdate_2_branchMask = branchOps_valid ? _GEN_25 : storeInstructions_2_branchMask; // @[scheduler.scala 176:10 177:27]
  wire  storeInstructionsUpdate_2_valid = branchOps_valid ? _GEN_26 : storeInstructions_2_valid; // @[scheduler.scala 176:10 177:27]
  wire [3:0] _T_30 = storeInstructions_3_branchMask & branchOps_branchMask; // @[scheduler.scala 178:29]
  wire  _T_31 = |_T_30; // @[scheduler.scala 178:53]
  wire [3:0] _storeInstructionsUpdate_3_branchMask_T = storeInstructions_3_branchMask ^ branchOps_branchMask; // @[scheduler.scala 178:96]
  wire [3:0] _GEN_29 = |_T_30 ? _storeInstructionsUpdate_3_branchMask_T : storeInstructions_3_branchMask; // @[scheduler.scala 176:10 178:{59,77}]
  wire  _GEN_30 = _T_80 & _T_31 ? 1'h0 : storeInstructions_3_valid; // @[scheduler.scala 176:10 179:{79,92}]
  wire [3:0] storeInstructionsUpdate_3_branchMask = branchOps_valid ? _GEN_29 : storeInstructions_3_branchMask; // @[scheduler.scala 176:10 177:27]
  wire  storeInstructionsUpdate_3_valid = branchOps_valid ? _GEN_30 : storeInstructions_3_valid; // @[scheduler.scala 176:10 177:27]
  wire [3:0] _storeInstructionsUpdate_4_branchMask_T = fromBuffer_branchMask ^ branchOps_branchMask; // @[scheduler.scala 178:96]
  wire [3:0] _GEN_33 = _T_82 ? _storeInstructionsUpdate_4_branchMask_T : fromBuffer_branchMask; // @[scheduler.scala 176:10 178:{59,77}]
  wire [3:0] storeInstructionsUpdate_4_branchMask = branchOps_valid ? _GEN_33 : fromBuffer_branchMask; // @[scheduler.scala 176:10 177:27]
  wire [3:0] _currDependentReads_newEntry_dependency_robAddr_T_16 = _currDependentReads_newEntry_valid_T_25 ?
    storeInstructions_0_robAddr : scheduledInstruction_query_robAddr; // @[Mux.scala 101:16]
  wire [3:0] _currDependentReads_newEntry_dependency_robAddr_T_17 = _currDependentReads_newEntry_valid_T_29 ?
    storeInstructions_1_robAddr : _currDependentReads_newEntry_dependency_robAddr_T_16; // @[Mux.scala 101:16]
  wire [3:0] _currDependentReads_newEntry_dependency_robAddr_T_18 = _currDependentReads_newEntry_valid_T_33 ?
    storeInstructions_2_robAddr : _currDependentReads_newEntry_dependency_robAddr_T_17; // @[Mux.scala 101:16]
  wire [3:0] currDependentReads_4_dependency_robAddr = _currDependentReads_newEntry_valid_T_37 ?
    storeInstructions_3_robAddr : _currDependentReads_newEntry_dependency_robAddr_T_18; // @[Mux.scala 101:16]
  wire [3:0] _T_50 = dependentReads_0_branchMask & branchOps_branchMask; // @[scheduler.scala 240:29]
  wire  _T_51 = |_T_50; // @[scheduler.scala 240:53]
  wire [3:0] _dependentReadsUpdate_0_branchMask_T = dependentReads_0_branchMask ^ branchOps_branchMask; // @[scheduler.scala 241:44]
  wire  _GEN_88 = ~branchOps_passed & _T_51 ? 1'h0 : dependentReads_0_valid; // @[scheduler.scala 238:10 243:{79,92}]
  wire  _GEN_90 = branchOps_valid ? _GEN_88 : dependentReads_0_valid; // @[scheduler.scala 238:10 239:27]
  reg  REG; // @[scheduler.scala 245:17]
  wire  _GEN_91 = dependentReads_0_dependency_robAddr == scheduledInstruction_query_robAddr |
    dependentReads_0_dependency_free; // @[scheduler.scala 238:10 247:{76,99}]
  wire [3:0] _T_57 = dependentReads_1_branchMask & branchOps_branchMask; // @[scheduler.scala 240:29]
  wire  _T_58 = |_T_57; // @[scheduler.scala 240:53]
  wire [3:0] _dependentReadsUpdate_1_branchMask_T = dependentReads_1_branchMask ^ branchOps_branchMask; // @[scheduler.scala 241:44]
  wire [3:0] _GEN_93 = |_T_57 ? _dependentReadsUpdate_1_branchMask_T : dependentReads_1_branchMask; // @[scheduler.scala 238:10 240:58 241:25]
  wire  _GEN_94 = ~branchOps_passed & _T_58 ? 1'h0 : dependentReads_1_valid; // @[scheduler.scala 238:10 243:{79,92}]
  wire [3:0] dependentReadsUpdate_1_branchMask = branchOps_valid ? _GEN_93 : dependentReads_1_branchMask; // @[scheduler.scala 238:10 239:27]
  wire  _GEN_96 = branchOps_valid ? _GEN_94 : dependentReads_1_valid; // @[scheduler.scala 238:10 239:27]
  reg  REG_1; // @[scheduler.scala 245:17]
  wire  _GEN_97 = dependentReads_1_dependency_robAddr == scheduledInstruction_query_robAddr |
    dependentReads_1_dependency_free; // @[scheduler.scala 238:10 247:{76,99}]
  wire  dependentReadsUpdate_1_dependency_free = REG_1 ? _GEN_97 : dependentReads_1_dependency_free; // @[scheduler.scala 238:10 245:38]
  wire [3:0] _T_64 = dependentReads_2_branchMask & branchOps_branchMask; // @[scheduler.scala 240:29]
  wire  _T_65 = |_T_64; // @[scheduler.scala 240:53]
  wire [3:0] _dependentReadsUpdate_2_branchMask_T = dependentReads_2_branchMask ^ branchOps_branchMask; // @[scheduler.scala 241:44]
  wire [3:0] _GEN_99 = |_T_64 ? _dependentReadsUpdate_2_branchMask_T : dependentReads_2_branchMask; // @[scheduler.scala 238:10 240:58 241:25]
  wire  _GEN_100 = ~branchOps_passed & _T_65 ? 1'h0 : dependentReads_2_valid; // @[scheduler.scala 238:10 243:{79,92}]
  wire [3:0] dependentReadsUpdate_2_branchMask = branchOps_valid ? _GEN_99 : dependentReads_2_branchMask; // @[scheduler.scala 238:10 239:27]
  wire  _GEN_102 = branchOps_valid ? _GEN_100 : dependentReads_2_valid; // @[scheduler.scala 238:10 239:27]
  reg  REG_2; // @[scheduler.scala 245:17]
  wire  _GEN_103 = dependentReads_2_dependency_robAddr == scheduledInstruction_query_robAddr |
    dependentReads_2_dependency_free; // @[scheduler.scala 238:10 247:{76,99}]
  wire  dependentReadsUpdate_2_dependency_free = REG_2 ? _GEN_103 : dependentReads_2_dependency_free; // @[scheduler.scala 238:10 245:38]
  wire [3:0] _T_71 = dependentReads_3_branchMask & branchOps_branchMask; // @[scheduler.scala 240:29]
  wire  _T_72 = |_T_71; // @[scheduler.scala 240:53]
  wire [3:0] _dependentReadsUpdate_3_branchMask_T = dependentReads_3_branchMask ^ branchOps_branchMask; // @[scheduler.scala 241:44]
  wire [3:0] _GEN_105 = |_T_71 ? _dependentReadsUpdate_3_branchMask_T : dependentReads_3_branchMask; // @[scheduler.scala 238:10 240:58 241:25]
  wire  _GEN_106 = ~branchOps_passed & _T_72 ? 1'h0 : dependentReads_3_valid; // @[scheduler.scala 238:10 243:{79,92}]
  wire [3:0] dependentReadsUpdate_3_branchMask = branchOps_valid ? _GEN_105 : dependentReads_3_branchMask; // @[scheduler.scala 238:10 239:27]
  wire  _GEN_108 = branchOps_valid ? _GEN_106 : dependentReads_3_valid; // @[scheduler.scala 238:10 239:27]
  reg  REG_3; // @[scheduler.scala 245:17]
  wire  _GEN_109 = dependentReads_3_dependency_robAddr == scheduledInstruction_query_robAddr |
    dependentReads_3_dependency_free; // @[scheduler.scala 238:10 247:{76,99}]
  wire  dependentReadsUpdate_3_dependency_free = REG_3 ? _GEN_109 : dependentReads_3_dependency_free; // @[scheduler.scala 238:10 245:38]
  reg  REG_4; // @[scheduler.scala 245:17]
  wire  _T_84 = currDependentReads_4_dependency_robAddr == scheduledInstruction_query_robAddr; // @[scheduler.scala 247:36]
  wire  dependentReadsUpdate_4_dependency_free = REG_4 & _T_84; // @[scheduler.scala 238:10 245:38]
  wire  _T_91 = ~replaying & _T_4 & ~storeCommit_fired & dependentRead_valid & dependentRead_dependency_free; // @[scheduler.scala 252:81]
  wire  _T_92 = dependentReads_0_valid & dependentReads_0_dependency_free; // @[scheduler.scala 253:45]
  wire  _T_93 = dependentReads_1_valid & dependentReads_1_dependency_free; // @[scheduler.scala 253:45]
  wire  _T_94 = dependentReads_2_valid & dependentReads_2_dependency_free; // @[scheduler.scala 253:45]
  wire  _T_97 = _T_92 | _T_93; // @[scheduler.scala 254:26]
  wire  _T_98 = _T_92 | _T_93 | _T_94; // @[scheduler.scala 254:26]
  wire  _GEN_117 = dependentReads_0_dependency_free ? 1'h0 : _GEN_90; // @[scheduler.scala 256:{108,123}]
  wire  _GEN_118 = ~_T_92 & dependentReads_1_dependency_free ? 1'h0 : _GEN_96; // @[scheduler.scala 256:{108,123}]
  wire  _GEN_119 = ~_T_97 & dependentReads_2_dependency_free ? 1'h0 : _GEN_102; // @[scheduler.scala 256:{108,123}]
  wire  _GEN_120 = ~_T_98 & dependentReads_3_dependency_free ? 1'h0 : _GEN_108; // @[scheduler.scala 256:{108,123}]
  wire  dependentReadsUpdate_1_valid = ~replaying & _T_4 & ~storeCommit_fired & dependentRead_valid &
    dependentRead_dependency_free ? _GEN_118 : _GEN_96; // @[scheduler.scala 252:115]
  wire  dependentReadsUpdate_2_valid = ~replaying & _T_4 & ~storeCommit_fired & dependentRead_valid &
    dependentRead_dependency_free ? _GEN_119 : _GEN_102; // @[scheduler.scala 252:115]
  wire  dependentReadsUpdate_3_valid = ~replaying & _T_4 & ~storeCommit_fired & dependentRead_valid &
    dependentRead_dependency_free ? _GEN_120 : _GEN_108; // @[scheduler.scala 252:115]
  reg  bufferQueue_0_valid; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_0_address; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_0_instruction; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_0_branchMask; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_0_robAddr; // @[scheduler.scala 294:28]
  reg [5:0] bufferQueue_0_prfDest; // @[scheduler.scala 294:28]
  reg  bufferQueue_1_valid; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_1_address; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_1_instruction; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_1_branchMask; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_1_robAddr; // @[scheduler.scala 294:28]
  reg [5:0] bufferQueue_1_prfDest; // @[scheduler.scala 294:28]
  reg  bufferQueue_2_valid; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_2_address; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_2_instruction; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_2_branchMask; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_2_robAddr; // @[scheduler.scala 294:28]
  reg [5:0] bufferQueue_2_prfDest; // @[scheduler.scala 294:28]
  reg  bufferQueue_3_valid; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_3_address; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_3_instruction; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_3_branchMask; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_3_robAddr; // @[scheduler.scala 294:28]
  reg [5:0] bufferQueue_3_prfDest; // @[scheduler.scala 294:28]
  reg  bufferQueue_4_valid; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_4_address; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_4_instruction; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_4_branchMask; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_4_robAddr; // @[scheduler.scala 294:28]
  reg [5:0] bufferQueue_4_prfDest; // @[scheduler.scala 294:28]
  reg  bufferQueue_5_valid; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_5_address; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_5_instruction; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_5_branchMask; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_5_robAddr; // @[scheduler.scala 294:28]
  reg [5:0] bufferQueue_5_prfDest; // @[scheduler.scala 294:28]
  reg  bufferQueue_6_valid; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_6_address; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_6_instruction; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_6_branchMask; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_6_robAddr; // @[scheduler.scala 294:28]
  reg [5:0] bufferQueue_6_prfDest; // @[scheduler.scala 294:28]
  reg  bufferQueue_7_valid; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_7_address; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_7_instruction; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_7_branchMask; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_7_robAddr; // @[scheduler.scala 294:28]
  reg [5:0] bufferQueue_7_prfDest; // @[scheduler.scala 294:28]
  reg  bufferQueue_8_valid; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_8_address; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_8_instruction; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_8_branchMask; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_8_robAddr; // @[scheduler.scala 294:28]
  reg [5:0] bufferQueue_8_prfDest; // @[scheduler.scala 294:28]
  reg  bufferQueue_9_valid; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_9_address; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_9_instruction; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_9_branchMask; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_9_robAddr; // @[scheduler.scala 294:28]
  reg [5:0] bufferQueue_9_prfDest; // @[scheduler.scala 294:28]
  reg  bufferQueue_10_valid; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_10_address; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_10_instruction; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_10_branchMask; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_10_robAddr; // @[scheduler.scala 294:28]
  reg [5:0] bufferQueue_10_prfDest; // @[scheduler.scala 294:28]
  reg  bufferQueue_11_valid; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_11_address; // @[scheduler.scala 294:28]
  reg [31:0] bufferQueue_11_instruction; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_11_branchMask; // @[scheduler.scala 294:28]
  reg [3:0] bufferQueue_11_robAddr; // @[scheduler.scala 294:28]
  reg [5:0] bufferQueue_11_prfDest; // @[scheduler.scala 294:28]
  wire  _T_187 = bufferQueue_0_valid & bufferQueue_1_valid; // @[scheduler.scala 300:48]
  wire  _T_188 = bufferQueue_0_valid & bufferQueue_1_valid & bufferQueue_2_valid; // @[scheduler.scala 300:48]
  wire  _T_189 = bufferQueue_0_valid & bufferQueue_1_valid & bufferQueue_2_valid & bufferQueue_3_valid; // @[scheduler.scala 300:48]
  wire  _T_190 = bufferQueue_0_valid & bufferQueue_1_valid & bufferQueue_2_valid & bufferQueue_3_valid &
    bufferQueue_4_valid; // @[scheduler.scala 300:48]
  wire  _T_191 = bufferQueue_0_valid & bufferQueue_1_valid & bufferQueue_2_valid & bufferQueue_3_valid &
    bufferQueue_4_valid & bufferQueue_5_valid; // @[scheduler.scala 300:48]
  wire  _T_192 = bufferQueue_0_valid & bufferQueue_1_valid & bufferQueue_2_valid & bufferQueue_3_valid &
    bufferQueue_4_valid & bufferQueue_5_valid & bufferQueue_6_valid; // @[scheduler.scala 300:48]
  wire  _T_193 = bufferQueue_0_valid & bufferQueue_1_valid & bufferQueue_2_valid & bufferQueue_3_valid &
    bufferQueue_4_valid & bufferQueue_5_valid & bufferQueue_6_valid & bufferQueue_7_valid; // @[scheduler.scala 300:48]
  wire  _T_194 = bufferQueue_0_valid & bufferQueue_1_valid & bufferQueue_2_valid & bufferQueue_3_valid &
    bufferQueue_4_valid & bufferQueue_5_valid & bufferQueue_6_valid & bufferQueue_7_valid & bufferQueue_8_valid; // @[scheduler.scala 300:48]
  wire  _T_195 = bufferQueue_0_valid & bufferQueue_1_valid & bufferQueue_2_valid & bufferQueue_3_valid &
    bufferQueue_4_valid & bufferQueue_5_valid & bufferQueue_6_valid & bufferQueue_7_valid & bufferQueue_8_valid &
    bufferQueue_9_valid; // @[scheduler.scala 300:48]
  wire  _T_196 = bufferQueue_0_valid & bufferQueue_1_valid & bufferQueue_2_valid & bufferQueue_3_valid &
    bufferQueue_4_valid & bufferQueue_5_valid & bufferQueue_6_valid & bufferQueue_7_valid & bufferQueue_8_valid &
    bufferQueue_9_valid & bufferQueue_10_valid; // @[scheduler.scala 300:48]
  wire  _T_199 = ~bufferQueue_0_valid; // @[scheduler.scala 302:86]
  wire [3:0] _T_243 = bufferQueue_1_branchMask & branchOps_branchMask; // @[scheduler.scala 308:50]
  wire  _T_244 = |_T_243; // @[scheduler.scala 308:74]
  wire  _GEN_287 = _T_80 & |_T_243 ? 1'h0 : bufferQueue_1_valid; // @[scheduler.scala 305:12 308:{79,94}]
  wire  _GEN_289 = branchOps_valid ? _GEN_287 : bufferQueue_1_valid; // @[scheduler.scala 305:12 306:28]
  wire  _GEN_343 = _T_199 & bufferQueue_1_valid ? 1'h0 : _GEN_289; // @[scheduler.scala 341:{107,92}]
  wire  bufferQueueUpdate_1_valid = (dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1 ? _GEN_343 :
    _GEN_289; // @[scheduler.scala 334:90]
  wire [3:0] _T_237 = bufferQueue_0_branchMask & branchOps_branchMask; // @[scheduler.scala 308:50]
  wire  _T_238 = |_T_237; // @[scheduler.scala 308:74]
  wire  _GEN_283 = _T_80 & |_T_237 ? 1'h0 : bufferQueue_0_valid; // @[scheduler.scala 305:12 308:{79,94}]
  wire  _GEN_285 = branchOps_valid ? _GEN_283 : bufferQueue_0_valid; // @[scheduler.scala 305:12 306:28]
  wire  _GEN_342 = bufferQueue_0_valid ? 1'h0 : _GEN_285; // @[scheduler.scala 341:{107,92}]
  wire [3:0] _bufferQueueUpdate_1_branchMask_T = bufferQueue_1_branchMask ^ branchOps_branchMask; // @[scheduler.scala 307:96]
  wire [3:0] _GEN_286 = _T_244 ? _bufferQueueUpdate_1_branchMask_T : bufferQueue_1_branchMask; // @[scheduler.scala 305:12 307:{58,77}]
  wire [3:0] bufferQueueUpdate_1_branchMask = branchOps_valid ? _GEN_286 : bufferQueue_1_branchMask; // @[scheduler.scala 305:12 306:28]
  wire [3:0] _bufferQueueUpdate_0_branchMask_T = bufferQueue_0_branchMask ^ branchOps_branchMask; // @[scheduler.scala 307:96]
  wire  _T_332 = bufferQueue_0_valid | bufferQueue_1_valid; // @[scheduler.scala 339:50]
  wire [3:0] _T_249 = bufferQueue_2_branchMask & branchOps_branchMask; // @[scheduler.scala 308:50]
  wire  _T_250 = |_T_249; // @[scheduler.scala 308:74]
  wire  _GEN_291 = _T_80 & |_T_249 ? 1'h0 : bufferQueue_2_valid; // @[scheduler.scala 305:12 308:{79,94}]
  wire  _GEN_293 = branchOps_valid ? _GEN_291 : bufferQueue_2_valid; // @[scheduler.scala 305:12 306:28]
  wire  _GEN_344 = ~_T_332 & bufferQueue_2_valid ? 1'h0 : _GEN_293; // @[scheduler.scala 341:{107,92}]
  wire  bufferQueueUpdate_2_valid = (dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1 ? _GEN_344 :
    _GEN_293; // @[scheduler.scala 334:90]
  wire [3:0] _bufferQueueUpdate_2_branchMask_T = bufferQueue_2_branchMask ^ branchOps_branchMask; // @[scheduler.scala 307:96]
  wire [3:0] _GEN_290 = _T_250 ? _bufferQueueUpdate_2_branchMask_T : bufferQueue_2_branchMask; // @[scheduler.scala 305:12 307:{58,77}]
  wire [3:0] bufferQueueUpdate_2_branchMask = branchOps_valid ? _GEN_290 : bufferQueue_2_branchMask; // @[scheduler.scala 305:12 306:28]
  wire  _T_333 = bufferQueue_0_valid | bufferQueue_1_valid | bufferQueue_2_valid; // @[scheduler.scala 339:50]
  wire [3:0] _T_255 = bufferQueue_3_branchMask & branchOps_branchMask; // @[scheduler.scala 308:50]
  wire  _T_256 = |_T_255; // @[scheduler.scala 308:74]
  wire  _GEN_295 = _T_80 & |_T_255 ? 1'h0 : bufferQueue_3_valid; // @[scheduler.scala 305:12 308:{79,94}]
  wire  _GEN_297 = branchOps_valid ? _GEN_295 : bufferQueue_3_valid; // @[scheduler.scala 305:12 306:28]
  wire  _GEN_345 = ~_T_333 & bufferQueue_3_valid ? 1'h0 : _GEN_297; // @[scheduler.scala 341:{107,92}]
  wire  bufferQueueUpdate_3_valid = (dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1 ? _GEN_345 :
    _GEN_297; // @[scheduler.scala 334:90]
  wire [3:0] _bufferQueueUpdate_3_branchMask_T = bufferQueue_3_branchMask ^ branchOps_branchMask; // @[scheduler.scala 307:96]
  wire [3:0] _GEN_294 = _T_256 ? _bufferQueueUpdate_3_branchMask_T : bufferQueue_3_branchMask; // @[scheduler.scala 305:12 307:{58,77}]
  wire [3:0] bufferQueueUpdate_3_branchMask = branchOps_valid ? _GEN_294 : bufferQueue_3_branchMask; // @[scheduler.scala 305:12 306:28]
  wire  _T_334 = bufferQueue_0_valid | bufferQueue_1_valid | bufferQueue_2_valid | bufferQueue_3_valid; // @[scheduler.scala 339:50]
  wire [3:0] _T_261 = bufferQueue_4_branchMask & branchOps_branchMask; // @[scheduler.scala 308:50]
  wire  _T_262 = |_T_261; // @[scheduler.scala 308:74]
  wire  _GEN_299 = _T_80 & |_T_261 ? 1'h0 : bufferQueue_4_valid; // @[scheduler.scala 305:12 308:{79,94}]
  wire  _GEN_301 = branchOps_valid ? _GEN_299 : bufferQueue_4_valid; // @[scheduler.scala 305:12 306:28]
  wire  _GEN_346 = ~_T_334 & bufferQueue_4_valid ? 1'h0 : _GEN_301; // @[scheduler.scala 341:{107,92}]
  wire  bufferQueueUpdate_4_valid = (dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1 ? _GEN_346 :
    _GEN_301; // @[scheduler.scala 334:90]
  wire [3:0] _bufferQueueUpdate_4_branchMask_T = bufferQueue_4_branchMask ^ branchOps_branchMask; // @[scheduler.scala 307:96]
  wire [3:0] _GEN_298 = _T_262 ? _bufferQueueUpdate_4_branchMask_T : bufferQueue_4_branchMask; // @[scheduler.scala 305:12 307:{58,77}]
  wire [3:0] bufferQueueUpdate_4_branchMask = branchOps_valid ? _GEN_298 : bufferQueue_4_branchMask; // @[scheduler.scala 305:12 306:28]
  wire  _T_335 = bufferQueue_0_valid | bufferQueue_1_valid | bufferQueue_2_valid | bufferQueue_3_valid |
    bufferQueue_4_valid; // @[scheduler.scala 339:50]
  wire [3:0] _T_267 = bufferQueue_5_branchMask & branchOps_branchMask; // @[scheduler.scala 308:50]
  wire  _T_268 = |_T_267; // @[scheduler.scala 308:74]
  wire  _GEN_303 = _T_80 & |_T_267 ? 1'h0 : bufferQueue_5_valid; // @[scheduler.scala 305:12 308:{79,94}]
  wire  _GEN_305 = branchOps_valid ? _GEN_303 : bufferQueue_5_valid; // @[scheduler.scala 305:12 306:28]
  wire  _GEN_347 = ~_T_335 & bufferQueue_5_valid ? 1'h0 : _GEN_305; // @[scheduler.scala 341:{107,92}]
  wire  bufferQueueUpdate_5_valid = (dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1 ? _GEN_347 :
    _GEN_305; // @[scheduler.scala 334:90]
  wire [3:0] _bufferQueueUpdate_5_branchMask_T = bufferQueue_5_branchMask ^ branchOps_branchMask; // @[scheduler.scala 307:96]
  wire [3:0] _GEN_302 = _T_268 ? _bufferQueueUpdate_5_branchMask_T : bufferQueue_5_branchMask; // @[scheduler.scala 305:12 307:{58,77}]
  wire [3:0] bufferQueueUpdate_5_branchMask = branchOps_valid ? _GEN_302 : bufferQueue_5_branchMask; // @[scheduler.scala 305:12 306:28]
  wire  _T_336 = bufferQueue_0_valid | bufferQueue_1_valid | bufferQueue_2_valid | bufferQueue_3_valid |
    bufferQueue_4_valid | bufferQueue_5_valid; // @[scheduler.scala 339:50]
  wire [3:0] _T_273 = bufferQueue_6_branchMask & branchOps_branchMask; // @[scheduler.scala 308:50]
  wire  _T_274 = |_T_273; // @[scheduler.scala 308:74]
  wire  _GEN_307 = _T_80 & |_T_273 ? 1'h0 : bufferQueue_6_valid; // @[scheduler.scala 305:12 308:{79,94}]
  wire  _GEN_309 = branchOps_valid ? _GEN_307 : bufferQueue_6_valid; // @[scheduler.scala 305:12 306:28]
  wire  _GEN_348 = ~_T_336 & bufferQueue_6_valid ? 1'h0 : _GEN_309; // @[scheduler.scala 341:{107,92}]
  wire  bufferQueueUpdate_6_valid = (dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1 ? _GEN_348 :
    _GEN_309; // @[scheduler.scala 334:90]
  wire [3:0] _bufferQueueUpdate_6_branchMask_T = bufferQueue_6_branchMask ^ branchOps_branchMask; // @[scheduler.scala 307:96]
  wire [3:0] _GEN_306 = _T_274 ? _bufferQueueUpdate_6_branchMask_T : bufferQueue_6_branchMask; // @[scheduler.scala 305:12 307:{58,77}]
  wire [3:0] bufferQueueUpdate_6_branchMask = branchOps_valid ? _GEN_306 : bufferQueue_6_branchMask; // @[scheduler.scala 305:12 306:28]
  wire  _T_337 = bufferQueue_0_valid | bufferQueue_1_valid | bufferQueue_2_valid | bufferQueue_3_valid |
    bufferQueue_4_valid | bufferQueue_5_valid | bufferQueue_6_valid; // @[scheduler.scala 339:50]
  wire [3:0] _T_279 = bufferQueue_7_branchMask & branchOps_branchMask; // @[scheduler.scala 308:50]
  wire  _T_280 = |_T_279; // @[scheduler.scala 308:74]
  wire  _GEN_311 = _T_80 & |_T_279 ? 1'h0 : bufferQueue_7_valid; // @[scheduler.scala 305:12 308:{79,94}]
  wire  _GEN_313 = branchOps_valid ? _GEN_311 : bufferQueue_7_valid; // @[scheduler.scala 305:12 306:28]
  wire  _GEN_349 = ~_T_337 & bufferQueue_7_valid ? 1'h0 : _GEN_313; // @[scheduler.scala 341:{107,92}]
  wire  bufferQueueUpdate_7_valid = (dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1 ? _GEN_349 :
    _GEN_313; // @[scheduler.scala 334:90]
  wire [3:0] _bufferQueueUpdate_7_branchMask_T = bufferQueue_7_branchMask ^ branchOps_branchMask; // @[scheduler.scala 307:96]
  wire [3:0] _GEN_310 = _T_280 ? _bufferQueueUpdate_7_branchMask_T : bufferQueue_7_branchMask; // @[scheduler.scala 305:12 307:{58,77}]
  wire [3:0] bufferQueueUpdate_7_branchMask = branchOps_valid ? _GEN_310 : bufferQueue_7_branchMask; // @[scheduler.scala 305:12 306:28]
  wire  _T_338 = bufferQueue_0_valid | bufferQueue_1_valid | bufferQueue_2_valid | bufferQueue_3_valid |
    bufferQueue_4_valid | bufferQueue_5_valid | bufferQueue_6_valid | bufferQueue_7_valid; // @[scheduler.scala 339:50]
  wire [3:0] _T_285 = bufferQueue_8_branchMask & branchOps_branchMask; // @[scheduler.scala 308:50]
  wire  _T_286 = |_T_285; // @[scheduler.scala 308:74]
  wire  _GEN_315 = _T_80 & |_T_285 ? 1'h0 : bufferQueue_8_valid; // @[scheduler.scala 305:12 308:{79,94}]
  wire  _GEN_317 = branchOps_valid ? _GEN_315 : bufferQueue_8_valid; // @[scheduler.scala 305:12 306:28]
  wire  _GEN_350 = ~_T_338 & bufferQueue_8_valid ? 1'h0 : _GEN_317; // @[scheduler.scala 341:{107,92}]
  wire  bufferQueueUpdate_8_valid = (dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1 ? _GEN_350 :
    _GEN_317; // @[scheduler.scala 334:90]
  wire [3:0] _bufferQueueUpdate_8_branchMask_T = bufferQueue_8_branchMask ^ branchOps_branchMask; // @[scheduler.scala 307:96]
  wire [3:0] _GEN_314 = _T_286 ? _bufferQueueUpdate_8_branchMask_T : bufferQueue_8_branchMask; // @[scheduler.scala 305:12 307:{58,77}]
  wire [3:0] bufferQueueUpdate_8_branchMask = branchOps_valid ? _GEN_314 : bufferQueue_8_branchMask; // @[scheduler.scala 305:12 306:28]
  wire  _T_339 = bufferQueue_0_valid | bufferQueue_1_valid | bufferQueue_2_valid | bufferQueue_3_valid |
    bufferQueue_4_valid | bufferQueue_5_valid | bufferQueue_6_valid | bufferQueue_7_valid | bufferQueue_8_valid; // @[scheduler.scala 339:50]
  wire [3:0] _T_291 = bufferQueue_9_branchMask & branchOps_branchMask; // @[scheduler.scala 308:50]
  wire  _T_292 = |_T_291; // @[scheduler.scala 308:74]
  wire  _GEN_319 = _T_80 & |_T_291 ? 1'h0 : bufferQueue_9_valid; // @[scheduler.scala 305:12 308:{79,94}]
  wire  _GEN_321 = branchOps_valid ? _GEN_319 : bufferQueue_9_valid; // @[scheduler.scala 305:12 306:28]
  wire  _GEN_351 = ~_T_339 & bufferQueue_9_valid ? 1'h0 : _GEN_321; // @[scheduler.scala 341:{107,92}]
  wire  bufferQueueUpdate_9_valid = (dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1 ? _GEN_351 :
    _GEN_321; // @[scheduler.scala 334:90]
  wire [3:0] _bufferQueueUpdate_9_branchMask_T = bufferQueue_9_branchMask ^ branchOps_branchMask; // @[scheduler.scala 307:96]
  wire [3:0] _GEN_318 = _T_292 ? _bufferQueueUpdate_9_branchMask_T : bufferQueue_9_branchMask; // @[scheduler.scala 305:12 307:{58,77}]
  wire [3:0] bufferQueueUpdate_9_branchMask = branchOps_valid ? _GEN_318 : bufferQueue_9_branchMask; // @[scheduler.scala 305:12 306:28]
  wire  _T_340 = bufferQueue_0_valid | bufferQueue_1_valid | bufferQueue_2_valid | bufferQueue_3_valid |
    bufferQueue_4_valid | bufferQueue_5_valid | bufferQueue_6_valid | bufferQueue_7_valid | bufferQueue_8_valid |
    bufferQueue_9_valid; // @[scheduler.scala 339:50]
  wire [3:0] _T_297 = bufferQueue_10_branchMask & branchOps_branchMask; // @[scheduler.scala 308:50]
  wire  _T_298 = |_T_297; // @[scheduler.scala 308:74]
  wire  _GEN_323 = _T_80 & |_T_297 ? 1'h0 : bufferQueue_10_valid; // @[scheduler.scala 305:12 308:{79,94}]
  wire  _GEN_325 = branchOps_valid ? _GEN_323 : bufferQueue_10_valid; // @[scheduler.scala 305:12 306:28]
  wire  _GEN_352 = ~_T_340 & bufferQueue_10_valid ? 1'h0 : _GEN_325; // @[scheduler.scala 341:{107,92}]
  wire  bufferQueueUpdate_10_valid = (dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1 ? _GEN_352 :
    _GEN_325; // @[scheduler.scala 334:90]
  wire [3:0] _bufferQueueUpdate_10_branchMask_T = bufferQueue_10_branchMask ^ branchOps_branchMask; // @[scheduler.scala 307:96]
  wire [3:0] _GEN_322 = _T_298 ? _bufferQueueUpdate_10_branchMask_T : bufferQueue_10_branchMask; // @[scheduler.scala 305:12 307:{58,77}]
  wire [3:0] bufferQueueUpdate_10_branchMask = branchOps_valid ? _GEN_322 : bufferQueue_10_branchMask; // @[scheduler.scala 305:12 306:28]
  wire  _T_341 = bufferQueue_0_valid | bufferQueue_1_valid | bufferQueue_2_valid | bufferQueue_3_valid |
    bufferQueue_4_valid | bufferQueue_5_valid | bufferQueue_6_valid | bufferQueue_7_valid | bufferQueue_8_valid |
    bufferQueue_9_valid | bufferQueue_10_valid; // @[scheduler.scala 339:50]
  wire [3:0] _T_303 = bufferQueue_11_branchMask & branchOps_branchMask; // @[scheduler.scala 308:50]
  wire  _T_304 = |_T_303; // @[scheduler.scala 308:74]
  wire  _GEN_327 = _T_80 & |_T_303 ? 1'h0 : bufferQueue_11_valid; // @[scheduler.scala 305:12 308:{79,94}]
  wire  _GEN_329 = branchOps_valid ? _GEN_327 : bufferQueue_11_valid; // @[scheduler.scala 305:12 306:28]
  wire  _GEN_353 = ~_T_341 & bufferQueue_11_valid ? 1'h0 : _GEN_329; // @[scheduler.scala 341:{107,92}]
  wire  bufferQueueUpdate_11_valid = (dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1 ? _GEN_353 :
    _GEN_329; // @[scheduler.scala 334:90]
  wire [3:0] _bufferQueueUpdate_11_branchMask_T = bufferQueue_11_branchMask ^ branchOps_branchMask; // @[scheduler.scala 307:96]
  wire [3:0] _GEN_326 = _T_304 ? _bufferQueueUpdate_11_branchMask_T : bufferQueue_11_branchMask; // @[scheduler.scala 305:12 307:{58,77}]
  wire [3:0] bufferQueueUpdate_11_branchMask = branchOps_valid ? _GEN_326 : bufferQueue_11_branchMask; // @[scheduler.scala 305:12 306:28]
  wire  _T_377 = _T_341 | bufferQueue_11_valid; // @[scheduler.scala 344:45]
  wire [3:0] _T_309 = newInstruction_branchMask & branchOps_branchMask; // @[scheduler.scala 308:50]
  wire  _T_310 = |_T_309; // @[scheduler.scala 308:74]
  wire  _GEN_331 = _T_80 & |_T_309 ? 1'h0 : newInstruction_valid; // @[scheduler.scala 305:12 308:{79,94}]
  wire  _GEN_333 = branchOps_valid ? _GEN_331 : newInstruction_valid; // @[scheduler.scala 305:12 306:28]
  wire  _GEN_354 = ~(_T_341 | bufferQueue_11_valid) ? 1'h0 : _GEN_333; // @[scheduler.scala 344:{52,98}]
  wire  bufferQueueUpdate_12_valid = (dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1 ? _GEN_354 :
    _GEN_333; // @[scheduler.scala 334:90]
  wire [3:0] _bufferQueueUpdate_12_branchMask_T = newInstruction_branchMask ^ branchOps_branchMask; // @[scheduler.scala 307:96]
  wire [3:0] _GEN_330 = _T_310 ? _bufferQueueUpdate_12_branchMask_T : newInstruction_branchMask; // @[scheduler.scala 305:12 307:{58,77}]
  wire [3:0] bufferQueueUpdate_12_branchMask = branchOps_valid ? _GEN_330 : newInstruction_branchMask; // @[scheduler.scala 305:12 306:28]
  wire  _GEN_334 = peripheral_ready ? 1'h0 : toPeripheral; // @[scheduler.scala 312:25 313:18 117:25]
  wire  _nextFrmBuffer_T_11_valid = bufferQueue_10_valid ? bufferQueue_10_valid : bufferQueue_11_valid; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_11_address = bufferQueue_10_valid ? bufferQueue_10_address : bufferQueue_11_address; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_11_instruction = bufferQueue_10_valid ? bufferQueue_10_instruction :
    bufferQueue_11_instruction; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_11_branchMask = bufferQueue_10_valid ? bufferQueue_10_branchMask :
    bufferQueue_11_branchMask; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_11_robAddr = bufferQueue_10_valid ? bufferQueue_10_robAddr : bufferQueue_11_robAddr; // @[Mux.scala 101:16]
  wire [5:0] _nextFrmBuffer_T_11_prfDest = bufferQueue_10_valid ? bufferQueue_10_prfDest : bufferQueue_11_prfDest; // @[Mux.scala 101:16]
  wire  _nextFrmBuffer_T_12_valid = bufferQueue_9_valid ? bufferQueue_9_valid : _nextFrmBuffer_T_11_valid; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_12_address = bufferQueue_9_valid ? bufferQueue_9_address : _nextFrmBuffer_T_11_address; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_12_instruction = bufferQueue_9_valid ? bufferQueue_9_instruction :
    _nextFrmBuffer_T_11_instruction; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_12_branchMask = bufferQueue_9_valid ? bufferQueue_9_branchMask :
    _nextFrmBuffer_T_11_branchMask; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_12_robAddr = bufferQueue_9_valid ? bufferQueue_9_robAddr : _nextFrmBuffer_T_11_robAddr; // @[Mux.scala 101:16]
  wire [5:0] _nextFrmBuffer_T_12_prfDest = bufferQueue_9_valid ? bufferQueue_9_prfDest : _nextFrmBuffer_T_11_prfDest; // @[Mux.scala 101:16]
  wire  _nextFrmBuffer_T_13_valid = bufferQueue_8_valid ? bufferQueue_8_valid : _nextFrmBuffer_T_12_valid; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_13_address = bufferQueue_8_valid ? bufferQueue_8_address : _nextFrmBuffer_T_12_address; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_13_instruction = bufferQueue_8_valid ? bufferQueue_8_instruction :
    _nextFrmBuffer_T_12_instruction; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_13_branchMask = bufferQueue_8_valid ? bufferQueue_8_branchMask :
    _nextFrmBuffer_T_12_branchMask; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_13_robAddr = bufferQueue_8_valid ? bufferQueue_8_robAddr : _nextFrmBuffer_T_12_robAddr; // @[Mux.scala 101:16]
  wire [5:0] _nextFrmBuffer_T_13_prfDest = bufferQueue_8_valid ? bufferQueue_8_prfDest : _nextFrmBuffer_T_12_prfDest; // @[Mux.scala 101:16]
  wire  _nextFrmBuffer_T_14_valid = bufferQueue_7_valid ? bufferQueue_7_valid : _nextFrmBuffer_T_13_valid; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_14_address = bufferQueue_7_valid ? bufferQueue_7_address : _nextFrmBuffer_T_13_address; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_14_instruction = bufferQueue_7_valid ? bufferQueue_7_instruction :
    _nextFrmBuffer_T_13_instruction; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_14_branchMask = bufferQueue_7_valid ? bufferQueue_7_branchMask :
    _nextFrmBuffer_T_13_branchMask; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_14_robAddr = bufferQueue_7_valid ? bufferQueue_7_robAddr : _nextFrmBuffer_T_13_robAddr; // @[Mux.scala 101:16]
  wire [5:0] _nextFrmBuffer_T_14_prfDest = bufferQueue_7_valid ? bufferQueue_7_prfDest : _nextFrmBuffer_T_13_prfDest; // @[Mux.scala 101:16]
  wire  _nextFrmBuffer_T_15_valid = bufferQueue_6_valid ? bufferQueue_6_valid : _nextFrmBuffer_T_14_valid; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_15_address = bufferQueue_6_valid ? bufferQueue_6_address : _nextFrmBuffer_T_14_address; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_15_instruction = bufferQueue_6_valid ? bufferQueue_6_instruction :
    _nextFrmBuffer_T_14_instruction; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_15_branchMask = bufferQueue_6_valid ? bufferQueue_6_branchMask :
    _nextFrmBuffer_T_14_branchMask; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_15_robAddr = bufferQueue_6_valid ? bufferQueue_6_robAddr : _nextFrmBuffer_T_14_robAddr; // @[Mux.scala 101:16]
  wire [5:0] _nextFrmBuffer_T_15_prfDest = bufferQueue_6_valid ? bufferQueue_6_prfDest : _nextFrmBuffer_T_14_prfDest; // @[Mux.scala 101:16]
  wire  _nextFrmBuffer_T_16_valid = bufferQueue_5_valid ? bufferQueue_5_valid : _nextFrmBuffer_T_15_valid; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_16_address = bufferQueue_5_valid ? bufferQueue_5_address : _nextFrmBuffer_T_15_address; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_16_instruction = bufferQueue_5_valid ? bufferQueue_5_instruction :
    _nextFrmBuffer_T_15_instruction; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_16_branchMask = bufferQueue_5_valid ? bufferQueue_5_branchMask :
    _nextFrmBuffer_T_15_branchMask; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_16_robAddr = bufferQueue_5_valid ? bufferQueue_5_robAddr : _nextFrmBuffer_T_15_robAddr; // @[Mux.scala 101:16]
  wire [5:0] _nextFrmBuffer_T_16_prfDest = bufferQueue_5_valid ? bufferQueue_5_prfDest : _nextFrmBuffer_T_15_prfDest; // @[Mux.scala 101:16]
  wire  _nextFrmBuffer_T_17_valid = bufferQueue_4_valid ? bufferQueue_4_valid : _nextFrmBuffer_T_16_valid; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_17_address = bufferQueue_4_valid ? bufferQueue_4_address : _nextFrmBuffer_T_16_address; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_17_instruction = bufferQueue_4_valid ? bufferQueue_4_instruction :
    _nextFrmBuffer_T_16_instruction; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_17_branchMask = bufferQueue_4_valid ? bufferQueue_4_branchMask :
    _nextFrmBuffer_T_16_branchMask; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_17_robAddr = bufferQueue_4_valid ? bufferQueue_4_robAddr : _nextFrmBuffer_T_16_robAddr; // @[Mux.scala 101:16]
  wire [5:0] _nextFrmBuffer_T_17_prfDest = bufferQueue_4_valid ? bufferQueue_4_prfDest : _nextFrmBuffer_T_16_prfDest; // @[Mux.scala 101:16]
  wire  _nextFrmBuffer_T_18_valid = bufferQueue_3_valid ? bufferQueue_3_valid : _nextFrmBuffer_T_17_valid; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_18_address = bufferQueue_3_valid ? bufferQueue_3_address : _nextFrmBuffer_T_17_address; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_18_instruction = bufferQueue_3_valid ? bufferQueue_3_instruction :
    _nextFrmBuffer_T_17_instruction; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_18_branchMask = bufferQueue_3_valid ? bufferQueue_3_branchMask :
    _nextFrmBuffer_T_17_branchMask; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_18_robAddr = bufferQueue_3_valid ? bufferQueue_3_robAddr : _nextFrmBuffer_T_17_robAddr; // @[Mux.scala 101:16]
  wire [5:0] _nextFrmBuffer_T_18_prfDest = bufferQueue_3_valid ? bufferQueue_3_prfDest : _nextFrmBuffer_T_17_prfDest; // @[Mux.scala 101:16]
  wire  _nextFrmBuffer_T_19_valid = bufferQueue_2_valid ? bufferQueue_2_valid : _nextFrmBuffer_T_18_valid; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_19_address = bufferQueue_2_valid ? bufferQueue_2_address : _nextFrmBuffer_T_18_address; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_19_instruction = bufferQueue_2_valid ? bufferQueue_2_instruction :
    _nextFrmBuffer_T_18_instruction; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_19_branchMask = bufferQueue_2_valid ? bufferQueue_2_branchMask :
    _nextFrmBuffer_T_18_branchMask; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_19_robAddr = bufferQueue_2_valid ? bufferQueue_2_robAddr : _nextFrmBuffer_T_18_robAddr; // @[Mux.scala 101:16]
  wire [5:0] _nextFrmBuffer_T_19_prfDest = bufferQueue_2_valid ? bufferQueue_2_prfDest : _nextFrmBuffer_T_18_prfDest; // @[Mux.scala 101:16]
  wire  _nextFrmBuffer_T_20_valid = bufferQueue_1_valid ? bufferQueue_1_valid : _nextFrmBuffer_T_19_valid; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_20_address = bufferQueue_1_valid ? bufferQueue_1_address : _nextFrmBuffer_T_19_address; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_20_instruction = bufferQueue_1_valid ? bufferQueue_1_instruction :
    _nextFrmBuffer_T_19_instruction; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_20_branchMask = bufferQueue_1_valid ? bufferQueue_1_branchMask :
    _nextFrmBuffer_T_19_branchMask; // @[Mux.scala 101:16]
  wire  _nextFrmBuffer_T_21_valid = bufferQueue_0_valid ? bufferQueue_0_valid : _nextFrmBuffer_T_20_valid; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_21_address = bufferQueue_0_valid ? bufferQueue_0_address : _nextFrmBuffer_T_20_address; // @[Mux.scala 101:16]
  wire [31:0] _nextFrmBuffer_T_21_instruction = bufferQueue_0_valid ? bufferQueue_0_instruction :
    _nextFrmBuffer_T_20_instruction; // @[Mux.scala 101:16]
  wire [3:0] _nextFrmBuffer_T_21_branchMask = bufferQueue_0_valid ? bufferQueue_0_branchMask :
    _nextFrmBuffer_T_20_branchMask; // @[Mux.scala 101:16]
  wire  nextFrmBuffer_valid = _T_377 ? _nextFrmBuffer_T_21_valid : newInstruction_valid; // @[scheduler.scala 315:26]
  wire [31:0] nextFrmBuffer_address = _T_377 ? _nextFrmBuffer_T_21_address : newInstruction_address; // @[scheduler.scala 315:26]
  wire [31:0] nextFrmBuffer_instruction = _T_377 ? _nextFrmBuffer_T_21_instruction : newInstruction_instruction; // @[scheduler.scala 315:26]
  wire [3:0] nextFrmBuffer_branchMask = _T_377 ? _nextFrmBuffer_T_21_branchMask : newInstruction_branchMask; // @[scheduler.scala 315:26]
  wire  _T_323 = nextFrmBuffer_address >= 32'h80000000; // @[configuration.scala 41:44]
  wire  _T_326 = ~_T_323; // @[scheduler.scala 336:10]
  wire  _GEN_341 = ~_T_323 & ~nextFrmBuffer_instruction[5] ? 1'h0 : nextFrmBuffer_valid; // @[scheduler.scala 336:{100,119} 335:16]
  wire [3:0] _T_379 = branchOps_branchMask & nextFrmBuffer_branchMask; // @[scheduler.scala 349:34]
  wire  _T_380 = |_T_379; // @[scheduler.scala 349:62]
  wire [3:0] _fromBuffer_branchMask_T_1 = branchOps_branchMask ^ nextFrmBuffer_branchMask; // @[scheduler.scala 349:114]
  assign toCache_queryWithData_query_valid = scheduledInstruction_query_valid; // @[scheduler.scala 60:25]
  assign toCache_queryWithData_query_address = scheduledInstruction_query_address; // @[scheduler.scala 60:25]
  assign toCache_queryWithData_query_instruction = scheduledInstruction_query_instruction; // @[scheduler.scala 60:25]
  assign toCache_queryWithData_query_branchMask = scheduledInstruction_query_branchMask; // @[scheduler.scala 60:25]
  assign toCache_queryWithData_query_robAddr = scheduledInstruction_query_robAddr; // @[scheduler.scala 60:25]
  assign toCache_queryWithData_query_prfDest = scheduledInstruction_query_prfDest; // @[scheduler.scala 60:25]
  assign toCache_queryWithData_data = scheduledInstruction_data; // @[scheduler.scala 60:25]
  assign toCache_replaying = toCache_replaying_REG; // @[scheduler.scala 92:21]
  assign storeCommit_ready = storeInstructions_0_valid; // @[scheduler.scala 84:21]
  assign peripheral_bits_valid = toPeripheral; // @[scheduler.scala 358:25]
  assign peripheral_bits_address = fromBuffer_address; // @[scheduler.scala 357:19]
  assign peripheral_bits_instruction = fromBuffer_instruction; // @[scheduler.scala 357:19]
  assign peripheral_bits_branchMask = fromBuffer_branchMask; // @[scheduler.scala 357:19]
  assign peripheral_bits_robAddr = fromBuffer_robAddr; // @[scheduler.scala 357:19]
  assign peripheral_bits_prfDest = fromBuffer_prfDest; // @[scheduler.scala 357:19]
  assign canAllocate = ~(bufferQueue_7_valid | bufferQueue_6_valid | bufferQueue_5_valid | bufferQueue_4_valid |
    bufferQueue_3_valid | bufferQueue_2_valid | bufferQueue_1_valid | bufferQueue_0_valid); // @[scheduler.scala 363:18]
  assign clean = ~(_T_377 | dependentReads_0_valid | dependentReads_1_valid | dependentReads_2_valid |
    dependentReads_3_valid | storeInstructions_0_valid | storeInstructions_1_valid | storeInstructions_2_valid |
    storeInstructions_3_valid | fromBuffer_valid); // @[scheduler.scala 367:12]
  always @(posedge clock) begin
    if (reset) begin // @[scheduler.scala 52:37]
      scheduledInstruction_query_valid <= 1'h0; // @[scheduler.scala 52:37]
    end else if (branchOps_valid) begin // @[scheduler.scala 165:25]
      if (_T_80 & _T_7) begin // @[scheduler.scala 169:92]
        scheduledInstruction_query_valid <= 1'h0; // @[scheduler.scala 169:127]
      end else begin
        scheduledInstruction_query_valid <= _GEN_6;
      end
    end else begin
      scheduledInstruction_query_valid <= _GEN_6;
    end
    if (replaying | ~cacheStalled) begin // @[scheduler.scala 163:38]
      if (replaying) begin // @[scheduler.scala 270:19]
        scheduledInstruction_query_address <= replayQueue_query_address; // @[scheduler.scala 270:35]
      end else if (storeCommit_fired) begin // @[scheduler.scala 271:32]
        if (storeInstructions_0_valid) begin // @[Mux.scala 101:16]
          scheduledInstruction_query_address <= storeInstructions_0_address;
        end else begin
          scheduledInstruction_query_address <= _storeInstruction_T_2_address;
        end
      end else if (_readCanDequeue_T_4) begin // @[scheduler.scala 272:67]
        scheduledInstruction_query_address <= dependentRead_address; // @[scheduler.scala 273:33]
      end else begin
        scheduledInstruction_query_address <= fromBuffer_address; // @[scheduler.scala 281:25]
      end
    end
    if (replaying | ~cacheStalled) begin // @[scheduler.scala 163:38]
      if (replaying) begin // @[scheduler.scala 270:19]
        scheduledInstruction_query_instruction <= replayQueue_query_instruction; // @[scheduler.scala 270:35]
      end else if (storeCommit_fired) begin // @[scheduler.scala 271:32]
        if (storeInstructions_0_valid) begin // @[Mux.scala 101:16]
          scheduledInstruction_query_instruction <= storeInstructions_0_instruction;
        end else begin
          scheduledInstruction_query_instruction <= _storeInstruction_T_2_instruction;
        end
      end else if (_readCanDequeue_T_4) begin // @[scheduler.scala 272:67]
        scheduledInstruction_query_instruction <= dependentRead_instruction; // @[scheduler.scala 275:37]
      end else begin
        scheduledInstruction_query_instruction <= _GEN_190;
      end
    end
    if (branchOps_valid) begin // @[scheduler.scala 165:25]
      if (|_T_6) begin // @[scheduler.scala 166:70]
        scheduledInstruction_query_branchMask <= _scheduledInstruction_query_branchMask_T; // @[scheduler.scala 167:45]
      end else begin
        scheduledInstruction_query_branchMask <= _GEN_9;
      end
    end else begin
      scheduledInstruction_query_branchMask <= _GEN_9;
    end
    if (replaying | ~cacheStalled) begin // @[scheduler.scala 163:38]
      if (replaying) begin // @[scheduler.scala 270:19]
        scheduledInstruction_query_robAddr <= replayQueue_query_robAddr; // @[scheduler.scala 270:35]
      end else if (storeCommit_fired) begin // @[scheduler.scala 271:32]
        if (storeInstructions_0_valid) begin // @[Mux.scala 101:16]
          scheduledInstruction_query_robAddr <= storeInstructions_0_robAddr;
        end else begin
          scheduledInstruction_query_robAddr <= _storeInstruction_T_2_robAddr;
        end
      end else if (_readCanDequeue_T_4) begin // @[scheduler.scala 272:67]
        scheduledInstruction_query_robAddr <= dependentRead_robAddr; // @[scheduler.scala 277:33]
      end else begin
        scheduledInstruction_query_robAddr <= fromBuffer_robAddr; // @[scheduler.scala 281:25]
      end
    end
    if (replaying | ~cacheStalled) begin // @[scheduler.scala 163:38]
      if (replaying) begin // @[scheduler.scala 270:19]
        scheduledInstruction_query_prfDest <= replayQueue_query_prfDest; // @[scheduler.scala 270:35]
      end else if (storeCommit_fired) begin // @[scheduler.scala 271:32]
        if (storeInstructions_0_valid) begin // @[Mux.scala 101:16]
          scheduledInstruction_query_prfDest <= storeInstructions_0_prfDest;
        end else begin
          scheduledInstruction_query_prfDest <= _storeInstruction_T_2_prfDest;
        end
      end else if (_readCanDequeue_T_4) begin // @[scheduler.scala 272:67]
        scheduledInstruction_query_prfDest <= dependentRead_prfDest; // @[scheduler.scala 276:33]
      end else begin
        scheduledInstruction_query_prfDest <= fromBuffer_prfDest; // @[scheduler.scala 281:25]
      end
    end
    if (replaying | ~cacheStalled) begin // @[scheduler.scala 163:38]
      scheduledInstruction_data <= replayQueue_data; // @[scheduler.scala 163:61]
    end
    if (reset) begin // @[scheduler.scala 65:31]
      dependentReads_0_valid <= 1'h0; // @[scheduler.scala 65:31]
    end else if (~dependentReads_0_valid) begin // @[scheduler.scala 263:47]
      dependentReads_0_valid <= dependentReadsUpdate_1_valid; // @[scheduler.scala 263:53]
    end else if (dependentReads_0_dependency_free & dependentReads_0_valid & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_0_valid <= dependentReadsUpdate_1_valid; // @[scheduler.scala 266:11]
    end else if (~replaying & _T_4 & ~storeCommit_fired & dependentRead_valid & dependentRead_dependency_free) begin // @[scheduler.scala 252:115]
      dependentReads_0_valid <= _GEN_117;
    end else begin
      dependentReads_0_valid <= _GEN_90;
    end
    if (~dependentReads_0_valid) begin // @[scheduler.scala 263:47]
      dependentReads_0_address <= dependentReads_1_address; // @[scheduler.scala 263:53]
    end else if (dependentReads_0_dependency_free & dependentReads_0_valid & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_0_address <= dependentReads_1_address; // @[scheduler.scala 266:11]
    end
    if (~dependentReads_0_valid) begin // @[scheduler.scala 263:47]
      dependentReads_0_instruction <= dependentReads_1_instruction; // @[scheduler.scala 263:53]
    end else if (dependentReads_0_dependency_free & dependentReads_0_valid & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_0_instruction <= dependentReads_1_instruction; // @[scheduler.scala 266:11]
    end
    if (~dependentReads_0_valid) begin // @[scheduler.scala 263:47]
      dependentReads_0_branchMask <= dependentReadsUpdate_1_branchMask; // @[scheduler.scala 263:53]
    end else if (dependentReads_0_dependency_free & dependentReads_0_valid & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_0_branchMask <= dependentReadsUpdate_1_branchMask; // @[scheduler.scala 266:11]
    end else if (branchOps_valid) begin // @[scheduler.scala 239:27]
      if (|_T_50) begin // @[scheduler.scala 240:58]
        dependentReads_0_branchMask <= _dependentReadsUpdate_0_branchMask_T; // @[scheduler.scala 241:25]
      end
    end
    if (~dependentReads_0_valid) begin // @[scheduler.scala 263:47]
      dependentReads_0_robAddr <= dependentReads_1_robAddr; // @[scheduler.scala 263:53]
    end else if (dependentReads_0_dependency_free & dependentReads_0_valid & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_0_robAddr <= dependentReads_1_robAddr; // @[scheduler.scala 266:11]
    end
    if (~dependentReads_0_valid) begin // @[scheduler.scala 263:47]
      dependentReads_0_prfDest <= dependentReads_1_prfDest; // @[scheduler.scala 263:53]
    end else if (dependentReads_0_dependency_free & dependentReads_0_valid & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_0_prfDest <= dependentReads_1_prfDest; // @[scheduler.scala 266:11]
    end
    if (~dependentReads_0_valid) begin // @[scheduler.scala 263:47]
      dependentReads_0_dependency_free <= dependentReadsUpdate_1_dependency_free; // @[scheduler.scala 263:53]
    end else if (dependentReads_0_dependency_free & dependentReads_0_valid & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_0_dependency_free <= dependentReadsUpdate_1_dependency_free; // @[scheduler.scala 266:11]
    end else if (REG) begin // @[scheduler.scala 245:38]
      dependentReads_0_dependency_free <= _GEN_91;
    end
    if (~dependentReads_0_valid) begin // @[scheduler.scala 263:47]
      dependentReads_0_dependency_robAddr <= dependentReads_1_dependency_robAddr; // @[scheduler.scala 263:53]
    end else if (dependentReads_0_dependency_free & dependentReads_0_valid & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_0_dependency_robAddr <= dependentReads_1_dependency_robAddr; // @[scheduler.scala 266:11]
    end
    if (reset) begin // @[scheduler.scala 65:31]
      dependentReads_1_valid <= 1'h0; // @[scheduler.scala 65:31]
    end else if (~dependentReads_0_valid | ~dependentReads_1_valid) begin // @[scheduler.scala 263:47]
      dependentReads_1_valid <= dependentReadsUpdate_2_valid; // @[scheduler.scala 263:53]
    end else if ((_T_92 | dependentReads_1_dependency_free & dependentReads_1_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_1_valid <= dependentReadsUpdate_2_valid; // @[scheduler.scala 266:11]
    end else if (~replaying & _T_4 & ~storeCommit_fired & dependentRead_valid & dependentRead_dependency_free) begin // @[scheduler.scala 252:115]
      dependentReads_1_valid <= _GEN_118;
    end else begin
      dependentReads_1_valid <= _GEN_96;
    end
    if (~dependentReads_0_valid | ~dependentReads_1_valid) begin // @[scheduler.scala 263:47]
      dependentReads_1_address <= dependentReads_2_address; // @[scheduler.scala 263:53]
    end else if ((_T_92 | dependentReads_1_dependency_free & dependentReads_1_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_1_address <= dependentReads_2_address; // @[scheduler.scala 266:11]
    end
    if (~dependentReads_0_valid | ~dependentReads_1_valid) begin // @[scheduler.scala 263:47]
      dependentReads_1_instruction <= dependentReads_2_instruction; // @[scheduler.scala 263:53]
    end else if ((_T_92 | dependentReads_1_dependency_free & dependentReads_1_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_1_instruction <= dependentReads_2_instruction; // @[scheduler.scala 266:11]
    end
    if (~dependentReads_0_valid | ~dependentReads_1_valid) begin // @[scheduler.scala 263:47]
      dependentReads_1_branchMask <= dependentReadsUpdate_2_branchMask; // @[scheduler.scala 263:53]
    end else if ((_T_92 | dependentReads_1_dependency_free & dependentReads_1_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_1_branchMask <= dependentReadsUpdate_2_branchMask; // @[scheduler.scala 266:11]
    end else if (branchOps_valid) begin // @[scheduler.scala 239:27]
      if (|_T_57) begin // @[scheduler.scala 240:58]
        dependentReads_1_branchMask <= _dependentReadsUpdate_1_branchMask_T; // @[scheduler.scala 241:25]
      end
    end
    if (~dependentReads_0_valid | ~dependentReads_1_valid) begin // @[scheduler.scala 263:47]
      dependentReads_1_robAddr <= dependentReads_2_robAddr; // @[scheduler.scala 263:53]
    end else if ((_T_92 | dependentReads_1_dependency_free & dependentReads_1_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_1_robAddr <= dependentReads_2_robAddr; // @[scheduler.scala 266:11]
    end
    if (~dependentReads_0_valid | ~dependentReads_1_valid) begin // @[scheduler.scala 263:47]
      dependentReads_1_prfDest <= dependentReads_2_prfDest; // @[scheduler.scala 263:53]
    end else if ((_T_92 | dependentReads_1_dependency_free & dependentReads_1_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_1_prfDest <= dependentReads_2_prfDest; // @[scheduler.scala 266:11]
    end
    if (~dependentReads_0_valid | ~dependentReads_1_valid) begin // @[scheduler.scala 263:47]
      dependentReads_1_dependency_free <= dependentReadsUpdate_2_dependency_free; // @[scheduler.scala 263:53]
    end else if ((_T_92 | dependentReads_1_dependency_free & dependentReads_1_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_1_dependency_free <= dependentReadsUpdate_2_dependency_free; // @[scheduler.scala 266:11]
    end else if (REG_1) begin // @[scheduler.scala 245:38]
      dependentReads_1_dependency_free <= _GEN_97;
    end
    if (~dependentReads_0_valid | ~dependentReads_1_valid) begin // @[scheduler.scala 263:47]
      dependentReads_1_dependency_robAddr <= dependentReads_2_dependency_robAddr; // @[scheduler.scala 263:53]
    end else if ((_T_92 | dependentReads_1_dependency_free & dependentReads_1_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_1_dependency_robAddr <= dependentReads_2_dependency_robAddr; // @[scheduler.scala 266:11]
    end
    if (reset) begin // @[scheduler.scala 65:31]
      dependentReads_2_valid <= 1'h0; // @[scheduler.scala 65:31]
    end else if (~_readCanDequeue_T | ~dependentReads_2_valid) begin // @[scheduler.scala 263:47]
      dependentReads_2_valid <= dependentReadsUpdate_3_valid; // @[scheduler.scala 263:53]
    end else if ((_T_97 | dependentReads_2_dependency_free & dependentReads_2_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_2_valid <= dependentReadsUpdate_3_valid; // @[scheduler.scala 266:11]
    end else if (~replaying & _T_4 & ~storeCommit_fired & dependentRead_valid & dependentRead_dependency_free) begin // @[scheduler.scala 252:115]
      dependentReads_2_valid <= _GEN_119;
    end else begin
      dependentReads_2_valid <= _GEN_102;
    end
    if (~_readCanDequeue_T | ~dependentReads_2_valid) begin // @[scheduler.scala 263:47]
      dependentReads_2_address <= dependentReads_3_address; // @[scheduler.scala 263:53]
    end else if ((_T_97 | dependentReads_2_dependency_free & dependentReads_2_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_2_address <= dependentReads_3_address; // @[scheduler.scala 266:11]
    end
    if (~_readCanDequeue_T | ~dependentReads_2_valid) begin // @[scheduler.scala 263:47]
      dependentReads_2_instruction <= dependentReads_3_instruction; // @[scheduler.scala 263:53]
    end else if ((_T_97 | dependentReads_2_dependency_free & dependentReads_2_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_2_instruction <= dependentReads_3_instruction; // @[scheduler.scala 266:11]
    end
    if (~_readCanDequeue_T | ~dependentReads_2_valid) begin // @[scheduler.scala 263:47]
      dependentReads_2_branchMask <= dependentReadsUpdate_3_branchMask; // @[scheduler.scala 263:53]
    end else if ((_T_97 | dependentReads_2_dependency_free & dependentReads_2_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_2_branchMask <= dependentReadsUpdate_3_branchMask; // @[scheduler.scala 266:11]
    end else if (branchOps_valid) begin // @[scheduler.scala 239:27]
      if (|_T_64) begin // @[scheduler.scala 240:58]
        dependentReads_2_branchMask <= _dependentReadsUpdate_2_branchMask_T; // @[scheduler.scala 241:25]
      end
    end
    if (~_readCanDequeue_T | ~dependentReads_2_valid) begin // @[scheduler.scala 263:47]
      dependentReads_2_robAddr <= dependentReads_3_robAddr; // @[scheduler.scala 263:53]
    end else if ((_T_97 | dependentReads_2_dependency_free & dependentReads_2_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_2_robAddr <= dependentReads_3_robAddr; // @[scheduler.scala 266:11]
    end
    if (~_readCanDequeue_T | ~dependentReads_2_valid) begin // @[scheduler.scala 263:47]
      dependentReads_2_prfDest <= dependentReads_3_prfDest; // @[scheduler.scala 263:53]
    end else if ((_T_97 | dependentReads_2_dependency_free & dependentReads_2_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_2_prfDest <= dependentReads_3_prfDest; // @[scheduler.scala 266:11]
    end
    if (~_readCanDequeue_T | ~dependentReads_2_valid) begin // @[scheduler.scala 263:47]
      dependentReads_2_dependency_free <= dependentReadsUpdate_3_dependency_free; // @[scheduler.scala 263:53]
    end else if ((_T_97 | dependentReads_2_dependency_free & dependentReads_2_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_2_dependency_free <= dependentReadsUpdate_3_dependency_free; // @[scheduler.scala 266:11]
    end else if (REG_2) begin // @[scheduler.scala 245:38]
      dependentReads_2_dependency_free <= _GEN_103;
    end
    if (~_readCanDequeue_T | ~dependentReads_2_valid) begin // @[scheduler.scala 263:47]
      dependentReads_2_dependency_robAddr <= dependentReads_3_dependency_robAddr; // @[scheduler.scala 263:53]
    end else if ((_T_97 | dependentReads_2_dependency_free & dependentReads_2_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_2_dependency_robAddr <= dependentReads_3_dependency_robAddr; // @[scheduler.scala 266:11]
    end
    if (reset) begin // @[scheduler.scala 65:31]
      dependentReads_3_valid <= 1'h0; // @[scheduler.scala 65:31]
    end else if (~_readCanDequeue_T_1 | ~dependentReads_3_valid) begin // @[scheduler.scala 263:47]
      dependentReads_3_valid <= dependentReadsUpdate_4_valid; // @[scheduler.scala 263:53]
    end else if ((_T_98 | dependentReads_3_dependency_free & dependentReads_3_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_3_valid <= dependentReadsUpdate_4_valid; // @[scheduler.scala 266:11]
    end else if (~replaying & _T_4 & ~storeCommit_fired & dependentRead_valid & dependentRead_dependency_free) begin // @[scheduler.scala 252:115]
      dependentReads_3_valid <= _GEN_120;
    end else begin
      dependentReads_3_valid <= _GEN_108;
    end
    if (~_readCanDequeue_T_1 | ~dependentReads_3_valid) begin // @[scheduler.scala 263:47]
      dependentReads_3_address <= fromBuffer_address; // @[scheduler.scala 263:53]
    end else if ((_T_98 | dependentReads_3_dependency_free & dependentReads_3_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_3_address <= fromBuffer_address; // @[scheduler.scala 266:11]
    end
    if (~_readCanDequeue_T_1 | ~dependentReads_3_valid) begin // @[scheduler.scala 263:47]
      dependentReads_3_instruction <= _GEN_190; // @[scheduler.scala 263:53]
    end else if ((_T_98 | dependentReads_3_dependency_free & dependentReads_3_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_3_instruction <= _GEN_190; // @[scheduler.scala 266:11]
    end
    if (~_readCanDequeue_T_1 | ~dependentReads_3_valid) begin // @[scheduler.scala 263:47]
      dependentReads_3_branchMask <= storeInstructionsUpdate_4_branchMask; // @[scheduler.scala 263:53]
    end else if ((_T_98 | dependentReads_3_dependency_free & dependentReads_3_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_3_branchMask <= storeInstructionsUpdate_4_branchMask; // @[scheduler.scala 266:11]
    end else if (branchOps_valid) begin // @[scheduler.scala 239:27]
      if (|_T_71) begin // @[scheduler.scala 240:58]
        dependentReads_3_branchMask <= _dependentReadsUpdate_3_branchMask_T; // @[scheduler.scala 241:25]
      end
    end
    if (~_readCanDequeue_T_1 | ~dependentReads_3_valid) begin // @[scheduler.scala 263:47]
      dependentReads_3_robAddr <= fromBuffer_robAddr; // @[scheduler.scala 263:53]
    end else if ((_T_98 | dependentReads_3_dependency_free & dependentReads_3_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_3_robAddr <= fromBuffer_robAddr; // @[scheduler.scala 266:11]
    end
    if (~_readCanDequeue_T_1 | ~dependentReads_3_valid) begin // @[scheduler.scala 263:47]
      dependentReads_3_prfDest <= fromBuffer_prfDest; // @[scheduler.scala 263:53]
    end else if ((_T_98 | dependentReads_3_dependency_free & dependentReads_3_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_3_prfDest <= fromBuffer_prfDest; // @[scheduler.scala 266:11]
    end
    if (~_readCanDequeue_T_1 | ~dependentReads_3_valid) begin // @[scheduler.scala 263:47]
      dependentReads_3_dependency_free <= dependentReadsUpdate_4_dependency_free; // @[scheduler.scala 263:53]
    end else if ((_T_98 | dependentReads_3_dependency_free & dependentReads_3_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_3_dependency_free <= dependentReadsUpdate_4_dependency_free; // @[scheduler.scala 266:11]
    end else if (REG_3) begin // @[scheduler.scala 245:38]
      dependentReads_3_dependency_free <= _GEN_109;
    end
    if (~_readCanDequeue_T_1 | ~dependentReads_3_valid) begin // @[scheduler.scala 263:47]
      dependentReads_3_dependency_robAddr <= currDependentReads_4_dependency_robAddr; // @[scheduler.scala 263:53]
    end else if ((_T_98 | dependentReads_3_dependency_free & dependentReads_3_valid) & _T_91) begin // @[scheduler.scala 264:186]
      dependentReads_3_dependency_robAddr <= currDependentReads_4_dependency_robAddr; // @[scheduler.scala 266:11]
    end
    if (reset) begin // @[scheduler.scala 76:34]
      storeInstructions_0_valid <= 1'h0; // @[scheduler.scala 76:34]
    end else if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_0_valid <= storeInstructionsUpdate_1_valid; // @[scheduler.scala 201:91]
    end else if (storeInstructions_0_valid) begin // @[scheduler.scala 197:96]
      if (storeCommit_fired) begin // @[scheduler.scala 189:27]
        storeInstructions_0_valid <= 1'h0; // @[scheduler.scala 190:40]
      end else begin
        storeInstructions_0_valid <= _GEN_20;
      end
    end else begin
      storeInstructions_0_valid <= storeInstructionsUpdate_1_valid; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_0_address <= storeInstructions_1_address; // @[scheduler.scala 201:91]
    end else if (!(storeInstructions_0_valid)) begin // @[scheduler.scala 197:96]
      storeInstructions_0_address <= storeInstructions_1_address; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_0_instruction <= storeInstructions_1_instruction; // @[scheduler.scala 201:91]
    end else if (!(storeInstructions_0_valid)) begin // @[scheduler.scala 197:96]
      storeInstructions_0_instruction <= storeInstructions_1_instruction; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_0_branchMask <= storeInstructionsUpdate_1_branchMask; // @[scheduler.scala 201:91]
    end else if (storeInstructions_0_valid) begin // @[scheduler.scala 197:96]
      if (branchOps_valid) begin // @[scheduler.scala 177:27]
        if (|_T_12) begin // @[scheduler.scala 178:59]
          storeInstructions_0_branchMask <= _storeInstructionsUpdate_0_branchMask_T; // @[scheduler.scala 178:77]
        end
      end
    end else begin
      storeInstructions_0_branchMask <= storeInstructionsUpdate_1_branchMask; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_0_robAddr <= storeInstructions_1_robAddr; // @[scheduler.scala 201:91]
    end else if (!(storeInstructions_0_valid)) begin // @[scheduler.scala 197:96]
      storeInstructions_0_robAddr <= storeInstructions_1_robAddr; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_0_prfDest <= storeInstructions_1_prfDest; // @[scheduler.scala 201:91]
    end else if (!(storeInstructions_0_valid)) begin // @[scheduler.scala 197:96]
      storeInstructions_0_prfDest <= storeInstructions_1_prfDest; // @[scheduler.scala 197:127]
    end
    if (reset) begin // @[scheduler.scala 76:34]
      storeInstructions_1_valid <= 1'h0; // @[scheduler.scala 76:34]
    end else if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_1_valid <= storeInstructionsUpdate_2_valid; // @[scheduler.scala 201:91]
    end else if (_storeInstructionsFree_T) begin // @[scheduler.scala 197:96]
      if (branchOps_valid) begin // @[scheduler.scala 177:27]
        storeInstructions_1_valid <= _GEN_22;
      end
    end else begin
      storeInstructions_1_valid <= storeInstructionsUpdate_2_valid; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_1_address <= storeInstructions_2_address; // @[scheduler.scala 201:91]
    end else if (!(_storeInstructionsFree_T)) begin // @[scheduler.scala 197:96]
      storeInstructions_1_address <= storeInstructions_2_address; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_1_instruction <= storeInstructions_2_instruction; // @[scheduler.scala 201:91]
    end else if (!(_storeInstructionsFree_T)) begin // @[scheduler.scala 197:96]
      storeInstructions_1_instruction <= storeInstructions_2_instruction; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_1_branchMask <= storeInstructionsUpdate_2_branchMask; // @[scheduler.scala 201:91]
    end else if (_storeInstructionsFree_T) begin // @[scheduler.scala 197:96]
      if (branchOps_valid) begin // @[scheduler.scala 177:27]
        if (|_T_18) begin // @[scheduler.scala 178:59]
          storeInstructions_1_branchMask <= _storeInstructionsUpdate_1_branchMask_T; // @[scheduler.scala 178:77]
        end
      end
    end else begin
      storeInstructions_1_branchMask <= storeInstructionsUpdate_2_branchMask; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_1_robAddr <= storeInstructions_2_robAddr; // @[scheduler.scala 201:91]
    end else if (!(_storeInstructionsFree_T)) begin // @[scheduler.scala 197:96]
      storeInstructions_1_robAddr <= storeInstructions_2_robAddr; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_1_prfDest <= storeInstructions_2_prfDest; // @[scheduler.scala 201:91]
    end else if (!(_storeInstructionsFree_T)) begin // @[scheduler.scala 197:96]
      storeInstructions_1_prfDest <= storeInstructions_2_prfDest; // @[scheduler.scala 197:127]
    end
    if (reset) begin // @[scheduler.scala 76:34]
      storeInstructions_2_valid <= 1'h0; // @[scheduler.scala 76:34]
    end else if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_2_valid <= storeInstructionsUpdate_3_valid; // @[scheduler.scala 201:91]
    end else if (_storeInstructionsFree_T_1) begin // @[scheduler.scala 197:96]
      if (branchOps_valid) begin // @[scheduler.scala 177:27]
        storeInstructions_2_valid <= _GEN_26;
      end
    end else begin
      storeInstructions_2_valid <= storeInstructionsUpdate_3_valid; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_2_address <= storeInstructions_3_address; // @[scheduler.scala 201:91]
    end else if (!(_storeInstructionsFree_T_1)) begin // @[scheduler.scala 197:96]
      storeInstructions_2_address <= storeInstructions_3_address; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_2_instruction <= storeInstructions_3_instruction; // @[scheduler.scala 201:91]
    end else if (!(_storeInstructionsFree_T_1)) begin // @[scheduler.scala 197:96]
      storeInstructions_2_instruction <= storeInstructions_3_instruction; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_2_branchMask <= storeInstructionsUpdate_3_branchMask; // @[scheduler.scala 201:91]
    end else if (_storeInstructionsFree_T_1) begin // @[scheduler.scala 197:96]
      if (branchOps_valid) begin // @[scheduler.scala 177:27]
        if (|_T_24) begin // @[scheduler.scala 178:59]
          storeInstructions_2_branchMask <= _storeInstructionsUpdate_2_branchMask_T; // @[scheduler.scala 178:77]
        end
      end
    end else begin
      storeInstructions_2_branchMask <= storeInstructionsUpdate_3_branchMask; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_2_robAddr <= storeInstructions_3_robAddr; // @[scheduler.scala 201:91]
    end else if (!(_storeInstructionsFree_T_1)) begin // @[scheduler.scala 197:96]
      storeInstructions_2_robAddr <= storeInstructions_3_robAddr; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_2_prfDest <= storeInstructions_3_prfDest; // @[scheduler.scala 201:91]
    end else if (!(_storeInstructionsFree_T_1)) begin // @[scheduler.scala 197:96]
      storeInstructions_2_prfDest <= storeInstructions_3_prfDest; // @[scheduler.scala 197:127]
    end
    if (reset) begin // @[scheduler.scala 76:34]
      storeInstructions_3_valid <= 1'h0; // @[scheduler.scala 76:34]
    end else if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_3_valid <= storeInstructionsUpdate_4_valid; // @[scheduler.scala 201:91]
    end else if (_storeInstructionsFree_T_2) begin // @[scheduler.scala 197:96]
      if (branchOps_valid) begin // @[scheduler.scala 177:27]
        storeInstructions_3_valid <= _GEN_30;
      end
    end else begin
      storeInstructions_3_valid <= storeInstructionsUpdate_4_valid; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_3_address <= fromBuffer_address; // @[scheduler.scala 201:91]
    end else if (!(_storeInstructionsFree_T_2)) begin // @[scheduler.scala 197:96]
      storeInstructions_3_address <= fromBuffer_address; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_3_instruction <= fromBuffer_instruction; // @[scheduler.scala 201:91]
    end else if (!(_storeInstructionsFree_T_2)) begin // @[scheduler.scala 197:96]
      storeInstructions_3_instruction <= fromBuffer_instruction; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_3_branchMask <= storeInstructionsUpdate_4_branchMask; // @[scheduler.scala 201:91]
    end else if (_storeInstructionsFree_T_2) begin // @[scheduler.scala 197:96]
      if (branchOps_valid) begin // @[scheduler.scala 177:27]
        if (|_T_30) begin // @[scheduler.scala 178:59]
          storeInstructions_3_branchMask <= _storeInstructionsUpdate_3_branchMask_T; // @[scheduler.scala 178:77]
        end
      end
    end else begin
      storeInstructions_3_branchMask <= storeInstructionsUpdate_4_branchMask; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_3_robAddr <= fromBuffer_robAddr; // @[scheduler.scala 201:91]
    end else if (!(_storeInstructionsFree_T_2)) begin // @[scheduler.scala 197:96]
      storeInstructions_3_robAddr <= fromBuffer_robAddr; // @[scheduler.scala 197:127]
    end
    if (storeCommit_fired) begin // @[scheduler.scala 198:27]
      storeInstructions_3_prfDest <= fromBuffer_prfDest; // @[scheduler.scala 201:91]
    end else if (!(_storeInstructionsFree_T_2)) begin // @[scheduler.scala 197:96]
      storeInstructions_3_prfDest <= fromBuffer_prfDest; // @[scheduler.scala 197:127]
    end
    if (reset) begin // @[scheduler.scala 86:27]
      fromBuffer_valid <= 1'h0; // @[scheduler.scala 86:27]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      if (branchOps_valid) begin // @[scheduler.scala 348:27]
        if (_T_80 & _T_380) begin // @[scheduler.scala 350:88]
          fromBuffer_valid <= 1'h0; // @[scheduler.scala 351:26]
        end else begin
          fromBuffer_valid <= _GEN_341;
        end
      end else begin
        fromBuffer_valid <= _GEN_341;
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 318:25]
      if (_T_83) begin // @[scheduler.scala 322:83]
        fromBuffer_valid <= 1'h0; // @[scheduler.scala 323:24]
      end
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      if (_T_377) begin // @[scheduler.scala 315:26]
        if (bufferQueue_0_valid) begin // @[Mux.scala 101:16]
          fromBuffer_address <= bufferQueue_0_address;
        end else if (bufferQueue_1_valid) begin // @[Mux.scala 101:16]
          fromBuffer_address <= bufferQueue_1_address;
        end else begin
          fromBuffer_address <= _nextFrmBuffer_T_19_address;
        end
      end else begin
        fromBuffer_address <= newInstruction_address;
      end
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      if (_T_377) begin // @[scheduler.scala 315:26]
        if (bufferQueue_0_valid) begin // @[Mux.scala 101:16]
          fromBuffer_instruction <= bufferQueue_0_instruction;
        end else if (bufferQueue_1_valid) begin // @[Mux.scala 101:16]
          fromBuffer_instruction <= bufferQueue_1_instruction;
        end else begin
          fromBuffer_instruction <= _nextFrmBuffer_T_19_instruction;
        end
      end else begin
        fromBuffer_instruction <= newInstruction_instruction;
      end
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      if (branchOps_valid) begin // @[scheduler.scala 348:27]
        if (|_T_379) begin // @[scheduler.scala 349:67]
          fromBuffer_branchMask <= _fromBuffer_branchMask_T_1; // @[scheduler.scala 349:90]
        end else begin
          fromBuffer_branchMask <= nextFrmBuffer_branchMask; // @[scheduler.scala 335:16]
        end
      end else begin
        fromBuffer_branchMask <= nextFrmBuffer_branchMask; // @[scheduler.scala 335:16]
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 177:27]
      if (_T_82) begin // @[scheduler.scala 178:59]
        fromBuffer_branchMask <= _storeInstructionsUpdate_4_branchMask_T; // @[scheduler.scala 178:77]
      end
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      if (_T_377) begin // @[scheduler.scala 315:26]
        if (bufferQueue_0_valid) begin // @[Mux.scala 101:16]
          fromBuffer_robAddr <= bufferQueue_0_robAddr;
        end else if (bufferQueue_1_valid) begin // @[Mux.scala 101:16]
          fromBuffer_robAddr <= bufferQueue_1_robAddr;
        end else begin
          fromBuffer_robAddr <= _nextFrmBuffer_T_19_robAddr;
        end
      end else begin
        fromBuffer_robAddr <= newInstruction_robAddr;
      end
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      if (_T_377) begin // @[scheduler.scala 315:26]
        if (bufferQueue_0_valid) begin // @[Mux.scala 101:16]
          fromBuffer_prfDest <= bufferQueue_0_prfDest;
        end else if (bufferQueue_1_valid) begin // @[Mux.scala 101:16]
          fromBuffer_prfDest <= bufferQueue_1_prfDest;
        end else begin
          fromBuffer_prfDest <= _nextFrmBuffer_T_19_prfDest;
        end
      end else begin
        fromBuffer_prfDest <= newInstruction_prfDest;
      end
    end
    toCache_replaying_REG <= replaying; // @[scheduler.scala 92:31]
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      if (branchOps_valid) begin // @[scheduler.scala 348:27]
        if (_T_80 & _T_380) begin // @[scheduler.scala 350:88]
          toPeripheral <= 1'h0; // @[scheduler.scala 352:22]
        end else begin
          toPeripheral <= nextFrmBuffer_valid & _T_326; // @[scheduler.scala 337:18]
        end
      end else begin
        toPeripheral <= nextFrmBuffer_valid & _T_326; // @[scheduler.scala 337:18]
      end
    end else if (branchOps_valid) begin // @[scheduler.scala 318:25]
      if (_T_83) begin // @[scheduler.scala 322:83]
        toPeripheral <= 1'h0; // @[scheduler.scala 324:20]
      end else begin
        toPeripheral <= _GEN_334;
      end
    end else begin
      toPeripheral <= _GEN_334;
    end
    REG <= storeCommit_fired; // @[scheduler.scala 245:17]
    REG_1 <= storeCommit_fired; // @[scheduler.scala 245:17]
    REG_2 <= storeCommit_fired; // @[scheduler.scala 245:17]
    REG_3 <= storeCommit_fired; // @[scheduler.scala 245:17]
    REG_4 <= storeCommit_fired; // @[scheduler.scala 245:17]
    if (reset) begin // @[scheduler.scala 294:28]
      bufferQueue_0_valid <= 1'h0; // @[scheduler.scala 294:28]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_0_valid <= bufferQueueUpdate_1_valid; // @[scheduler.scala 346:81]
    end else if (~bufferQueue_0_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_0_valid <= bufferQueueUpdate_1_valid; // @[scheduler.scala 302:103]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_0_valid <= _GEN_342;
    end else begin
      bufferQueue_0_valid <= _GEN_285;
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_0_address <= bufferQueue_1_address; // @[scheduler.scala 346:81]
    end else if (~bufferQueue_0_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_0_address <= bufferQueue_1_address; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_0_instruction <= bufferQueue_1_instruction; // @[scheduler.scala 346:81]
    end else if (~bufferQueue_0_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_0_instruction <= bufferQueue_1_instruction; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_0_branchMask <= bufferQueueUpdate_1_branchMask; // @[scheduler.scala 346:81]
    end else if (~bufferQueue_0_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_0_branchMask <= bufferQueueUpdate_1_branchMask; // @[scheduler.scala 302:103]
    end else if (branchOps_valid) begin // @[scheduler.scala 306:28]
      if (_T_238) begin // @[scheduler.scala 307:58]
        bufferQueue_0_branchMask <= _bufferQueueUpdate_0_branchMask_T; // @[scheduler.scala 307:77]
      end
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_0_robAddr <= bufferQueue_1_robAddr; // @[scheduler.scala 346:81]
    end else if (~bufferQueue_0_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_0_robAddr <= bufferQueue_1_robAddr; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_0_prfDest <= bufferQueue_1_prfDest; // @[scheduler.scala 346:81]
    end else if (~bufferQueue_0_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_0_prfDest <= bufferQueue_1_prfDest; // @[scheduler.scala 302:103]
    end
    if (reset) begin // @[scheduler.scala 294:28]
      bufferQueue_1_valid <= 1'h0; // @[scheduler.scala 294:28]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_1_valid <= bufferQueueUpdate_2_valid; // @[scheduler.scala 346:81]
    end else if (~bufferQueue_0_valid | ~bufferQueue_1_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_1_valid <= bufferQueueUpdate_2_valid; // @[scheduler.scala 302:103]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_1_valid <= _GEN_343;
    end else begin
      bufferQueue_1_valid <= _GEN_289;
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_1_address <= bufferQueue_2_address; // @[scheduler.scala 346:81]
    end else if (~bufferQueue_0_valid | ~bufferQueue_1_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_1_address <= bufferQueue_2_address; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_1_instruction <= bufferQueue_2_instruction; // @[scheduler.scala 346:81]
    end else if (~bufferQueue_0_valid | ~bufferQueue_1_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_1_instruction <= bufferQueue_2_instruction; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_1_branchMask <= bufferQueueUpdate_2_branchMask; // @[scheduler.scala 346:81]
    end else if (~bufferQueue_0_valid | ~bufferQueue_1_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_1_branchMask <= bufferQueueUpdate_2_branchMask; // @[scheduler.scala 302:103]
    end else if (branchOps_valid) begin // @[scheduler.scala 306:28]
      if (_T_244) begin // @[scheduler.scala 307:58]
        bufferQueue_1_branchMask <= _bufferQueueUpdate_1_branchMask_T; // @[scheduler.scala 307:77]
      end
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_1_robAddr <= bufferQueue_2_robAddr; // @[scheduler.scala 346:81]
    end else if (~bufferQueue_0_valid | ~bufferQueue_1_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_1_robAddr <= bufferQueue_2_robAddr; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_1_prfDest <= bufferQueue_2_prfDest; // @[scheduler.scala 346:81]
    end else if (~bufferQueue_0_valid | ~bufferQueue_1_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_1_prfDest <= bufferQueue_2_prfDest; // @[scheduler.scala 302:103]
    end
    if (reset) begin // @[scheduler.scala 294:28]
      bufferQueue_2_valid <= 1'h0; // @[scheduler.scala 294:28]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_2_valid <= bufferQueueUpdate_3_valid; // @[scheduler.scala 346:81]
    end else if (~_T_187 | ~bufferQueue_2_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_2_valid <= bufferQueueUpdate_3_valid; // @[scheduler.scala 302:103]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_2_valid <= _GEN_344;
    end else begin
      bufferQueue_2_valid <= _GEN_293;
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_2_address <= bufferQueue_3_address; // @[scheduler.scala 346:81]
    end else if (~_T_187 | ~bufferQueue_2_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_2_address <= bufferQueue_3_address; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_2_instruction <= bufferQueue_3_instruction; // @[scheduler.scala 346:81]
    end else if (~_T_187 | ~bufferQueue_2_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_2_instruction <= bufferQueue_3_instruction; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_2_branchMask <= bufferQueueUpdate_3_branchMask; // @[scheduler.scala 346:81]
    end else if (~_T_187 | ~bufferQueue_2_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_2_branchMask <= bufferQueueUpdate_3_branchMask; // @[scheduler.scala 302:103]
    end else if (branchOps_valid) begin // @[scheduler.scala 306:28]
      if (_T_250) begin // @[scheduler.scala 307:58]
        bufferQueue_2_branchMask <= _bufferQueueUpdate_2_branchMask_T; // @[scheduler.scala 307:77]
      end
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_2_robAddr <= bufferQueue_3_robAddr; // @[scheduler.scala 346:81]
    end else if (~_T_187 | ~bufferQueue_2_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_2_robAddr <= bufferQueue_3_robAddr; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_2_prfDest <= bufferQueue_3_prfDest; // @[scheduler.scala 346:81]
    end else if (~_T_187 | ~bufferQueue_2_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_2_prfDest <= bufferQueue_3_prfDest; // @[scheduler.scala 302:103]
    end
    if (reset) begin // @[scheduler.scala 294:28]
      bufferQueue_3_valid <= 1'h0; // @[scheduler.scala 294:28]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_3_valid <= bufferQueueUpdate_4_valid; // @[scheduler.scala 346:81]
    end else if (~_T_188 | ~bufferQueue_3_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_3_valid <= bufferQueueUpdate_4_valid; // @[scheduler.scala 302:103]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_3_valid <= _GEN_345;
    end else begin
      bufferQueue_3_valid <= _GEN_297;
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_3_address <= bufferQueue_4_address; // @[scheduler.scala 346:81]
    end else if (~_T_188 | ~bufferQueue_3_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_3_address <= bufferQueue_4_address; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_3_instruction <= bufferQueue_4_instruction; // @[scheduler.scala 346:81]
    end else if (~_T_188 | ~bufferQueue_3_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_3_instruction <= bufferQueue_4_instruction; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_3_branchMask <= bufferQueueUpdate_4_branchMask; // @[scheduler.scala 346:81]
    end else if (~_T_188 | ~bufferQueue_3_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_3_branchMask <= bufferQueueUpdate_4_branchMask; // @[scheduler.scala 302:103]
    end else if (branchOps_valid) begin // @[scheduler.scala 306:28]
      if (_T_256) begin // @[scheduler.scala 307:58]
        bufferQueue_3_branchMask <= _bufferQueueUpdate_3_branchMask_T; // @[scheduler.scala 307:77]
      end
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_3_robAddr <= bufferQueue_4_robAddr; // @[scheduler.scala 346:81]
    end else if (~_T_188 | ~bufferQueue_3_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_3_robAddr <= bufferQueue_4_robAddr; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_3_prfDest <= bufferQueue_4_prfDest; // @[scheduler.scala 346:81]
    end else if (~_T_188 | ~bufferQueue_3_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_3_prfDest <= bufferQueue_4_prfDest; // @[scheduler.scala 302:103]
    end
    if (reset) begin // @[scheduler.scala 294:28]
      bufferQueue_4_valid <= 1'h0; // @[scheduler.scala 294:28]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_4_valid <= bufferQueueUpdate_5_valid; // @[scheduler.scala 346:81]
    end else if (~_T_189 | ~bufferQueue_4_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_4_valid <= bufferQueueUpdate_5_valid; // @[scheduler.scala 302:103]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_4_valid <= _GEN_346;
    end else begin
      bufferQueue_4_valid <= _GEN_301;
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_4_address <= bufferQueue_5_address; // @[scheduler.scala 346:81]
    end else if (~_T_189 | ~bufferQueue_4_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_4_address <= bufferQueue_5_address; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_4_instruction <= bufferQueue_5_instruction; // @[scheduler.scala 346:81]
    end else if (~_T_189 | ~bufferQueue_4_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_4_instruction <= bufferQueue_5_instruction; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_4_branchMask <= bufferQueueUpdate_5_branchMask; // @[scheduler.scala 346:81]
    end else if (~_T_189 | ~bufferQueue_4_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_4_branchMask <= bufferQueueUpdate_5_branchMask; // @[scheduler.scala 302:103]
    end else if (branchOps_valid) begin // @[scheduler.scala 306:28]
      if (_T_262) begin // @[scheduler.scala 307:58]
        bufferQueue_4_branchMask <= _bufferQueueUpdate_4_branchMask_T; // @[scheduler.scala 307:77]
      end
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_4_robAddr <= bufferQueue_5_robAddr; // @[scheduler.scala 346:81]
    end else if (~_T_189 | ~bufferQueue_4_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_4_robAddr <= bufferQueue_5_robAddr; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_4_prfDest <= bufferQueue_5_prfDest; // @[scheduler.scala 346:81]
    end else if (~_T_189 | ~bufferQueue_4_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_4_prfDest <= bufferQueue_5_prfDest; // @[scheduler.scala 302:103]
    end
    if (reset) begin // @[scheduler.scala 294:28]
      bufferQueue_5_valid <= 1'h0; // @[scheduler.scala 294:28]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_5_valid <= bufferQueueUpdate_6_valid; // @[scheduler.scala 346:81]
    end else if (~_T_190 | ~bufferQueue_5_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_5_valid <= bufferQueueUpdate_6_valid; // @[scheduler.scala 302:103]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_5_valid <= _GEN_347;
    end else begin
      bufferQueue_5_valid <= _GEN_305;
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_5_address <= bufferQueue_6_address; // @[scheduler.scala 346:81]
    end else if (~_T_190 | ~bufferQueue_5_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_5_address <= bufferQueue_6_address; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_5_instruction <= bufferQueue_6_instruction; // @[scheduler.scala 346:81]
    end else if (~_T_190 | ~bufferQueue_5_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_5_instruction <= bufferQueue_6_instruction; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_5_branchMask <= bufferQueueUpdate_6_branchMask; // @[scheduler.scala 346:81]
    end else if (~_T_190 | ~bufferQueue_5_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_5_branchMask <= bufferQueueUpdate_6_branchMask; // @[scheduler.scala 302:103]
    end else if (branchOps_valid) begin // @[scheduler.scala 306:28]
      if (_T_268) begin // @[scheduler.scala 307:58]
        bufferQueue_5_branchMask <= _bufferQueueUpdate_5_branchMask_T; // @[scheduler.scala 307:77]
      end
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_5_robAddr <= bufferQueue_6_robAddr; // @[scheduler.scala 346:81]
    end else if (~_T_190 | ~bufferQueue_5_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_5_robAddr <= bufferQueue_6_robAddr; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_5_prfDest <= bufferQueue_6_prfDest; // @[scheduler.scala 346:81]
    end else if (~_T_190 | ~bufferQueue_5_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_5_prfDest <= bufferQueue_6_prfDest; // @[scheduler.scala 302:103]
    end
    if (reset) begin // @[scheduler.scala 294:28]
      bufferQueue_6_valid <= 1'h0; // @[scheduler.scala 294:28]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_6_valid <= bufferQueueUpdate_7_valid; // @[scheduler.scala 346:81]
    end else if (~_T_191 | ~bufferQueue_6_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_6_valid <= bufferQueueUpdate_7_valid; // @[scheduler.scala 302:103]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_6_valid <= _GEN_348;
    end else begin
      bufferQueue_6_valid <= _GEN_309;
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_6_address <= bufferQueue_7_address; // @[scheduler.scala 346:81]
    end else if (~_T_191 | ~bufferQueue_6_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_6_address <= bufferQueue_7_address; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_6_instruction <= bufferQueue_7_instruction; // @[scheduler.scala 346:81]
    end else if (~_T_191 | ~bufferQueue_6_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_6_instruction <= bufferQueue_7_instruction; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_6_branchMask <= bufferQueueUpdate_7_branchMask; // @[scheduler.scala 346:81]
    end else if (~_T_191 | ~bufferQueue_6_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_6_branchMask <= bufferQueueUpdate_7_branchMask; // @[scheduler.scala 302:103]
    end else if (branchOps_valid) begin // @[scheduler.scala 306:28]
      if (_T_274) begin // @[scheduler.scala 307:58]
        bufferQueue_6_branchMask <= _bufferQueueUpdate_6_branchMask_T; // @[scheduler.scala 307:77]
      end
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_6_robAddr <= bufferQueue_7_robAddr; // @[scheduler.scala 346:81]
    end else if (~_T_191 | ~bufferQueue_6_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_6_robAddr <= bufferQueue_7_robAddr; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_6_prfDest <= bufferQueue_7_prfDest; // @[scheduler.scala 346:81]
    end else if (~_T_191 | ~bufferQueue_6_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_6_prfDest <= bufferQueue_7_prfDest; // @[scheduler.scala 302:103]
    end
    if (reset) begin // @[scheduler.scala 294:28]
      bufferQueue_7_valid <= 1'h0; // @[scheduler.scala 294:28]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_7_valid <= bufferQueueUpdate_8_valid; // @[scheduler.scala 346:81]
    end else if (~_T_192 | ~bufferQueue_7_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_7_valid <= bufferQueueUpdate_8_valid; // @[scheduler.scala 302:103]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_7_valid <= _GEN_349;
    end else begin
      bufferQueue_7_valid <= _GEN_313;
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_7_address <= bufferQueue_8_address; // @[scheduler.scala 346:81]
    end else if (~_T_192 | ~bufferQueue_7_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_7_address <= bufferQueue_8_address; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_7_instruction <= bufferQueue_8_instruction; // @[scheduler.scala 346:81]
    end else if (~_T_192 | ~bufferQueue_7_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_7_instruction <= bufferQueue_8_instruction; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_7_branchMask <= bufferQueueUpdate_8_branchMask; // @[scheduler.scala 346:81]
    end else if (~_T_192 | ~bufferQueue_7_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_7_branchMask <= bufferQueueUpdate_8_branchMask; // @[scheduler.scala 302:103]
    end else if (branchOps_valid) begin // @[scheduler.scala 306:28]
      if (_T_280) begin // @[scheduler.scala 307:58]
        bufferQueue_7_branchMask <= _bufferQueueUpdate_7_branchMask_T; // @[scheduler.scala 307:77]
      end
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_7_robAddr <= bufferQueue_8_robAddr; // @[scheduler.scala 346:81]
    end else if (~_T_192 | ~bufferQueue_7_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_7_robAddr <= bufferQueue_8_robAddr; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_7_prfDest <= bufferQueue_8_prfDest; // @[scheduler.scala 346:81]
    end else if (~_T_192 | ~bufferQueue_7_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_7_prfDest <= bufferQueue_8_prfDest; // @[scheduler.scala 302:103]
    end
    if (reset) begin // @[scheduler.scala 294:28]
      bufferQueue_8_valid <= 1'h0; // @[scheduler.scala 294:28]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_8_valid <= bufferQueueUpdate_9_valid; // @[scheduler.scala 346:81]
    end else if (~_T_193 | ~bufferQueue_8_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_8_valid <= bufferQueueUpdate_9_valid; // @[scheduler.scala 302:103]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_8_valid <= _GEN_350;
    end else begin
      bufferQueue_8_valid <= _GEN_317;
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_8_address <= bufferQueue_9_address; // @[scheduler.scala 346:81]
    end else if (~_T_193 | ~bufferQueue_8_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_8_address <= bufferQueue_9_address; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_8_instruction <= bufferQueue_9_instruction; // @[scheduler.scala 346:81]
    end else if (~_T_193 | ~bufferQueue_8_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_8_instruction <= bufferQueue_9_instruction; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_8_branchMask <= bufferQueueUpdate_9_branchMask; // @[scheduler.scala 346:81]
    end else if (~_T_193 | ~bufferQueue_8_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_8_branchMask <= bufferQueueUpdate_9_branchMask; // @[scheduler.scala 302:103]
    end else if (branchOps_valid) begin // @[scheduler.scala 306:28]
      if (_T_286) begin // @[scheduler.scala 307:58]
        bufferQueue_8_branchMask <= _bufferQueueUpdate_8_branchMask_T; // @[scheduler.scala 307:77]
      end
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_8_robAddr <= bufferQueue_9_robAddr; // @[scheduler.scala 346:81]
    end else if (~_T_193 | ~bufferQueue_8_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_8_robAddr <= bufferQueue_9_robAddr; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_8_prfDest <= bufferQueue_9_prfDest; // @[scheduler.scala 346:81]
    end else if (~_T_193 | ~bufferQueue_8_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_8_prfDest <= bufferQueue_9_prfDest; // @[scheduler.scala 302:103]
    end
    if (reset) begin // @[scheduler.scala 294:28]
      bufferQueue_9_valid <= 1'h0; // @[scheduler.scala 294:28]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_9_valid <= bufferQueueUpdate_10_valid; // @[scheduler.scala 346:81]
    end else if (~_T_194 | ~bufferQueue_9_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_9_valid <= bufferQueueUpdate_10_valid; // @[scheduler.scala 302:103]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_9_valid <= _GEN_351;
    end else begin
      bufferQueue_9_valid <= _GEN_321;
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_9_address <= bufferQueue_10_address; // @[scheduler.scala 346:81]
    end else if (~_T_194 | ~bufferQueue_9_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_9_address <= bufferQueue_10_address; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_9_instruction <= bufferQueue_10_instruction; // @[scheduler.scala 346:81]
    end else if (~_T_194 | ~bufferQueue_9_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_9_instruction <= bufferQueue_10_instruction; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_9_branchMask <= bufferQueueUpdate_10_branchMask; // @[scheduler.scala 346:81]
    end else if (~_T_194 | ~bufferQueue_9_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_9_branchMask <= bufferQueueUpdate_10_branchMask; // @[scheduler.scala 302:103]
    end else if (branchOps_valid) begin // @[scheduler.scala 306:28]
      if (_T_292) begin // @[scheduler.scala 307:58]
        bufferQueue_9_branchMask <= _bufferQueueUpdate_9_branchMask_T; // @[scheduler.scala 307:77]
      end
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_9_robAddr <= bufferQueue_10_robAddr; // @[scheduler.scala 346:81]
    end else if (~_T_194 | ~bufferQueue_9_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_9_robAddr <= bufferQueue_10_robAddr; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_9_prfDest <= bufferQueue_10_prfDest; // @[scheduler.scala 346:81]
    end else if (~_T_194 | ~bufferQueue_9_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_9_prfDest <= bufferQueue_10_prfDest; // @[scheduler.scala 302:103]
    end
    if (reset) begin // @[scheduler.scala 294:28]
      bufferQueue_10_valid <= 1'h0; // @[scheduler.scala 294:28]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_10_valid <= bufferQueueUpdate_11_valid; // @[scheduler.scala 346:81]
    end else if (~_T_195 | ~bufferQueue_10_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_10_valid <= bufferQueueUpdate_11_valid; // @[scheduler.scala 302:103]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_10_valid <= _GEN_352;
    end else begin
      bufferQueue_10_valid <= _GEN_325;
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_10_address <= bufferQueue_11_address; // @[scheduler.scala 346:81]
    end else if (~_T_195 | ~bufferQueue_10_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_10_address <= bufferQueue_11_address; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_10_instruction <= bufferQueue_11_instruction; // @[scheduler.scala 346:81]
    end else if (~_T_195 | ~bufferQueue_10_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_10_instruction <= bufferQueue_11_instruction; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_10_branchMask <= bufferQueueUpdate_11_branchMask; // @[scheduler.scala 346:81]
    end else if (~_T_195 | ~bufferQueue_10_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_10_branchMask <= bufferQueueUpdate_11_branchMask; // @[scheduler.scala 302:103]
    end else if (branchOps_valid) begin // @[scheduler.scala 306:28]
      if (_T_298) begin // @[scheduler.scala 307:58]
        bufferQueue_10_branchMask <= _bufferQueueUpdate_10_branchMask_T; // @[scheduler.scala 307:77]
      end
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_10_robAddr <= bufferQueue_11_robAddr; // @[scheduler.scala 346:81]
    end else if (~_T_195 | ~bufferQueue_10_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_10_robAddr <= bufferQueue_11_robAddr; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_10_prfDest <= bufferQueue_11_prfDest; // @[scheduler.scala 346:81]
    end else if (~_T_195 | ~bufferQueue_10_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_10_prfDest <= bufferQueue_11_prfDest; // @[scheduler.scala 302:103]
    end
    if (reset) begin // @[scheduler.scala 294:28]
      bufferQueue_11_valid <= 1'h0; // @[scheduler.scala 294:28]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_11_valid <= bufferQueueUpdate_12_valid; // @[scheduler.scala 346:81]
    end else if (~_T_196 | ~bufferQueue_11_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_11_valid <= bufferQueueUpdate_12_valid; // @[scheduler.scala 302:103]
    end else if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_11_valid <= _GEN_353;
    end else begin
      bufferQueue_11_valid <= _GEN_329;
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_11_address <= newInstruction_address; // @[scheduler.scala 346:81]
    end else if (~_T_196 | ~bufferQueue_11_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_11_address <= newInstruction_address; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_11_instruction <= newInstruction_instruction; // @[scheduler.scala 346:81]
    end else if (~_T_196 | ~bufferQueue_11_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_11_instruction <= newInstruction_instruction; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_11_branchMask <= bufferQueueUpdate_12_branchMask; // @[scheduler.scala 346:81]
    end else if (~_T_196 | ~bufferQueue_11_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_11_branchMask <= bufferQueueUpdate_12_branchMask; // @[scheduler.scala 302:103]
    end else if (branchOps_valid) begin // @[scheduler.scala 306:28]
      if (_T_304) begin // @[scheduler.scala 307:58]
        bufferQueue_11_branchMask <= _bufferQueueUpdate_11_branchMask_T; // @[scheduler.scala 307:77]
      end
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_11_robAddr <= newInstruction_robAddr; // @[scheduler.scala 346:81]
    end else if (~_T_196 | ~bufferQueue_11_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_11_robAddr <= newInstruction_robAddr; // @[scheduler.scala 302:103]
    end
    if ((dequeuedFromBuffer | ~fromBuffer_valid) & _dequeuedFromBuffer_T_1) begin // @[scheduler.scala 334:90]
      bufferQueue_11_prfDest <= newInstruction_prfDest; // @[scheduler.scala 346:81]
    end else if (~_T_196 | ~bufferQueue_11_valid) begin // @[scheduler.scala 302:98]
      bufferQueue_11_prfDest <= newInstruction_prfDest; // @[scheduler.scala 302:103]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  scheduledInstruction_query_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  scheduledInstruction_query_address = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  scheduledInstruction_query_instruction = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  scheduledInstruction_query_branchMask = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  scheduledInstruction_query_robAddr = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  scheduledInstruction_query_prfDest = _RAND_5[5:0];
  _RAND_6 = {2{`RANDOM}};
  scheduledInstruction_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  dependentReads_0_valid = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  dependentReads_0_address = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  dependentReads_0_instruction = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  dependentReads_0_branchMask = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  dependentReads_0_robAddr = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  dependentReads_0_prfDest = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  dependentReads_0_dependency_free = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  dependentReads_0_dependency_robAddr = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  dependentReads_1_valid = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  dependentReads_1_address = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  dependentReads_1_instruction = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  dependentReads_1_branchMask = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  dependentReads_1_robAddr = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  dependentReads_1_prfDest = _RAND_20[5:0];
  _RAND_21 = {1{`RANDOM}};
  dependentReads_1_dependency_free = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  dependentReads_1_dependency_robAddr = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  dependentReads_2_valid = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  dependentReads_2_address = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  dependentReads_2_instruction = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  dependentReads_2_branchMask = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  dependentReads_2_robAddr = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  dependentReads_2_prfDest = _RAND_28[5:0];
  _RAND_29 = {1{`RANDOM}};
  dependentReads_2_dependency_free = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  dependentReads_2_dependency_robAddr = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  dependentReads_3_valid = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  dependentReads_3_address = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  dependentReads_3_instruction = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  dependentReads_3_branchMask = _RAND_34[3:0];
  _RAND_35 = {1{`RANDOM}};
  dependentReads_3_robAddr = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  dependentReads_3_prfDest = _RAND_36[5:0];
  _RAND_37 = {1{`RANDOM}};
  dependentReads_3_dependency_free = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  dependentReads_3_dependency_robAddr = _RAND_38[3:0];
  _RAND_39 = {1{`RANDOM}};
  storeInstructions_0_valid = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  storeInstructions_0_address = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  storeInstructions_0_instruction = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  storeInstructions_0_branchMask = _RAND_42[3:0];
  _RAND_43 = {1{`RANDOM}};
  storeInstructions_0_robAddr = _RAND_43[3:0];
  _RAND_44 = {1{`RANDOM}};
  storeInstructions_0_prfDest = _RAND_44[5:0];
  _RAND_45 = {1{`RANDOM}};
  storeInstructions_1_valid = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  storeInstructions_1_address = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  storeInstructions_1_instruction = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  storeInstructions_1_branchMask = _RAND_48[3:0];
  _RAND_49 = {1{`RANDOM}};
  storeInstructions_1_robAddr = _RAND_49[3:0];
  _RAND_50 = {1{`RANDOM}};
  storeInstructions_1_prfDest = _RAND_50[5:0];
  _RAND_51 = {1{`RANDOM}};
  storeInstructions_2_valid = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  storeInstructions_2_address = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  storeInstructions_2_instruction = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  storeInstructions_2_branchMask = _RAND_54[3:0];
  _RAND_55 = {1{`RANDOM}};
  storeInstructions_2_robAddr = _RAND_55[3:0];
  _RAND_56 = {1{`RANDOM}};
  storeInstructions_2_prfDest = _RAND_56[5:0];
  _RAND_57 = {1{`RANDOM}};
  storeInstructions_3_valid = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  storeInstructions_3_address = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  storeInstructions_3_instruction = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  storeInstructions_3_branchMask = _RAND_60[3:0];
  _RAND_61 = {1{`RANDOM}};
  storeInstructions_3_robAddr = _RAND_61[3:0];
  _RAND_62 = {1{`RANDOM}};
  storeInstructions_3_prfDest = _RAND_62[5:0];
  _RAND_63 = {1{`RANDOM}};
  fromBuffer_valid = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  fromBuffer_address = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  fromBuffer_instruction = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  fromBuffer_branchMask = _RAND_66[3:0];
  _RAND_67 = {1{`RANDOM}};
  fromBuffer_robAddr = _RAND_67[3:0];
  _RAND_68 = {1{`RANDOM}};
  fromBuffer_prfDest = _RAND_68[5:0];
  _RAND_69 = {1{`RANDOM}};
  toCache_replaying_REG = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  toPeripheral = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  REG = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  REG_1 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  REG_2 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  REG_3 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  REG_4 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  bufferQueue_0_valid = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  bufferQueue_0_address = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  bufferQueue_0_instruction = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  bufferQueue_0_branchMask = _RAND_79[3:0];
  _RAND_80 = {1{`RANDOM}};
  bufferQueue_0_robAddr = _RAND_80[3:0];
  _RAND_81 = {1{`RANDOM}};
  bufferQueue_0_prfDest = _RAND_81[5:0];
  _RAND_82 = {1{`RANDOM}};
  bufferQueue_1_valid = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  bufferQueue_1_address = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  bufferQueue_1_instruction = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  bufferQueue_1_branchMask = _RAND_85[3:0];
  _RAND_86 = {1{`RANDOM}};
  bufferQueue_1_robAddr = _RAND_86[3:0];
  _RAND_87 = {1{`RANDOM}};
  bufferQueue_1_prfDest = _RAND_87[5:0];
  _RAND_88 = {1{`RANDOM}};
  bufferQueue_2_valid = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  bufferQueue_2_address = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  bufferQueue_2_instruction = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  bufferQueue_2_branchMask = _RAND_91[3:0];
  _RAND_92 = {1{`RANDOM}};
  bufferQueue_2_robAddr = _RAND_92[3:0];
  _RAND_93 = {1{`RANDOM}};
  bufferQueue_2_prfDest = _RAND_93[5:0];
  _RAND_94 = {1{`RANDOM}};
  bufferQueue_3_valid = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  bufferQueue_3_address = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  bufferQueue_3_instruction = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  bufferQueue_3_branchMask = _RAND_97[3:0];
  _RAND_98 = {1{`RANDOM}};
  bufferQueue_3_robAddr = _RAND_98[3:0];
  _RAND_99 = {1{`RANDOM}};
  bufferQueue_3_prfDest = _RAND_99[5:0];
  _RAND_100 = {1{`RANDOM}};
  bufferQueue_4_valid = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  bufferQueue_4_address = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  bufferQueue_4_instruction = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  bufferQueue_4_branchMask = _RAND_103[3:0];
  _RAND_104 = {1{`RANDOM}};
  bufferQueue_4_robAddr = _RAND_104[3:0];
  _RAND_105 = {1{`RANDOM}};
  bufferQueue_4_prfDest = _RAND_105[5:0];
  _RAND_106 = {1{`RANDOM}};
  bufferQueue_5_valid = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  bufferQueue_5_address = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  bufferQueue_5_instruction = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  bufferQueue_5_branchMask = _RAND_109[3:0];
  _RAND_110 = {1{`RANDOM}};
  bufferQueue_5_robAddr = _RAND_110[3:0];
  _RAND_111 = {1{`RANDOM}};
  bufferQueue_5_prfDest = _RAND_111[5:0];
  _RAND_112 = {1{`RANDOM}};
  bufferQueue_6_valid = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  bufferQueue_6_address = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  bufferQueue_6_instruction = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  bufferQueue_6_branchMask = _RAND_115[3:0];
  _RAND_116 = {1{`RANDOM}};
  bufferQueue_6_robAddr = _RAND_116[3:0];
  _RAND_117 = {1{`RANDOM}};
  bufferQueue_6_prfDest = _RAND_117[5:0];
  _RAND_118 = {1{`RANDOM}};
  bufferQueue_7_valid = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  bufferQueue_7_address = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  bufferQueue_7_instruction = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  bufferQueue_7_branchMask = _RAND_121[3:0];
  _RAND_122 = {1{`RANDOM}};
  bufferQueue_7_robAddr = _RAND_122[3:0];
  _RAND_123 = {1{`RANDOM}};
  bufferQueue_7_prfDest = _RAND_123[5:0];
  _RAND_124 = {1{`RANDOM}};
  bufferQueue_8_valid = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  bufferQueue_8_address = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  bufferQueue_8_instruction = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  bufferQueue_8_branchMask = _RAND_127[3:0];
  _RAND_128 = {1{`RANDOM}};
  bufferQueue_8_robAddr = _RAND_128[3:0];
  _RAND_129 = {1{`RANDOM}};
  bufferQueue_8_prfDest = _RAND_129[5:0];
  _RAND_130 = {1{`RANDOM}};
  bufferQueue_9_valid = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  bufferQueue_9_address = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  bufferQueue_9_instruction = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  bufferQueue_9_branchMask = _RAND_133[3:0];
  _RAND_134 = {1{`RANDOM}};
  bufferQueue_9_robAddr = _RAND_134[3:0];
  _RAND_135 = {1{`RANDOM}};
  bufferQueue_9_prfDest = _RAND_135[5:0];
  _RAND_136 = {1{`RANDOM}};
  bufferQueue_10_valid = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  bufferQueue_10_address = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  bufferQueue_10_instruction = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  bufferQueue_10_branchMask = _RAND_139[3:0];
  _RAND_140 = {1{`RANDOM}};
  bufferQueue_10_robAddr = _RAND_140[3:0];
  _RAND_141 = {1{`RANDOM}};
  bufferQueue_10_prfDest = _RAND_141[5:0];
  _RAND_142 = {1{`RANDOM}};
  bufferQueue_11_valid = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  bufferQueue_11_address = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  bufferQueue_11_instruction = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  bufferQueue_11_branchMask = _RAND_145[3:0];
  _RAND_146 = {1{`RANDOM}};
  bufferQueue_11_robAddr = _RAND_146[3:0];
  _RAND_147 = {1{`RANDOM}};
  bufferQueue_11_prfDest = _RAND_147[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module peripheralHandler(
  input         clock,
  input         reset,
  input         request_valid,
  input  [31:0] request_address,
  input  [31:0] request_instruction,
  input  [3:0]  request_branchMask,
  input  [3:0]  request_robAddr,
  input  [5:0]  request_prfDest,
  output        finishedRequest_valid,
  output [31:0] finishedRequest_address,
  output [31:0] finishedRequest_instruction,
  output [3:0]  finishedRequest_robAddr,
  output [5:0]  finishedRequest_prfDest,
  output        ready,
  input         branchOps_valid,
  input  [3:0]  branchOps_branchMask,
  input         branchOps_passed,
  output [31:0] axi_AWADDR,
  output [7:0]  axi_AWLEN,
  output [2:0]  axi_AWSIZE,
  output        axi_AWVALID,
  input         axi_AWREADY,
  output [31:0] axi_WDATA,
  output [3:0]  axi_WSTRB,
  output        axi_WLAST,
  output        axi_WVALID,
  input         axi_WREADY,
  input         axi_BVALID,
  output        axi_BREADY,
  output [31:0] axi_ARADDR,
  output [7:0]  axi_ARLEN,
  output [2:0]  axi_ARSIZE,
  output        axi_ARVALID,
  input         axi_ARREADY,
  input  [31:0] axi_RDATA,
  input         axi_RLAST,
  input         axi_RVALID,
  output        axi_RREADY,
  output        readFinished_ready,
  input         readFinished_fired,
  output [63:0] readDataOut,
  input         writeIn_valid,
  input  [63:0] writeIn_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  reg  servicing_valid; // @[peripheralHandler.scala 12:26]
  reg [31:0] servicing_address; // @[peripheralHandler.scala 12:26]
  reg [31:0] servicing_instruction; // @[peripheralHandler.scala 12:26]
  reg [3:0] servicing_branchMask; // @[peripheralHandler.scala 12:26]
  reg [3:0] servicing_robAddr; // @[peripheralHandler.scala 12:26]
  reg [5:0] servicing_prfDest; // @[peripheralHandler.scala 12:26]
  reg  arvalid; // @[peripheralHandler.scala 17:71]
  reg  rready; // @[peripheralHandler.scala 17:71]
  reg  awvalid; // @[peripheralHandler.scala 17:71]
  reg  wvalid; // @[peripheralHandler.scala 17:71]
  reg  wlast; // @[peripheralHandler.scala 17:71]
  reg  bready; // @[peripheralHandler.scala 17:71]
  reg  stall; // @[peripheralHandler.scala 17:71]
  reg [63:0] rdata; // @[peripheralHandler.scala 22:18]
  reg  writeCleared; // @[peripheralHandler.scala 30:29]
  wire  _GEN_0 = request_instruction[5] | awvalid; // @[peripheralHandler.scala 34:{41,51} 17:71]
  wire  _GEN_1 = request_instruction[5] ? arvalid : 1'h1; // @[peripheralHandler.scala 34:41 17:71 35:26]
  wire [3:0] _T_3 = branchOps_branchMask & request_branchMask; // @[peripheralHandler.scala 37:34]
  wire  _T_4 = |_T_3; // @[peripheralHandler.scala 37:56]
  wire [3:0] _servicing_branchMask_T = branchOps_branchMask ^ request_branchMask; // @[peripheralHandler.scala 38:54]
  wire [3:0] _GEN_2 = |_T_3 ? _servicing_branchMask_T : request_branchMask; // @[peripheralHandler.scala 33:15 37:61 38:30]
  wire  _T_5 = ~branchOps_passed; // @[peripheralHandler.scala 40:12]
  wire  _GEN_3 = ~branchOps_passed & _T_4 ? 1'h0 : _GEN_0; // @[peripheralHandler.scala 40:82 41:17]
  wire  _GEN_4 = ~branchOps_passed & _T_4 ? 1'h0 : _GEN_1; // @[peripheralHandler.scala 40:82 42:17]
  wire  _GEN_5 = ~branchOps_passed & _T_4 ? 1'h0 : request_valid; // @[peripheralHandler.scala 33:15 40:82 43:25]
  wire [3:0] _GEN_6 = branchOps_valid ? _GEN_2 : request_branchMask; // @[peripheralHandler.scala 33:15 36:27]
  wire  _GEN_7 = branchOps_valid ? _GEN_3 : _GEN_0; // @[peripheralHandler.scala 36:27]
  wire  _GEN_8 = branchOps_valid ? _GEN_4 : _GEN_1; // @[peripheralHandler.scala 36:27]
  wire  _GEN_9 = branchOps_valid ? _GEN_5 : request_valid; // @[peripheralHandler.scala 33:15 36:27]
  wire  _GEN_10 = request_valid & ready ? _GEN_9 : servicing_valid; // @[peripheralHandler.scala 12:26 32:32]
  wire [3:0] _GEN_13 = request_valid & ready ? _GEN_6 : servicing_branchMask; // @[peripheralHandler.scala 12:26 32:32]
  wire  _GEN_16 = request_valid & ready ? _GEN_7 : awvalid; // @[peripheralHandler.scala 32:32 17:71]
  wire  _GEN_17 = request_valid & ready ? _GEN_8 : arvalid; // @[peripheralHandler.scala 32:32 17:71]
  wire  _GEN_18 = axi_ARVALID & axi_ARREADY ? 1'h0 : _GEN_17; // @[peripheralHandler.scala 50:36 51:13]
  wire  _GEN_19 = axi_ARVALID & axi_ARREADY | rready; // @[peripheralHandler.scala 50:36 52:12 17:71]
  wire  _T_10 = axi_RVALID & axi_RREADY; // @[peripheralHandler.scala 55:19]
  wire  _T_11 = axi_RVALID & axi_RREADY & axi_RLAST; // @[peripheralHandler.scala 55:33]
  wire  _GEN_20 = servicing_valid | stall; // @[peripheralHandler.scala 57:27 58:13 17:71]
  wire  _GEN_22 = axi_RVALID & axi_RREADY & axi_RLAST ? _GEN_20 : stall; // @[peripheralHandler.scala 55:47 17:71]
  wire  _GEN_23 = readFinished_fired ? 1'h0 : _GEN_22; // @[peripheralHandler.scala 65:28 66:11]
  wire  _GEN_24 = readFinished_fired ? 1'h0 : _GEN_10; // @[peripheralHandler.scala 65:28 67:21]
  wire  _T_15 = servicing_instruction[13:12] == 2'h3; // @[peripheralHandler.scala 74:40]
  wire [63:0] _rdata_T_1 = {axi_RDATA,rdata[31:0]}; // @[Cat.scala 33:92]
  wire  _GEN_26 = 2'h1 == servicing_address[1:0] ? axi_RDATA[15] : axi_RDATA[7]; // @[peripheralHandler.scala 78:{26,26}]
  wire  _GEN_27 = 2'h2 == servicing_address[1:0] ? axi_RDATA[23] : _GEN_26; // @[peripheralHandler.scala 78:{26,26}]
  wire  _GEN_28 = 2'h3 == servicing_address[1:0] ? axi_RDATA[31] : _GEN_27; // @[peripheralHandler.scala 78:{26,26}]
  wire  _GEN_30 = servicing_address[2] ? axi_RDATA[31] : axi_RDATA[15]; // @[peripheralHandler.scala 78:{26,26}]
  wire  _rdata_T_4 = ~servicing_instruction[14]; // @[peripheralHandler.scala 84:28]
  wire  _GEN_32 = servicing_instruction[12] ? _GEN_30 : _GEN_28; // @[peripheralHandler.scala 84:{27,27}]
  wire  _rdata_T_5 = ~servicing_instruction[14] & _GEN_32; // @[peripheralHandler.scala 84:27]
  wire [55:0] _rdata_T_7 = _rdata_T_5 ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _GEN_34 = 2'h1 == servicing_address[1:0] ? axi_RDATA[15:8] : axi_RDATA[7:0]; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_35 = 2'h2 == servicing_address[1:0] ? axi_RDATA[23:16] : _GEN_34; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_36 = 2'h3 == servicing_address[1:0] ? axi_RDATA[31:24] : _GEN_35; // @[Cat.scala 33:{92,92}]
  wire [63:0] _rdata_T_13 = {_rdata_T_7,_GEN_36}; // @[Cat.scala 33:92]
  wire [47:0] _rdata_T_19 = _rdata_T_5 ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 77:12]
  wire [15:0] _GEN_38 = servicing_address[2] ? axi_RDATA[31:16] : axi_RDATA[15:0]; // @[Cat.scala 33:{92,92}]
  wire [63:0] _rdata_T_23 = {_rdata_T_19,_GEN_38}; // @[Cat.scala 33:92]
  wire  _rdata_T_28 = _rdata_T_4 & axi_RDATA[31]; // @[peripheralHandler.scala 86:27]
  wire [31:0] _rdata_T_30 = _rdata_T_28 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _rdata_T_31 = {_rdata_T_30,axi_RDATA}; // @[Cat.scala 33:92]
  wire [63:0] _GEN_40 = 2'h1 == servicing_instruction[13:12] ? _rdata_T_23 : _rdata_T_13; // @[peripheralHandler.scala 77:{13,13}]
  wire [63:0] _rdata_WIRE_2_3 = {{32'd0}, axi_RDATA}; // @[peripheralHandler.scala 83:{16,16}]
  wire [63:0] _rdata_T_33 = {32'h0,axi_RDATA}; // @[Cat.scala 33:92]
  reg [63:0] wdata; // @[peripheralHandler.scala 95:18]
  reg [3:0] wstrb; // @[peripheralHandler.scala 96:18]
  wire [4:0] _GEN_47 = 2'h1 == servicing_address[1:0] ? 5'h8 : 5'h0; // @[peripheralHandler.scala 103:{27,27}]
  wire [4:0] _GEN_48 = 2'h2 == servicing_address[1:0] ? 5'h10 : _GEN_47; // @[peripheralHandler.scala 103:{27,27}]
  wire [4:0] _GEN_49 = 2'h3 == servicing_address[1:0] ? 5'h18 : _GEN_48; // @[peripheralHandler.scala 103:{27,27}]
  wire [94:0] _GEN_80 = {{31'd0}, writeIn_data}; // @[peripheralHandler.scala 103:27]
  wire [94:0] _wdata_T_1 = _GEN_80 << _GEN_49; // @[peripheralHandler.scala 103:27]
  wire [3:0] _GEN_51 = 2'h1 == servicing_instruction[13:12] ? 4'h3 : 4'h1; // @[peripheralHandler.scala 105:{75,75}]
  wire [3:0] _GEN_52 = 2'h2 == servicing_instruction[13:12] ? 4'hf : _GEN_51; // @[peripheralHandler.scala 105:{75,75}]
  wire [3:0] _GEN_53 = 2'h3 == servicing_instruction[13:12] ? 4'hf : _GEN_52; // @[peripheralHandler.scala 105:{75,75}]
  wire [6:0] _GEN_81 = {{3'd0}, _GEN_53}; // @[peripheralHandler.scala 105:75]
  wire [6:0] _wstrb_T_2 = _GEN_81 << servicing_address[1:0]; // @[peripheralHandler.scala 105:75]
  wire  _GEN_54 = servicing_instruction[13:12] != 2'h3 | wlast; // @[peripheralHandler.scala 107:{49,57} 17:71]
  wire [94:0] _GEN_55 = writeIn_valid ? _wdata_T_1 : {{31'd0}, wdata}; // @[peripheralHandler.scala 102:23 103:11 95:18]
  wire  _GEN_56 = writeIn_valid | wvalid; // @[peripheralHandler.scala 102:23 104:12 17:71]
  wire [6:0] _GEN_57 = writeIn_valid ? _wstrb_T_2 : {{3'd0}, wstrb}; // @[peripheralHandler.scala 102:23 105:11 96:18]
  wire  _GEN_58 = writeIn_valid | writeCleared; // @[peripheralHandler.scala 102:23 106:18 30:29]
  wire  _GEN_59 = writeIn_valid ? _GEN_54 : wlast; // @[peripheralHandler.scala 102:23 17:71]
  wire  _GEN_60 = axi_AWVALID & axi_AWREADY ? 1'h0 : _GEN_16; // @[peripheralHandler.scala 110:36 111:13]
  wire  _GEN_62 = axi_AWVALID & axi_AWREADY | bready; // @[peripheralHandler.scala 110:36 113:12 17:71]
  wire  _T_20 = axi_WVALID & axi_WREADY; // @[peripheralHandler.scala 116:19]
  wire  _GEN_63 = _T_20 | _GEN_59; // @[peripheralHandler.scala 119:40 120:11]
  wire [94:0] _GEN_64 = _T_20 ? {{63'd0}, wdata[63:32]} : _GEN_55; // @[peripheralHandler.scala 119:40 121:11]
  wire [94:0] _GEN_67 = axi_WVALID & axi_WREADY & axi_WLAST ? _GEN_55 : _GEN_64; // @[peripheralHandler.scala 116:47]
  wire  _GEN_69 = axi_BREADY & axi_BVALID ? 1'h0 : _GEN_24; // @[peripheralHandler.scala 124:34 126:21]
  wire [3:0] _T_25 = servicing_branchMask & branchOps_branchMask; // @[peripheralHandler.scala 130:32]
  wire  _T_26 = |_T_25; // @[peripheralHandler.scala 130:56]
  wire [3:0] _servicing_branchMask_T_1 = servicing_branchMask ^ branchOps_branchMask; // @[peripheralHandler.scala 131:52]
  wire [1:0] _axi_ARSIZE_T_3 = _T_15 ? 2'h2 : servicing_instruction[13:12]; // @[peripheralHandler.scala 149:21]
  assign finishedRequest_valid = servicing_valid; // @[peripheralHandler.scala 15:19]
  assign finishedRequest_address = servicing_address; // @[peripheralHandler.scala 15:19]
  assign finishedRequest_instruction = servicing_instruction; // @[peripheralHandler.scala 15:19]
  assign finishedRequest_robAddr = servicing_robAddr; // @[peripheralHandler.scala 15:19]
  assign finishedRequest_prfDest = servicing_prfDest; // @[peripheralHandler.scala 15:19]
  assign ready = ~(arvalid | rready | awvalid | wvalid | bready | stall); // @[peripheralHandler.scala 20:12]
  assign axi_AWADDR = servicing_address; // @[peripheralHandler.scala 151:15]
  assign axi_AWLEN = {{7'd0}, _T_15}; // @[peripheralHandler.scala 155:15]
  assign axi_AWSIZE = {{1'd0}, _axi_ARSIZE_T_3}; // @[peripheralHandler.scala 159:15]
  assign axi_AWVALID = awvalid & writeCleared; // @[peripheralHandler.scala 160:26]
  assign axi_WDATA = wdata[31:0]; // @[peripheralHandler.scala 163:23]
  assign axi_WSTRB = wstrb; // @[peripheralHandler.scala 165:15]
  assign axi_WLAST = wlast; // @[peripheralHandler.scala 164:15]
  assign axi_WVALID = wvalid; // @[peripheralHandler.scala 166:15]
  assign axi_BREADY = bready; // @[peripheralHandler.scala 161:15]
  assign axi_ARADDR = servicing_address; // @[peripheralHandler.scala 141:15]
  assign axi_ARLEN = {{7'd0}, _T_15}; // @[peripheralHandler.scala 145:15]
  assign axi_ARSIZE = {{1'd0}, _axi_ARSIZE_T_3}; // @[peripheralHandler.scala 149:15]
  assign axi_ARVALID = arvalid & ~(|servicing_branchMask); // @[peripheralHandler.scala 150:26]
  assign axi_RREADY = rready; // @[peripheralHandler.scala 162:15]
  assign readFinished_ready = stall; // @[peripheralHandler.scala 63:22]
  assign readDataOut = rdata; // @[peripheralHandler.scala 71:15]
  always @(posedge clock) begin
    if (reset) begin // @[peripheralHandler.scala 12:26]
      servicing_valid <= 1'h0; // @[peripheralHandler.scala 12:26]
    end else if (branchOps_valid & servicing_valid) begin // @[peripheralHandler.scala 129:44]
      if (_T_5 & _T_26) begin // @[peripheralHandler.scala 133:82]
        servicing_valid <= 1'h0; // @[peripheralHandler.scala 134:23]
      end else begin
        servicing_valid <= _GEN_69;
      end
    end else begin
      servicing_valid <= _GEN_69;
    end
    if (request_valid & ready) begin // @[peripheralHandler.scala 32:32]
      servicing_address <= request_address; // @[peripheralHandler.scala 33:15]
    end
    if (request_valid & ready) begin // @[peripheralHandler.scala 32:32]
      servicing_instruction <= request_instruction; // @[peripheralHandler.scala 33:15]
    end
    if (branchOps_valid & servicing_valid) begin // @[peripheralHandler.scala 129:44]
      if (|_T_25) begin // @[peripheralHandler.scala 130:61]
        servicing_branchMask <= _servicing_branchMask_T_1; // @[peripheralHandler.scala 131:28]
      end else begin
        servicing_branchMask <= _GEN_13;
      end
    end else begin
      servicing_branchMask <= _GEN_13;
    end
    if (request_valid & ready) begin // @[peripheralHandler.scala 32:32]
      servicing_robAddr <= request_robAddr; // @[peripheralHandler.scala 33:15]
    end
    if (request_valid & ready) begin // @[peripheralHandler.scala 32:32]
      servicing_prfDest <= request_prfDest; // @[peripheralHandler.scala 33:15]
    end
    if (reset) begin // @[peripheralHandler.scala 17:71]
      arvalid <= 1'h0; // @[peripheralHandler.scala 17:71]
    end else if (branchOps_valid & servicing_valid) begin // @[peripheralHandler.scala 129:44]
      if (_T_5 & _T_26) begin // @[peripheralHandler.scala 133:82]
        arvalid <= 1'h0; // @[peripheralHandler.scala 137:15]
      end else begin
        arvalid <= _GEN_18;
      end
    end else begin
      arvalid <= _GEN_18;
    end
    if (reset) begin // @[peripheralHandler.scala 17:71]
      rready <= 1'h0; // @[peripheralHandler.scala 17:71]
    end else if (axi_RVALID & axi_RREADY & axi_RLAST) begin // @[peripheralHandler.scala 55:47]
      rready <= 1'h0; // @[peripheralHandler.scala 56:12]
    end else begin
      rready <= _GEN_19;
    end
    if (reset) begin // @[peripheralHandler.scala 17:71]
      awvalid <= 1'h0; // @[peripheralHandler.scala 17:71]
    end else if (branchOps_valid & servicing_valid) begin // @[peripheralHandler.scala 129:44]
      if (_T_5 & _T_26) begin // @[peripheralHandler.scala 133:82]
        awvalid <= 1'h0; // @[peripheralHandler.scala 135:15]
      end else begin
        awvalid <= _GEN_60;
      end
    end else begin
      awvalid <= _GEN_60;
    end
    if (reset) begin // @[peripheralHandler.scala 17:71]
      wvalid <= 1'h0; // @[peripheralHandler.scala 17:71]
    end else if (axi_WVALID & axi_WREADY & axi_WLAST) begin // @[peripheralHandler.scala 116:47]
      wvalid <= 1'h0; // @[peripheralHandler.scala 117:12]
    end else begin
      wvalid <= _GEN_56;
    end
    if (reset) begin // @[peripheralHandler.scala 17:71]
      wlast <= 1'h0; // @[peripheralHandler.scala 17:71]
    end else if (axi_WVALID & axi_WREADY & axi_WLAST) begin // @[peripheralHandler.scala 116:47]
      wlast <= 1'h0; // @[peripheralHandler.scala 118:11]
    end else begin
      wlast <= _GEN_63;
    end
    if (reset) begin // @[peripheralHandler.scala 17:71]
      bready <= 1'h0; // @[peripheralHandler.scala 17:71]
    end else if (axi_BREADY & axi_BVALID) begin // @[peripheralHandler.scala 124:34]
      bready <= 1'h0; // @[peripheralHandler.scala 125:12]
    end else begin
      bready <= _GEN_62;
    end
    if (reset) begin // @[peripheralHandler.scala 17:71]
      stall <= 1'h0; // @[peripheralHandler.scala 17:71]
    end else if (branchOps_valid & servicing_valid) begin // @[peripheralHandler.scala 129:44]
      if (_T_5 & _T_26) begin // @[peripheralHandler.scala 133:82]
        stall <= 1'h0; // @[peripheralHandler.scala 136:13]
      end else begin
        stall <= _GEN_23;
      end
    end else begin
      stall <= _GEN_23;
    end
    if (_T_11) begin // @[peripheralHandler.scala 73:47]
      if (servicing_instruction[13:12] == 2'h3) begin // @[peripheralHandler.scala 74:49]
        rdata <= _rdata_T_1; // @[peripheralHandler.scala 75:13]
      end else if (2'h3 == servicing_instruction[13:12]) begin // @[peripheralHandler.scala 77:13]
        rdata <= _rdata_WIRE_2_3; // @[peripheralHandler.scala 77:13]
      end else if (2'h2 == servicing_instruction[13:12]) begin // @[peripheralHandler.scala 77:13]
        rdata <= _rdata_T_31; // @[peripheralHandler.scala 77:13]
      end else begin
        rdata <= _GEN_40;
      end
    end else if (_T_10) begin // @[peripheralHandler.scala 91:40]
      rdata <= _rdata_T_33; // @[peripheralHandler.scala 92:11]
    end
    if (reset) begin // @[peripheralHandler.scala 30:29]
      writeCleared <= 1'h0; // @[peripheralHandler.scala 30:29]
    end else if (axi_AWVALID & axi_AWREADY) begin // @[peripheralHandler.scala 110:36]
      writeCleared <= 1'h0; // @[peripheralHandler.scala 112:18]
    end else begin
      writeCleared <= _GEN_58;
    end
    wdata <= _GEN_67[63:0];
    wstrb <= _GEN_57[3:0];
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  servicing_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  servicing_address = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  servicing_instruction = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  servicing_branchMask = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  servicing_robAddr = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  servicing_prfDest = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  arvalid = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  rready = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  awvalid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  wvalid = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  wlast = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  bready = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  stall = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  rdata = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  writeCleared = _RAND_14[0:0];
  _RAND_15 = {2{`RANDOM}};
  wdata = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  wstrb = _RAND_16[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module zeroWriteLatencyCache(
  input         clock,
  input         reset,
  input  [31:0] readAddress,
  output [63:0] readOut_0_data,
  output [19:0] readOut_0_tag,
  output        readOut_0_valid,
  output [63:0] readOut_1_data,
  output [19:0] readOut_1_tag,
  output        readOut_1_valid,
  input         writePorts_0_enable,
  input  [31:0] writePorts_0_cacheAddress,
  input  [63:0] writePorts_0_data,
  input         writePorts_1_enable,
  input  [31:0] writePorts_1_cacheAddress,
  input  [63:0] writePorts_1_data,
  input         invalidateSet_valid,
  input  [5:0]  invalidateSet_cacheIndex,
  input         invalidateSet_invalidateVector_0,
  input         invalidateSet_invalidateVector_1,
  input         cacheFillDone_valid,
  input  [5:0]  cacheFillDone_cacheIndex,
  input         cacheFillDone_validateVector_0,
  input         cacheFillDone_validateVector_1,
  input  [19:0] cacheFillDone_tag
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [63:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [31:0] _RAND_145;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] cacheSets_0 [0:511]; // @[writeToReadNoLatencyBRAM.scala 11:60]
  wire  cacheSets_0_readOut_0_data_MPORT_en; // @[writeToReadNoLatencyBRAM.scala 11:60]
  wire [8:0] cacheSets_0_readOut_0_data_MPORT_addr; // @[writeToReadNoLatencyBRAM.scala 11:60]
  wire [63:0] cacheSets_0_readOut_0_data_MPORT_data; // @[writeToReadNoLatencyBRAM.scala 11:60]
  wire [63:0] cacheSets_0_MPORT_data; // @[writeToReadNoLatencyBRAM.scala 11:60]
  wire [8:0] cacheSets_0_MPORT_addr; // @[writeToReadNoLatencyBRAM.scala 11:60]
  wire  cacheSets_0_MPORT_mask; // @[writeToReadNoLatencyBRAM.scala 11:60]
  wire  cacheSets_0_MPORT_en; // @[writeToReadNoLatencyBRAM.scala 11:60]
  reg  cacheSets_0_readOut_0_data_MPORT_en_pipe_0;
  reg [8:0] cacheSets_0_readOut_0_data_MPORT_addr_pipe_0;
  reg [63:0] cacheSets_1 [0:511]; // @[writeToReadNoLatencyBRAM.scala 11:60]
  wire  cacheSets_1_readOut_1_data_MPORT_en; // @[writeToReadNoLatencyBRAM.scala 11:60]
  wire [8:0] cacheSets_1_readOut_1_data_MPORT_addr; // @[writeToReadNoLatencyBRAM.scala 11:60]
  wire [63:0] cacheSets_1_readOut_1_data_MPORT_data; // @[writeToReadNoLatencyBRAM.scala 11:60]
  wire [63:0] cacheSets_1_MPORT_1_data; // @[writeToReadNoLatencyBRAM.scala 11:60]
  wire [8:0] cacheSets_1_MPORT_1_addr; // @[writeToReadNoLatencyBRAM.scala 11:60]
  wire  cacheSets_1_MPORT_1_mask; // @[writeToReadNoLatencyBRAM.scala 11:60]
  wire  cacheSets_1_MPORT_1_en; // @[writeToReadNoLatencyBRAM.scala 11:60]
  reg  cacheSets_1_readOut_1_data_MPORT_en_pipe_0;
  reg [8:0] cacheSets_1_readOut_1_data_MPORT_addr_pipe_0;
  reg [19:0] tags_0 [0:63]; // @[writeToReadNoLatencyBRAM.scala 12:55]
  wire  tags_0_readOut_0_tag_MPORT_en; // @[writeToReadNoLatencyBRAM.scala 12:55]
  wire [5:0] tags_0_readOut_0_tag_MPORT_addr; // @[writeToReadNoLatencyBRAM.scala 12:55]
  wire [19:0] tags_0_readOut_0_tag_MPORT_data; // @[writeToReadNoLatencyBRAM.scala 12:55]
  wire [19:0] tags_0_MPORT_2_data; // @[writeToReadNoLatencyBRAM.scala 12:55]
  wire [5:0] tags_0_MPORT_2_addr; // @[writeToReadNoLatencyBRAM.scala 12:55]
  wire  tags_0_MPORT_2_mask; // @[writeToReadNoLatencyBRAM.scala 12:55]
  wire  tags_0_MPORT_2_en; // @[writeToReadNoLatencyBRAM.scala 12:55]
  reg  tags_0_readOut_0_tag_MPORT_en_pipe_0;
  reg [5:0] tags_0_readOut_0_tag_MPORT_addr_pipe_0;
  reg [19:0] tags_1 [0:63]; // @[writeToReadNoLatencyBRAM.scala 12:55]
  wire  tags_1_readOut_1_tag_MPORT_en; // @[writeToReadNoLatencyBRAM.scala 12:55]
  wire [5:0] tags_1_readOut_1_tag_MPORT_addr; // @[writeToReadNoLatencyBRAM.scala 12:55]
  wire [19:0] tags_1_readOut_1_tag_MPORT_data; // @[writeToReadNoLatencyBRAM.scala 12:55]
  wire [19:0] tags_1_MPORT_3_data; // @[writeToReadNoLatencyBRAM.scala 12:55]
  wire [5:0] tags_1_MPORT_3_addr; // @[writeToReadNoLatencyBRAM.scala 12:55]
  wire  tags_1_MPORT_3_mask; // @[writeToReadNoLatencyBRAM.scala 12:55]
  wire  tags_1_MPORT_3_en; // @[writeToReadNoLatencyBRAM.scala 12:55]
  reg  tags_1_readOut_1_tag_MPORT_en_pipe_0;
  reg [5:0] tags_1_readOut_1_tag_MPORT_addr_pipe_0;
  reg  validBits_0_0; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_1; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_2; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_3; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_4; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_5; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_6; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_7; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_8; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_9; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_10; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_11; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_12; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_13; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_14; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_15; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_16; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_17; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_18; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_19; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_20; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_21; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_22; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_23; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_24; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_25; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_26; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_27; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_28; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_29; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_30; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_31; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_32; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_33; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_34; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_35; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_36; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_37; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_38; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_39; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_40; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_41; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_42; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_43; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_44; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_45; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_46; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_47; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_48; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_49; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_50; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_51; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_52; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_53; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_54; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_55; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_56; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_57; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_58; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_59; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_60; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_61; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_62; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_0_63; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_0; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_1; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_2; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_3; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_4; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_5; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_6; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_7; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_8; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_9; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_10; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_11; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_12; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_13; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_14; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_15; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_16; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_17; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_18; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_19; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_20; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_21; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_22; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_23; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_24; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_25; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_26; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_27; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_28; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_29; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_30; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_31; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_32; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_33; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_34; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_35; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_36; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_37; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_38; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_39; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_40; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_41; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_42; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_43; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_44; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_45; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_46; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_47; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_48; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_49; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_50; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_51; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_52; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_53; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_54; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_55; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_56; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_57; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_58; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_59; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_60; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_61; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_62; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  validBits_1_63; // @[writeToReadNoLatencyBRAM.scala 34:56]
  reg  doForward; // @[writeToReadNoLatencyBRAM.scala 40:28]
  reg [63:0] readOut_0_data_REG; // @[writeToReadNoLatencyBRAM.scala 42:40]
  reg  readOut_0_valid_REG; // @[writeToReadNoLatencyBRAM.scala 44:26]
  wire  _GEN_17 = 6'h1 == readAddress[11:6] ? validBits_0_1 : validBits_0_0; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_18 = 6'h2 == readAddress[11:6] ? validBits_0_2 : _GEN_17; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_19 = 6'h3 == readAddress[11:6] ? validBits_0_3 : _GEN_18; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_20 = 6'h4 == readAddress[11:6] ? validBits_0_4 : _GEN_19; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_21 = 6'h5 == readAddress[11:6] ? validBits_0_5 : _GEN_20; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_22 = 6'h6 == readAddress[11:6] ? validBits_0_6 : _GEN_21; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_23 = 6'h7 == readAddress[11:6] ? validBits_0_7 : _GEN_22; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_24 = 6'h8 == readAddress[11:6] ? validBits_0_8 : _GEN_23; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_25 = 6'h9 == readAddress[11:6] ? validBits_0_9 : _GEN_24; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_26 = 6'ha == readAddress[11:6] ? validBits_0_10 : _GEN_25; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_27 = 6'hb == readAddress[11:6] ? validBits_0_11 : _GEN_26; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_28 = 6'hc == readAddress[11:6] ? validBits_0_12 : _GEN_27; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_29 = 6'hd == readAddress[11:6] ? validBits_0_13 : _GEN_28; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_30 = 6'he == readAddress[11:6] ? validBits_0_14 : _GEN_29; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_31 = 6'hf == readAddress[11:6] ? validBits_0_15 : _GEN_30; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_32 = 6'h10 == readAddress[11:6] ? validBits_0_16 : _GEN_31; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_33 = 6'h11 == readAddress[11:6] ? validBits_0_17 : _GEN_32; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_34 = 6'h12 == readAddress[11:6] ? validBits_0_18 : _GEN_33; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_35 = 6'h13 == readAddress[11:6] ? validBits_0_19 : _GEN_34; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_36 = 6'h14 == readAddress[11:6] ? validBits_0_20 : _GEN_35; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_37 = 6'h15 == readAddress[11:6] ? validBits_0_21 : _GEN_36; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_38 = 6'h16 == readAddress[11:6] ? validBits_0_22 : _GEN_37; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_39 = 6'h17 == readAddress[11:6] ? validBits_0_23 : _GEN_38; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_40 = 6'h18 == readAddress[11:6] ? validBits_0_24 : _GEN_39; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_41 = 6'h19 == readAddress[11:6] ? validBits_0_25 : _GEN_40; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_42 = 6'h1a == readAddress[11:6] ? validBits_0_26 : _GEN_41; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_43 = 6'h1b == readAddress[11:6] ? validBits_0_27 : _GEN_42; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_44 = 6'h1c == readAddress[11:6] ? validBits_0_28 : _GEN_43; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_45 = 6'h1d == readAddress[11:6] ? validBits_0_29 : _GEN_44; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_46 = 6'h1e == readAddress[11:6] ? validBits_0_30 : _GEN_45; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_47 = 6'h1f == readAddress[11:6] ? validBits_0_31 : _GEN_46; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_48 = 6'h20 == readAddress[11:6] ? validBits_0_32 : _GEN_47; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_49 = 6'h21 == readAddress[11:6] ? validBits_0_33 : _GEN_48; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_50 = 6'h22 == readAddress[11:6] ? validBits_0_34 : _GEN_49; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_51 = 6'h23 == readAddress[11:6] ? validBits_0_35 : _GEN_50; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_52 = 6'h24 == readAddress[11:6] ? validBits_0_36 : _GEN_51; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_53 = 6'h25 == readAddress[11:6] ? validBits_0_37 : _GEN_52; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_54 = 6'h26 == readAddress[11:6] ? validBits_0_38 : _GEN_53; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_55 = 6'h27 == readAddress[11:6] ? validBits_0_39 : _GEN_54; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_56 = 6'h28 == readAddress[11:6] ? validBits_0_40 : _GEN_55; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_57 = 6'h29 == readAddress[11:6] ? validBits_0_41 : _GEN_56; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_58 = 6'h2a == readAddress[11:6] ? validBits_0_42 : _GEN_57; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_59 = 6'h2b == readAddress[11:6] ? validBits_0_43 : _GEN_58; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_60 = 6'h2c == readAddress[11:6] ? validBits_0_44 : _GEN_59; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_61 = 6'h2d == readAddress[11:6] ? validBits_0_45 : _GEN_60; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_62 = 6'h2e == readAddress[11:6] ? validBits_0_46 : _GEN_61; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_63 = 6'h2f == readAddress[11:6] ? validBits_0_47 : _GEN_62; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_64 = 6'h30 == readAddress[11:6] ? validBits_0_48 : _GEN_63; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_65 = 6'h31 == readAddress[11:6] ? validBits_0_49 : _GEN_64; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_66 = 6'h32 == readAddress[11:6] ? validBits_0_50 : _GEN_65; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_67 = 6'h33 == readAddress[11:6] ? validBits_0_51 : _GEN_66; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_68 = 6'h34 == readAddress[11:6] ? validBits_0_52 : _GEN_67; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_69 = 6'h35 == readAddress[11:6] ? validBits_0_53 : _GEN_68; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_70 = 6'h36 == readAddress[11:6] ? validBits_0_54 : _GEN_69; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_71 = 6'h37 == readAddress[11:6] ? validBits_0_55 : _GEN_70; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_72 = 6'h38 == readAddress[11:6] ? validBits_0_56 : _GEN_71; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_73 = 6'h39 == readAddress[11:6] ? validBits_0_57 : _GEN_72; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_74 = 6'h3a == readAddress[11:6] ? validBits_0_58 : _GEN_73; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_75 = 6'h3b == readAddress[11:6] ? validBits_0_59 : _GEN_74; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  reg  doForward_1; // @[writeToReadNoLatencyBRAM.scala 40:28]
  reg [63:0] readOut_1_data_REG; // @[writeToReadNoLatencyBRAM.scala 42:40]
  reg  readOut_1_valid_REG; // @[writeToReadNoLatencyBRAM.scala 44:26]
  wire  _GEN_85 = 6'h1 == readAddress[11:6] ? validBits_1_1 : validBits_1_0; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_86 = 6'h2 == readAddress[11:6] ? validBits_1_2 : _GEN_85; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_87 = 6'h3 == readAddress[11:6] ? validBits_1_3 : _GEN_86; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_88 = 6'h4 == readAddress[11:6] ? validBits_1_4 : _GEN_87; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_89 = 6'h5 == readAddress[11:6] ? validBits_1_5 : _GEN_88; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_90 = 6'h6 == readAddress[11:6] ? validBits_1_6 : _GEN_89; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_91 = 6'h7 == readAddress[11:6] ? validBits_1_7 : _GEN_90; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_92 = 6'h8 == readAddress[11:6] ? validBits_1_8 : _GEN_91; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_93 = 6'h9 == readAddress[11:6] ? validBits_1_9 : _GEN_92; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_94 = 6'ha == readAddress[11:6] ? validBits_1_10 : _GEN_93; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_95 = 6'hb == readAddress[11:6] ? validBits_1_11 : _GEN_94; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_96 = 6'hc == readAddress[11:6] ? validBits_1_12 : _GEN_95; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_97 = 6'hd == readAddress[11:6] ? validBits_1_13 : _GEN_96; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_98 = 6'he == readAddress[11:6] ? validBits_1_14 : _GEN_97; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_99 = 6'hf == readAddress[11:6] ? validBits_1_15 : _GEN_98; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_100 = 6'h10 == readAddress[11:6] ? validBits_1_16 : _GEN_99; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_101 = 6'h11 == readAddress[11:6] ? validBits_1_17 : _GEN_100; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_102 = 6'h12 == readAddress[11:6] ? validBits_1_18 : _GEN_101; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_103 = 6'h13 == readAddress[11:6] ? validBits_1_19 : _GEN_102; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_104 = 6'h14 == readAddress[11:6] ? validBits_1_20 : _GEN_103; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_105 = 6'h15 == readAddress[11:6] ? validBits_1_21 : _GEN_104; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_106 = 6'h16 == readAddress[11:6] ? validBits_1_22 : _GEN_105; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_107 = 6'h17 == readAddress[11:6] ? validBits_1_23 : _GEN_106; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_108 = 6'h18 == readAddress[11:6] ? validBits_1_24 : _GEN_107; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_109 = 6'h19 == readAddress[11:6] ? validBits_1_25 : _GEN_108; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_110 = 6'h1a == readAddress[11:6] ? validBits_1_26 : _GEN_109; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_111 = 6'h1b == readAddress[11:6] ? validBits_1_27 : _GEN_110; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_112 = 6'h1c == readAddress[11:6] ? validBits_1_28 : _GEN_111; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_113 = 6'h1d == readAddress[11:6] ? validBits_1_29 : _GEN_112; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_114 = 6'h1e == readAddress[11:6] ? validBits_1_30 : _GEN_113; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_115 = 6'h1f == readAddress[11:6] ? validBits_1_31 : _GEN_114; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_116 = 6'h20 == readAddress[11:6] ? validBits_1_32 : _GEN_115; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_117 = 6'h21 == readAddress[11:6] ? validBits_1_33 : _GEN_116; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_118 = 6'h22 == readAddress[11:6] ? validBits_1_34 : _GEN_117; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_119 = 6'h23 == readAddress[11:6] ? validBits_1_35 : _GEN_118; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_120 = 6'h24 == readAddress[11:6] ? validBits_1_36 : _GEN_119; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_121 = 6'h25 == readAddress[11:6] ? validBits_1_37 : _GEN_120; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_122 = 6'h26 == readAddress[11:6] ? validBits_1_38 : _GEN_121; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_123 = 6'h27 == readAddress[11:6] ? validBits_1_39 : _GEN_122; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_124 = 6'h28 == readAddress[11:6] ? validBits_1_40 : _GEN_123; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_125 = 6'h29 == readAddress[11:6] ? validBits_1_41 : _GEN_124; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_126 = 6'h2a == readAddress[11:6] ? validBits_1_42 : _GEN_125; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_127 = 6'h2b == readAddress[11:6] ? validBits_1_43 : _GEN_126; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_128 = 6'h2c == readAddress[11:6] ? validBits_1_44 : _GEN_127; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_129 = 6'h2d == readAddress[11:6] ? validBits_1_45 : _GEN_128; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_130 = 6'h2e == readAddress[11:6] ? validBits_1_46 : _GEN_129; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_131 = 6'h2f == readAddress[11:6] ? validBits_1_47 : _GEN_130; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_132 = 6'h30 == readAddress[11:6] ? validBits_1_48 : _GEN_131; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_133 = 6'h31 == readAddress[11:6] ? validBits_1_49 : _GEN_132; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_134 = 6'h32 == readAddress[11:6] ? validBits_1_50 : _GEN_133; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_135 = 6'h33 == readAddress[11:6] ? validBits_1_51 : _GEN_134; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_136 = 6'h34 == readAddress[11:6] ? validBits_1_52 : _GEN_135; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_137 = 6'h35 == readAddress[11:6] ? validBits_1_53 : _GEN_136; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_138 = 6'h36 == readAddress[11:6] ? validBits_1_54 : _GEN_137; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_139 = 6'h37 == readAddress[11:6] ? validBits_1_55 : _GEN_138; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_140 = 6'h38 == readAddress[11:6] ? validBits_1_56 : _GEN_139; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_141 = 6'h39 == readAddress[11:6] ? validBits_1_57 : _GEN_140; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_142 = 6'h3a == readAddress[11:6] ? validBits_1_58 : _GEN_141; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_143 = 6'h3b == readAddress[11:6] ? validBits_1_59 : _GEN_142; // @[writeToReadNoLatencyBRAM.scala 44:{26,26}]
  wire  _GEN_148 = 6'h0 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_0; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_149 = 6'h1 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_1; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_150 = 6'h2 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_2; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_151 = 6'h3 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_3; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_152 = 6'h4 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_4; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_153 = 6'h5 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_5; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_154 = 6'h6 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_6; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_155 = 6'h7 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_7; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_156 = 6'h8 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_8; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_157 = 6'h9 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_9; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_158 = 6'ha == invalidateSet_cacheIndex ? 1'h0 : validBits_0_10; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_159 = 6'hb == invalidateSet_cacheIndex ? 1'h0 : validBits_0_11; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_160 = 6'hc == invalidateSet_cacheIndex ? 1'h0 : validBits_0_12; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_161 = 6'hd == invalidateSet_cacheIndex ? 1'h0 : validBits_0_13; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_162 = 6'he == invalidateSet_cacheIndex ? 1'h0 : validBits_0_14; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_163 = 6'hf == invalidateSet_cacheIndex ? 1'h0 : validBits_0_15; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_164 = 6'h10 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_16; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_165 = 6'h11 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_17; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_166 = 6'h12 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_18; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_167 = 6'h13 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_19; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_168 = 6'h14 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_20; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_169 = 6'h15 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_21; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_170 = 6'h16 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_22; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_171 = 6'h17 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_23; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_172 = 6'h18 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_24; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_173 = 6'h19 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_25; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_174 = 6'h1a == invalidateSet_cacheIndex ? 1'h0 : validBits_0_26; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_175 = 6'h1b == invalidateSet_cacheIndex ? 1'h0 : validBits_0_27; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_176 = 6'h1c == invalidateSet_cacheIndex ? 1'h0 : validBits_0_28; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_177 = 6'h1d == invalidateSet_cacheIndex ? 1'h0 : validBits_0_29; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_178 = 6'h1e == invalidateSet_cacheIndex ? 1'h0 : validBits_0_30; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_179 = 6'h1f == invalidateSet_cacheIndex ? 1'h0 : validBits_0_31; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_180 = 6'h20 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_32; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_181 = 6'h21 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_33; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_182 = 6'h22 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_34; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_183 = 6'h23 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_35; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_184 = 6'h24 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_36; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_185 = 6'h25 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_37; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_186 = 6'h26 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_38; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_187 = 6'h27 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_39; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_188 = 6'h28 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_40; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_189 = 6'h29 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_41; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_190 = 6'h2a == invalidateSet_cacheIndex ? 1'h0 : validBits_0_42; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_191 = 6'h2b == invalidateSet_cacheIndex ? 1'h0 : validBits_0_43; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_192 = 6'h2c == invalidateSet_cacheIndex ? 1'h0 : validBits_0_44; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_193 = 6'h2d == invalidateSet_cacheIndex ? 1'h0 : validBits_0_45; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_194 = 6'h2e == invalidateSet_cacheIndex ? 1'h0 : validBits_0_46; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_195 = 6'h2f == invalidateSet_cacheIndex ? 1'h0 : validBits_0_47; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_196 = 6'h30 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_48; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_197 = 6'h31 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_49; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_198 = 6'h32 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_50; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_199 = 6'h33 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_51; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_200 = 6'h34 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_52; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_201 = 6'h35 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_53; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_202 = 6'h36 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_54; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_203 = 6'h37 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_55; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_204 = 6'h38 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_56; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_205 = 6'h39 == invalidateSet_cacheIndex ? 1'h0 : validBits_0_57; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_206 = 6'h3a == invalidateSet_cacheIndex ? 1'h0 : validBits_0_58; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_207 = 6'h3b == invalidateSet_cacheIndex ? 1'h0 : validBits_0_59; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_208 = 6'h3c == invalidateSet_cacheIndex ? 1'h0 : validBits_0_60; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_209 = 6'h3d == invalidateSet_cacheIndex ? 1'h0 : validBits_0_61; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_210 = 6'h3e == invalidateSet_cacheIndex ? 1'h0 : validBits_0_62; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_211 = 6'h3f == invalidateSet_cacheIndex ? 1'h0 : validBits_0_63; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_212 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_148 : validBits_0_0; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_213 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_149 : validBits_0_1; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_214 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_150 : validBits_0_2; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_215 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_151 : validBits_0_3; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_216 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_152 : validBits_0_4; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_217 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_153 : validBits_0_5; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_218 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_154 : validBits_0_6; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_219 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_155 : validBits_0_7; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_220 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_156 : validBits_0_8; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_221 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_157 : validBits_0_9; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_222 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_158 : validBits_0_10; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_223 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_159 : validBits_0_11; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_224 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_160 : validBits_0_12; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_225 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_161 : validBits_0_13; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_226 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_162 : validBits_0_14; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_227 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_163 : validBits_0_15; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_228 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_164 : validBits_0_16; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_229 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_165 : validBits_0_17; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_230 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_166 : validBits_0_18; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_231 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_167 : validBits_0_19; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_232 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_168 : validBits_0_20; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_233 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_169 : validBits_0_21; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_234 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_170 : validBits_0_22; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_235 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_171 : validBits_0_23; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_236 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_172 : validBits_0_24; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_237 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_173 : validBits_0_25; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_238 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_174 : validBits_0_26; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_239 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_175 : validBits_0_27; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_240 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_176 : validBits_0_28; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_241 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_177 : validBits_0_29; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_242 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_178 : validBits_0_30; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_243 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_179 : validBits_0_31; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_244 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_180 : validBits_0_32; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_245 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_181 : validBits_0_33; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_246 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_182 : validBits_0_34; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_247 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_183 : validBits_0_35; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_248 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_184 : validBits_0_36; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_249 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_185 : validBits_0_37; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_250 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_186 : validBits_0_38; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_251 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_187 : validBits_0_39; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_252 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_188 : validBits_0_40; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_253 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_189 : validBits_0_41; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_254 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_190 : validBits_0_42; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_255 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_191 : validBits_0_43; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_256 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_192 : validBits_0_44; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_257 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_193 : validBits_0_45; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_258 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_194 : validBits_0_46; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_259 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_195 : validBits_0_47; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_260 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_196 : validBits_0_48; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_261 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_197 : validBits_0_49; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_262 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_198 : validBits_0_50; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_263 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_199 : validBits_0_51; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_264 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_200 : validBits_0_52; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_265 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_201 : validBits_0_53; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_266 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_202 : validBits_0_54; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_267 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_203 : validBits_0_55; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_268 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_204 : validBits_0_56; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_269 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_205 : validBits_0_57; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_270 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_206 : validBits_0_58; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_271 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_207 : validBits_0_59; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_272 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_208 : validBits_0_60; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_273 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_209 : validBits_0_61; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_274 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_210 : validBits_0_62; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_275 = invalidateSet_valid & invalidateSet_invalidateVector_0 ? _GEN_211 : validBits_0_63; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_276 = 6'h0 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_0; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_277 = 6'h1 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_1; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_278 = 6'h2 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_2; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_279 = 6'h3 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_3; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_280 = 6'h4 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_4; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_281 = 6'h5 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_5; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_282 = 6'h6 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_6; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_283 = 6'h7 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_7; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_284 = 6'h8 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_8; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_285 = 6'h9 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_9; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_286 = 6'ha == invalidateSet_cacheIndex ? 1'h0 : validBits_1_10; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_287 = 6'hb == invalidateSet_cacheIndex ? 1'h0 : validBits_1_11; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_288 = 6'hc == invalidateSet_cacheIndex ? 1'h0 : validBits_1_12; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_289 = 6'hd == invalidateSet_cacheIndex ? 1'h0 : validBits_1_13; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_290 = 6'he == invalidateSet_cacheIndex ? 1'h0 : validBits_1_14; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_291 = 6'hf == invalidateSet_cacheIndex ? 1'h0 : validBits_1_15; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_292 = 6'h10 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_16; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_293 = 6'h11 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_17; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_294 = 6'h12 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_18; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_295 = 6'h13 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_19; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_296 = 6'h14 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_20; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_297 = 6'h15 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_21; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_298 = 6'h16 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_22; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_299 = 6'h17 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_23; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_300 = 6'h18 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_24; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_301 = 6'h19 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_25; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_302 = 6'h1a == invalidateSet_cacheIndex ? 1'h0 : validBits_1_26; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_303 = 6'h1b == invalidateSet_cacheIndex ? 1'h0 : validBits_1_27; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_304 = 6'h1c == invalidateSet_cacheIndex ? 1'h0 : validBits_1_28; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_305 = 6'h1d == invalidateSet_cacheIndex ? 1'h0 : validBits_1_29; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_306 = 6'h1e == invalidateSet_cacheIndex ? 1'h0 : validBits_1_30; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_307 = 6'h1f == invalidateSet_cacheIndex ? 1'h0 : validBits_1_31; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_308 = 6'h20 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_32; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_309 = 6'h21 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_33; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_310 = 6'h22 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_34; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_311 = 6'h23 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_35; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_312 = 6'h24 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_36; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_313 = 6'h25 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_37; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_314 = 6'h26 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_38; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_315 = 6'h27 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_39; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_316 = 6'h28 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_40; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_317 = 6'h29 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_41; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_318 = 6'h2a == invalidateSet_cacheIndex ? 1'h0 : validBits_1_42; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_319 = 6'h2b == invalidateSet_cacheIndex ? 1'h0 : validBits_1_43; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_320 = 6'h2c == invalidateSet_cacheIndex ? 1'h0 : validBits_1_44; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_321 = 6'h2d == invalidateSet_cacheIndex ? 1'h0 : validBits_1_45; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_322 = 6'h2e == invalidateSet_cacheIndex ? 1'h0 : validBits_1_46; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_323 = 6'h2f == invalidateSet_cacheIndex ? 1'h0 : validBits_1_47; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_324 = 6'h30 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_48; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_325 = 6'h31 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_49; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_326 = 6'h32 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_50; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_327 = 6'h33 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_51; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_328 = 6'h34 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_52; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_329 = 6'h35 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_53; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_330 = 6'h36 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_54; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_331 = 6'h37 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_55; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_332 = 6'h38 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_56; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_333 = 6'h39 == invalidateSet_cacheIndex ? 1'h0 : validBits_1_57; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_334 = 6'h3a == invalidateSet_cacheIndex ? 1'h0 : validBits_1_58; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_335 = 6'h3b == invalidateSet_cacheIndex ? 1'h0 : validBits_1_59; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_336 = 6'h3c == invalidateSet_cacheIndex ? 1'h0 : validBits_1_60; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_337 = 6'h3d == invalidateSet_cacheIndex ? 1'h0 : validBits_1_61; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_338 = 6'h3e == invalidateSet_cacheIndex ? 1'h0 : validBits_1_62; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_339 = 6'h3f == invalidateSet_cacheIndex ? 1'h0 : validBits_1_63; // @[writeToReadNoLatencyBRAM.scala 34:56 54:{82,82}]
  wire  _GEN_340 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_276 : validBits_1_0; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_341 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_277 : validBits_1_1; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_342 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_278 : validBits_1_2; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_343 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_279 : validBits_1_3; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_344 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_280 : validBits_1_4; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_345 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_281 : validBits_1_5; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_346 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_282 : validBits_1_6; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_347 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_283 : validBits_1_7; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_348 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_284 : validBits_1_8; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_349 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_285 : validBits_1_9; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_350 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_286 : validBits_1_10; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_351 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_287 : validBits_1_11; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_352 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_288 : validBits_1_12; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_353 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_289 : validBits_1_13; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_354 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_290 : validBits_1_14; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_355 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_291 : validBits_1_15; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_356 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_292 : validBits_1_16; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_357 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_293 : validBits_1_17; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_358 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_294 : validBits_1_18; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_359 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_295 : validBits_1_19; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_360 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_296 : validBits_1_20; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_361 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_297 : validBits_1_21; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_362 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_298 : validBits_1_22; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_363 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_299 : validBits_1_23; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_364 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_300 : validBits_1_24; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_365 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_301 : validBits_1_25; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_366 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_302 : validBits_1_26; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_367 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_303 : validBits_1_27; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_368 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_304 : validBits_1_28; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_369 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_305 : validBits_1_29; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_370 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_306 : validBits_1_30; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_371 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_307 : validBits_1_31; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_372 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_308 : validBits_1_32; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_373 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_309 : validBits_1_33; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_374 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_310 : validBits_1_34; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_375 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_311 : validBits_1_35; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_376 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_312 : validBits_1_36; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_377 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_313 : validBits_1_37; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_378 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_314 : validBits_1_38; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_379 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_315 : validBits_1_39; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_380 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_316 : validBits_1_40; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_381 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_317 : validBits_1_41; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_382 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_318 : validBits_1_42; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_383 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_319 : validBits_1_43; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_384 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_320 : validBits_1_44; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_385 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_321 : validBits_1_45; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_386 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_322 : validBits_1_46; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_387 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_323 : validBits_1_47; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_388 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_324 : validBits_1_48; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_389 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_325 : validBits_1_49; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_390 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_326 : validBits_1_50; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_391 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_327 : validBits_1_51; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_392 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_328 : validBits_1_52; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_393 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_329 : validBits_1_53; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_394 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_330 : validBits_1_54; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_395 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_331 : validBits_1_55; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_396 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_332 : validBits_1_56; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_397 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_333 : validBits_1_57; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_398 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_334 : validBits_1_58; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_399 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_335 : validBits_1_59; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_400 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_336 : validBits_1_60; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_401 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_337 : validBits_1_61; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_402 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_338 : validBits_1_62; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_403 = invalidateSet_valid & invalidateSet_invalidateVector_1 ? _GEN_339 : validBits_1_63; // @[writeToReadNoLatencyBRAM.scala 54:45 34:56]
  wire  _GEN_404 = 6'h0 == cacheFillDone_cacheIndex | _GEN_212; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_405 = 6'h1 == cacheFillDone_cacheIndex | _GEN_213; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_406 = 6'h2 == cacheFillDone_cacheIndex | _GEN_214; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_407 = 6'h3 == cacheFillDone_cacheIndex | _GEN_215; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_408 = 6'h4 == cacheFillDone_cacheIndex | _GEN_216; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_409 = 6'h5 == cacheFillDone_cacheIndex | _GEN_217; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_410 = 6'h6 == cacheFillDone_cacheIndex | _GEN_218; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_411 = 6'h7 == cacheFillDone_cacheIndex | _GEN_219; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_412 = 6'h8 == cacheFillDone_cacheIndex | _GEN_220; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_413 = 6'h9 == cacheFillDone_cacheIndex | _GEN_221; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_414 = 6'ha == cacheFillDone_cacheIndex | _GEN_222; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_415 = 6'hb == cacheFillDone_cacheIndex | _GEN_223; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_416 = 6'hc == cacheFillDone_cacheIndex | _GEN_224; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_417 = 6'hd == cacheFillDone_cacheIndex | _GEN_225; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_418 = 6'he == cacheFillDone_cacheIndex | _GEN_226; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_419 = 6'hf == cacheFillDone_cacheIndex | _GEN_227; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_420 = 6'h10 == cacheFillDone_cacheIndex | _GEN_228; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_421 = 6'h11 == cacheFillDone_cacheIndex | _GEN_229; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_422 = 6'h12 == cacheFillDone_cacheIndex | _GEN_230; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_423 = 6'h13 == cacheFillDone_cacheIndex | _GEN_231; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_424 = 6'h14 == cacheFillDone_cacheIndex | _GEN_232; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_425 = 6'h15 == cacheFillDone_cacheIndex | _GEN_233; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_426 = 6'h16 == cacheFillDone_cacheIndex | _GEN_234; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_427 = 6'h17 == cacheFillDone_cacheIndex | _GEN_235; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_428 = 6'h18 == cacheFillDone_cacheIndex | _GEN_236; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_429 = 6'h19 == cacheFillDone_cacheIndex | _GEN_237; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_430 = 6'h1a == cacheFillDone_cacheIndex | _GEN_238; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_431 = 6'h1b == cacheFillDone_cacheIndex | _GEN_239; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_432 = 6'h1c == cacheFillDone_cacheIndex | _GEN_240; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_433 = 6'h1d == cacheFillDone_cacheIndex | _GEN_241; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_434 = 6'h1e == cacheFillDone_cacheIndex | _GEN_242; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_435 = 6'h1f == cacheFillDone_cacheIndex | _GEN_243; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_436 = 6'h20 == cacheFillDone_cacheIndex | _GEN_244; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_437 = 6'h21 == cacheFillDone_cacheIndex | _GEN_245; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_438 = 6'h22 == cacheFillDone_cacheIndex | _GEN_246; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_439 = 6'h23 == cacheFillDone_cacheIndex | _GEN_247; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_440 = 6'h24 == cacheFillDone_cacheIndex | _GEN_248; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_441 = 6'h25 == cacheFillDone_cacheIndex | _GEN_249; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_442 = 6'h26 == cacheFillDone_cacheIndex | _GEN_250; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_443 = 6'h27 == cacheFillDone_cacheIndex | _GEN_251; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_444 = 6'h28 == cacheFillDone_cacheIndex | _GEN_252; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_445 = 6'h29 == cacheFillDone_cacheIndex | _GEN_253; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_446 = 6'h2a == cacheFillDone_cacheIndex | _GEN_254; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_447 = 6'h2b == cacheFillDone_cacheIndex | _GEN_255; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_448 = 6'h2c == cacheFillDone_cacheIndex | _GEN_256; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_449 = 6'h2d == cacheFillDone_cacheIndex | _GEN_257; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_450 = 6'h2e == cacheFillDone_cacheIndex | _GEN_258; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_451 = 6'h2f == cacheFillDone_cacheIndex | _GEN_259; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_452 = 6'h30 == cacheFillDone_cacheIndex | _GEN_260; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_453 = 6'h31 == cacheFillDone_cacheIndex | _GEN_261; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_454 = 6'h32 == cacheFillDone_cacheIndex | _GEN_262; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_455 = 6'h33 == cacheFillDone_cacheIndex | _GEN_263; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_456 = 6'h34 == cacheFillDone_cacheIndex | _GEN_264; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_457 = 6'h35 == cacheFillDone_cacheIndex | _GEN_265; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_458 = 6'h36 == cacheFillDone_cacheIndex | _GEN_266; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_459 = 6'h37 == cacheFillDone_cacheIndex | _GEN_267; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_460 = 6'h38 == cacheFillDone_cacheIndex | _GEN_268; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_461 = 6'h39 == cacheFillDone_cacheIndex | _GEN_269; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_462 = 6'h3a == cacheFillDone_cacheIndex | _GEN_270; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_463 = 6'h3b == cacheFillDone_cacheIndex | _GEN_271; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_464 = 6'h3c == cacheFillDone_cacheIndex | _GEN_272; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_465 = 6'h3d == cacheFillDone_cacheIndex | _GEN_273; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_466 = 6'h3e == cacheFillDone_cacheIndex | _GEN_274; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_467 = 6'h3f == cacheFillDone_cacheIndex | _GEN_275; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_537 = 6'h0 == cacheFillDone_cacheIndex | _GEN_340; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_538 = 6'h1 == cacheFillDone_cacheIndex | _GEN_341; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_539 = 6'h2 == cacheFillDone_cacheIndex | _GEN_342; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_540 = 6'h3 == cacheFillDone_cacheIndex | _GEN_343; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_541 = 6'h4 == cacheFillDone_cacheIndex | _GEN_344; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_542 = 6'h5 == cacheFillDone_cacheIndex | _GEN_345; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_543 = 6'h6 == cacheFillDone_cacheIndex | _GEN_346; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_544 = 6'h7 == cacheFillDone_cacheIndex | _GEN_347; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_545 = 6'h8 == cacheFillDone_cacheIndex | _GEN_348; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_546 = 6'h9 == cacheFillDone_cacheIndex | _GEN_349; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_547 = 6'ha == cacheFillDone_cacheIndex | _GEN_350; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_548 = 6'hb == cacheFillDone_cacheIndex | _GEN_351; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_549 = 6'hc == cacheFillDone_cacheIndex | _GEN_352; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_550 = 6'hd == cacheFillDone_cacheIndex | _GEN_353; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_551 = 6'he == cacheFillDone_cacheIndex | _GEN_354; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_552 = 6'hf == cacheFillDone_cacheIndex | _GEN_355; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_553 = 6'h10 == cacheFillDone_cacheIndex | _GEN_356; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_554 = 6'h11 == cacheFillDone_cacheIndex | _GEN_357; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_555 = 6'h12 == cacheFillDone_cacheIndex | _GEN_358; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_556 = 6'h13 == cacheFillDone_cacheIndex | _GEN_359; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_557 = 6'h14 == cacheFillDone_cacheIndex | _GEN_360; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_558 = 6'h15 == cacheFillDone_cacheIndex | _GEN_361; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_559 = 6'h16 == cacheFillDone_cacheIndex | _GEN_362; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_560 = 6'h17 == cacheFillDone_cacheIndex | _GEN_363; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_561 = 6'h18 == cacheFillDone_cacheIndex | _GEN_364; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_562 = 6'h19 == cacheFillDone_cacheIndex | _GEN_365; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_563 = 6'h1a == cacheFillDone_cacheIndex | _GEN_366; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_564 = 6'h1b == cacheFillDone_cacheIndex | _GEN_367; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_565 = 6'h1c == cacheFillDone_cacheIndex | _GEN_368; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_566 = 6'h1d == cacheFillDone_cacheIndex | _GEN_369; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_567 = 6'h1e == cacheFillDone_cacheIndex | _GEN_370; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_568 = 6'h1f == cacheFillDone_cacheIndex | _GEN_371; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_569 = 6'h20 == cacheFillDone_cacheIndex | _GEN_372; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_570 = 6'h21 == cacheFillDone_cacheIndex | _GEN_373; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_571 = 6'h22 == cacheFillDone_cacheIndex | _GEN_374; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_572 = 6'h23 == cacheFillDone_cacheIndex | _GEN_375; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_573 = 6'h24 == cacheFillDone_cacheIndex | _GEN_376; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_574 = 6'h25 == cacheFillDone_cacheIndex | _GEN_377; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_575 = 6'h26 == cacheFillDone_cacheIndex | _GEN_378; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_576 = 6'h27 == cacheFillDone_cacheIndex | _GEN_379; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_577 = 6'h28 == cacheFillDone_cacheIndex | _GEN_380; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_578 = 6'h29 == cacheFillDone_cacheIndex | _GEN_381; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_579 = 6'h2a == cacheFillDone_cacheIndex | _GEN_382; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_580 = 6'h2b == cacheFillDone_cacheIndex | _GEN_383; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_581 = 6'h2c == cacheFillDone_cacheIndex | _GEN_384; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_582 = 6'h2d == cacheFillDone_cacheIndex | _GEN_385; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_583 = 6'h2e == cacheFillDone_cacheIndex | _GEN_386; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_584 = 6'h2f == cacheFillDone_cacheIndex | _GEN_387; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_585 = 6'h30 == cacheFillDone_cacheIndex | _GEN_388; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_586 = 6'h31 == cacheFillDone_cacheIndex | _GEN_389; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_587 = 6'h32 == cacheFillDone_cacheIndex | _GEN_390; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_588 = 6'h33 == cacheFillDone_cacheIndex | _GEN_391; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_589 = 6'h34 == cacheFillDone_cacheIndex | _GEN_392; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_590 = 6'h35 == cacheFillDone_cacheIndex | _GEN_393; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_591 = 6'h36 == cacheFillDone_cacheIndex | _GEN_394; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_592 = 6'h37 == cacheFillDone_cacheIndex | _GEN_395; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_593 = 6'h38 == cacheFillDone_cacheIndex | _GEN_396; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_594 = 6'h39 == cacheFillDone_cacheIndex | _GEN_397; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_595 = 6'h3a == cacheFillDone_cacheIndex | _GEN_398; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_596 = 6'h3b == cacheFillDone_cacheIndex | _GEN_399; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_597 = 6'h3c == cacheFillDone_cacheIndex | _GEN_400; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_598 = 6'h3d == cacheFillDone_cacheIndex | _GEN_401; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_599 = 6'h3e == cacheFillDone_cacheIndex | _GEN_402; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  wire  _GEN_600 = 6'h3f == cacheFillDone_cacheIndex | _GEN_403; // @[writeToReadNoLatencyBRAM.scala 66:{42,42}]
  assign cacheSets_0_readOut_0_data_MPORT_en = cacheSets_0_readOut_0_data_MPORT_en_pipe_0;
  assign cacheSets_0_readOut_0_data_MPORT_addr = cacheSets_0_readOut_0_data_MPORT_addr_pipe_0;
  assign cacheSets_0_readOut_0_data_MPORT_data = cacheSets_0[cacheSets_0_readOut_0_data_MPORT_addr]; // @[writeToReadNoLatencyBRAM.scala 11:60]
  assign cacheSets_0_MPORT_data = writePorts_0_data;
  assign cacheSets_0_MPORT_addr = writePorts_0_cacheAddress[11:3];
  assign cacheSets_0_MPORT_mask = 1'h1;
  assign cacheSets_0_MPORT_en = writePorts_0_enable;
  assign cacheSets_1_readOut_1_data_MPORT_en = cacheSets_1_readOut_1_data_MPORT_en_pipe_0;
  assign cacheSets_1_readOut_1_data_MPORT_addr = cacheSets_1_readOut_1_data_MPORT_addr_pipe_0;
  assign cacheSets_1_readOut_1_data_MPORT_data = cacheSets_1[cacheSets_1_readOut_1_data_MPORT_addr]; // @[writeToReadNoLatencyBRAM.scala 11:60]
  assign cacheSets_1_MPORT_1_data = writePorts_1_data;
  assign cacheSets_1_MPORT_1_addr = writePorts_1_cacheAddress[11:3];
  assign cacheSets_1_MPORT_1_mask = 1'h1;
  assign cacheSets_1_MPORT_1_en = writePorts_1_enable;
  assign tags_0_readOut_0_tag_MPORT_en = tags_0_readOut_0_tag_MPORT_en_pipe_0;
  assign tags_0_readOut_0_tag_MPORT_addr = tags_0_readOut_0_tag_MPORT_addr_pipe_0;
  assign tags_0_readOut_0_tag_MPORT_data = tags_0[tags_0_readOut_0_tag_MPORT_addr]; // @[writeToReadNoLatencyBRAM.scala 12:55]
  assign tags_0_MPORT_2_data = cacheFillDone_tag;
  assign tags_0_MPORT_2_addr = cacheFillDone_cacheIndex;
  assign tags_0_MPORT_2_mask = 1'h1;
  assign tags_0_MPORT_2_en = cacheFillDone_valid & cacheFillDone_validateVector_0;
  assign tags_1_readOut_1_tag_MPORT_en = tags_1_readOut_1_tag_MPORT_en_pipe_0;
  assign tags_1_readOut_1_tag_MPORT_addr = tags_1_readOut_1_tag_MPORT_addr_pipe_0;
  assign tags_1_readOut_1_tag_MPORT_data = tags_1[tags_1_readOut_1_tag_MPORT_addr]; // @[writeToReadNoLatencyBRAM.scala 12:55]
  assign tags_1_MPORT_3_data = cacheFillDone_tag;
  assign tags_1_MPORT_3_addr = cacheFillDone_cacheIndex;
  assign tags_1_MPORT_3_mask = 1'h1;
  assign tags_1_MPORT_3_en = cacheFillDone_valid & cacheFillDone_validateVector_1;
  assign readOut_0_data = doForward ? readOut_0_data_REG : cacheSets_0_readOut_0_data_MPORT_data; // @[writeToReadNoLatencyBRAM.scala 42:21]
  assign readOut_0_tag = tags_0_readOut_0_tag_MPORT_data; // @[writeToReadNoLatencyBRAM.scala 43:14]
  assign readOut_0_valid = readOut_0_valid_REG; // @[writeToReadNoLatencyBRAM.scala 44:16]
  assign readOut_1_data = doForward_1 ? readOut_1_data_REG : cacheSets_1_readOut_1_data_MPORT_data; // @[writeToReadNoLatencyBRAM.scala 42:21]
  assign readOut_1_tag = tags_1_readOut_1_tag_MPORT_data; // @[writeToReadNoLatencyBRAM.scala 43:14]
  assign readOut_1_valid = readOut_1_valid_REG; // @[writeToReadNoLatencyBRAM.scala 44:16]
  always @(posedge clock) begin
    if (cacheSets_0_MPORT_en & cacheSets_0_MPORT_mask) begin
      cacheSets_0[cacheSets_0_MPORT_addr] <= cacheSets_0_MPORT_data; // @[writeToReadNoLatencyBRAM.scala 11:60]
    end
    cacheSets_0_readOut_0_data_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheSets_0_readOut_0_data_MPORT_addr_pipe_0 <= readAddress[11:3];
    end
    if (cacheSets_1_MPORT_1_en & cacheSets_1_MPORT_1_mask) begin
      cacheSets_1[cacheSets_1_MPORT_1_addr] <= cacheSets_1_MPORT_1_data; // @[writeToReadNoLatencyBRAM.scala 11:60]
    end
    cacheSets_1_readOut_1_data_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      cacheSets_1_readOut_1_data_MPORT_addr_pipe_0 <= readAddress[11:3];
    end
    if (tags_0_MPORT_2_en & tags_0_MPORT_2_mask) begin
      tags_0[tags_0_MPORT_2_addr] <= tags_0_MPORT_2_data; // @[writeToReadNoLatencyBRAM.scala 12:55]
    end
    tags_0_readOut_0_tag_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      tags_0_readOut_0_tag_MPORT_addr_pipe_0 <= readAddress[11:6];
    end
    if (tags_1_MPORT_3_en & tags_1_MPORT_3_mask) begin
      tags_1[tags_1_MPORT_3_addr] <= tags_1_MPORT_3_data; // @[writeToReadNoLatencyBRAM.scala 12:55]
    end
    tags_1_readOut_1_tag_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      tags_1_readOut_1_tag_MPORT_addr_pipe_0 <= readAddress[11:6];
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_0 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_0 <= _GEN_404;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h0 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_0 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_1 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_1 <= _GEN_405;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h1 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_1 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_2 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_2 <= _GEN_406;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h2 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_2 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_3 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_3 <= _GEN_407;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h3 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_3 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_4 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_4 <= _GEN_408;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h4 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_4 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_5 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_5 <= _GEN_409;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h5 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_5 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_6 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_6 <= _GEN_410;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h6 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_6 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_7 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_7 <= _GEN_411;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h7 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_7 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_8 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_8 <= _GEN_412;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h8 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_8 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_9 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_9 <= _GEN_413;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h9 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_9 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_10 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_10 <= _GEN_414;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'ha == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_10 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_11 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_11 <= _GEN_415;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'hb == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_11 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_12 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_12 <= _GEN_416;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'hc == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_12 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_13 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_13 <= _GEN_417;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'hd == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_13 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_14 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_14 <= _GEN_418;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'he == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_14 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_15 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_15 <= _GEN_419;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'hf == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_15 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_16 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_16 <= _GEN_420;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h10 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_16 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_17 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_17 <= _GEN_421;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h11 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_17 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_18 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_18 <= _GEN_422;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h12 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_18 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_19 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_19 <= _GEN_423;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h13 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_19 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_20 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_20 <= _GEN_424;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h14 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_20 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_21 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_21 <= _GEN_425;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h15 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_21 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_22 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_22 <= _GEN_426;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h16 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_22 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_23 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_23 <= _GEN_427;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h17 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_23 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_24 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_24 <= _GEN_428;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h18 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_24 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_25 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_25 <= _GEN_429;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h19 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_25 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_26 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_26 <= _GEN_430;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h1a == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_26 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_27 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_27 <= _GEN_431;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h1b == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_27 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_28 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_28 <= _GEN_432;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h1c == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_28 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_29 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_29 <= _GEN_433;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h1d == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_29 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_30 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_30 <= _GEN_434;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h1e == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_30 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_31 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_31 <= _GEN_435;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h1f == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_31 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_32 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_32 <= _GEN_436;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h20 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_32 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_33 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_33 <= _GEN_437;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h21 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_33 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_34 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_34 <= _GEN_438;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h22 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_34 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_35 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_35 <= _GEN_439;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h23 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_35 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_36 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_36 <= _GEN_440;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h24 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_36 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_37 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_37 <= _GEN_441;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h25 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_37 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_38 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_38 <= _GEN_442;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h26 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_38 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_39 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_39 <= _GEN_443;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h27 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_39 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_40 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_40 <= _GEN_444;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h28 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_40 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_41 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_41 <= _GEN_445;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h29 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_41 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_42 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_42 <= _GEN_446;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h2a == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_42 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_43 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_43 <= _GEN_447;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h2b == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_43 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_44 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_44 <= _GEN_448;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h2c == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_44 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_45 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_45 <= _GEN_449;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h2d == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_45 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_46 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_46 <= _GEN_450;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h2e == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_46 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_47 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_47 <= _GEN_451;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h2f == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_47 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_48 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_48 <= _GEN_452;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h30 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_48 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_49 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_49 <= _GEN_453;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h31 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_49 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_50 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_50 <= _GEN_454;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h32 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_50 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_51 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_51 <= _GEN_455;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h33 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_51 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_52 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_52 <= _GEN_456;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h34 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_52 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_53 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_53 <= _GEN_457;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h35 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_53 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_54 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_54 <= _GEN_458;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h36 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_54 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_55 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_55 <= _GEN_459;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h37 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_55 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_56 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_56 <= _GEN_460;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h38 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_56 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_57 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_57 <= _GEN_461;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h39 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_57 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_58 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_58 <= _GEN_462;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h3a == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_58 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_59 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_59 <= _GEN_463;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h3b == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_59 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_60 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_60 <= _GEN_464;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h3c == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_60 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_61 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_61 <= _GEN_465;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h3d == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_61 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_62 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_62 <= _GEN_466;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h3e == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_62 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_0_63 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_0_63 <= _GEN_467;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_0) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h3f == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_0_63 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_0 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_0 <= _GEN_537;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h0 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_0 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_1 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_1 <= _GEN_538;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h1 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_1 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_2 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_2 <= _GEN_539;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h2 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_2 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_3 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_3 <= _GEN_540;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h3 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_3 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_4 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_4 <= _GEN_541;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h4 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_4 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_5 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_5 <= _GEN_542;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h5 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_5 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_6 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_6 <= _GEN_543;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h6 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_6 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_7 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_7 <= _GEN_544;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h7 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_7 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_8 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_8 <= _GEN_545;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h8 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_8 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_9 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_9 <= _GEN_546;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h9 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_9 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_10 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_10 <= _GEN_547;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'ha == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_10 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_11 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_11 <= _GEN_548;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'hb == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_11 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_12 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_12 <= _GEN_549;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'hc == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_12 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_13 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_13 <= _GEN_550;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'hd == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_13 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_14 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_14 <= _GEN_551;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'he == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_14 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_15 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_15 <= _GEN_552;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'hf == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_15 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_16 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_16 <= _GEN_553;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h10 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_16 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_17 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_17 <= _GEN_554;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h11 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_17 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_18 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_18 <= _GEN_555;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h12 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_18 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_19 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_19 <= _GEN_556;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h13 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_19 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_20 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_20 <= _GEN_557;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h14 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_20 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_21 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_21 <= _GEN_558;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h15 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_21 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_22 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_22 <= _GEN_559;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h16 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_22 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_23 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_23 <= _GEN_560;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h17 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_23 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_24 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_24 <= _GEN_561;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h18 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_24 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_25 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_25 <= _GEN_562;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h19 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_25 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_26 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_26 <= _GEN_563;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h1a == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_26 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_27 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_27 <= _GEN_564;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h1b == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_27 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_28 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_28 <= _GEN_565;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h1c == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_28 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_29 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_29 <= _GEN_566;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h1d == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_29 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_30 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_30 <= _GEN_567;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h1e == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_30 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_31 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_31 <= _GEN_568;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h1f == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_31 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_32 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_32 <= _GEN_569;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h20 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_32 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_33 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_33 <= _GEN_570;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h21 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_33 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_34 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_34 <= _GEN_571;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h22 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_34 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_35 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_35 <= _GEN_572;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h23 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_35 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_36 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_36 <= _GEN_573;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h24 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_36 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_37 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_37 <= _GEN_574;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h25 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_37 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_38 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_38 <= _GEN_575;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h26 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_38 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_39 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_39 <= _GEN_576;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h27 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_39 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_40 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_40 <= _GEN_577;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h28 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_40 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_41 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_41 <= _GEN_578;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h29 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_41 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_42 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_42 <= _GEN_579;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h2a == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_42 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_43 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_43 <= _GEN_580;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h2b == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_43 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_44 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_44 <= _GEN_581;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h2c == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_44 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_45 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_45 <= _GEN_582;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h2d == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_45 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_46 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_46 <= _GEN_583;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h2e == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_46 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_47 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_47 <= _GEN_584;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h2f == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_47 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_48 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_48 <= _GEN_585;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h30 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_48 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_49 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_49 <= _GEN_586;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h31 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_49 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_50 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_50 <= _GEN_587;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h32 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_50 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_51 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_51 <= _GEN_588;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h33 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_51 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_52 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_52 <= _GEN_589;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h34 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_52 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_53 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_53 <= _GEN_590;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h35 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_53 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_54 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_54 <= _GEN_591;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h36 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_54 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_55 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_55 <= _GEN_592;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h37 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_55 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_56 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_56 <= _GEN_593;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h38 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_56 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_57 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_57 <= _GEN_594;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h39 == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_57 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_58 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_58 <= _GEN_595;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h3a == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_58 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_59 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_59 <= _GEN_596;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h3b == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_59 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_60 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_60 <= _GEN_597;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h3c == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_60 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_61 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_61 <= _GEN_598;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h3d == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_61 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_62 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_62 <= _GEN_599;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h3e == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_62 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    if (reset) begin // @[writeToReadNoLatencyBRAM.scala 34:56]
      validBits_1_63 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 34:56]
    end else if (cacheFillDone_valid & cacheFillDone_validateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 65:43]
      validBits_1_63 <= _GEN_600;
    end else if (invalidateSet_valid & invalidateSet_invalidateVector_1) begin // @[writeToReadNoLatencyBRAM.scala 54:45]
      if (6'h3f == invalidateSet_cacheIndex) begin // @[writeToReadNoLatencyBRAM.scala 54:82]
        validBits_1_63 <= 1'h0; // @[writeToReadNoLatencyBRAM.scala 54:82]
      end
    end
    doForward <= readAddress[31:2] == writePorts_0_cacheAddress[31:2] & writePorts_0_enable; // @[writeToReadNoLatencyBRAM.scala 40:78]
    readOut_0_data_REG <= writePorts_0_data; // @[writeToReadNoLatencyBRAM.scala 42:40]
    if (6'h3f == readAddress[11:6]) begin // @[writeToReadNoLatencyBRAM.scala 44:26]
      readOut_0_valid_REG <= validBits_0_63; // @[writeToReadNoLatencyBRAM.scala 44:26]
    end else if (6'h3e == readAddress[11:6]) begin // @[writeToReadNoLatencyBRAM.scala 44:26]
      readOut_0_valid_REG <= validBits_0_62; // @[writeToReadNoLatencyBRAM.scala 44:26]
    end else if (6'h3d == readAddress[11:6]) begin // @[writeToReadNoLatencyBRAM.scala 44:26]
      readOut_0_valid_REG <= validBits_0_61; // @[writeToReadNoLatencyBRAM.scala 44:26]
    end else if (6'h3c == readAddress[11:6]) begin // @[writeToReadNoLatencyBRAM.scala 44:26]
      readOut_0_valid_REG <= validBits_0_60; // @[writeToReadNoLatencyBRAM.scala 44:26]
    end else begin
      readOut_0_valid_REG <= _GEN_75;
    end
    doForward_1 <= readAddress[31:2] == writePorts_1_cacheAddress[31:2] & writePorts_1_enable; // @[writeToReadNoLatencyBRAM.scala 40:78]
    readOut_1_data_REG <= writePorts_1_data; // @[writeToReadNoLatencyBRAM.scala 42:40]
    if (6'h3f == readAddress[11:6]) begin // @[writeToReadNoLatencyBRAM.scala 44:26]
      readOut_1_valid_REG <= validBits_1_63; // @[writeToReadNoLatencyBRAM.scala 44:26]
    end else if (6'h3e == readAddress[11:6]) begin // @[writeToReadNoLatencyBRAM.scala 44:26]
      readOut_1_valid_REG <= validBits_1_62; // @[writeToReadNoLatencyBRAM.scala 44:26]
    end else if (6'h3d == readAddress[11:6]) begin // @[writeToReadNoLatencyBRAM.scala 44:26]
      readOut_1_valid_REG <= validBits_1_61; // @[writeToReadNoLatencyBRAM.scala 44:26]
    end else if (6'h3c == readAddress[11:6]) begin // @[writeToReadNoLatencyBRAM.scala 44:26]
      readOut_1_valid_REG <= validBits_1_60; // @[writeToReadNoLatencyBRAM.scala 44:26]
    end else begin
      readOut_1_valid_REG <= _GEN_143;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    cacheSets_0[initvar] = _RAND_0[63:0];
  _RAND_3 = {2{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    cacheSets_1[initvar] = _RAND_3[63:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tags_0[initvar] = _RAND_6[19:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tags_1[initvar] = _RAND_9[19:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cacheSets_0_readOut_0_data_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  cacheSets_0_readOut_0_data_MPORT_addr_pipe_0 = _RAND_2[8:0];
  _RAND_4 = {1{`RANDOM}};
  cacheSets_1_readOut_1_data_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cacheSets_1_readOut_1_data_MPORT_addr_pipe_0 = _RAND_5[8:0];
  _RAND_7 = {1{`RANDOM}};
  tags_0_readOut_0_tag_MPORT_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  tags_0_readOut_0_tag_MPORT_addr_pipe_0 = _RAND_8[5:0];
  _RAND_10 = {1{`RANDOM}};
  tags_1_readOut_1_tag_MPORT_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  tags_1_readOut_1_tag_MPORT_addr_pipe_0 = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  validBits_0_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  validBits_0_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  validBits_0_2 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  validBits_0_3 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  validBits_0_4 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  validBits_0_5 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  validBits_0_6 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  validBits_0_7 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  validBits_0_8 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  validBits_0_9 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  validBits_0_10 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  validBits_0_11 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  validBits_0_12 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  validBits_0_13 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  validBits_0_14 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  validBits_0_15 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  validBits_0_16 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  validBits_0_17 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  validBits_0_18 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  validBits_0_19 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  validBits_0_20 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  validBits_0_21 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  validBits_0_22 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  validBits_0_23 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  validBits_0_24 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  validBits_0_25 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  validBits_0_26 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  validBits_0_27 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  validBits_0_28 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  validBits_0_29 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  validBits_0_30 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  validBits_0_31 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  validBits_0_32 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  validBits_0_33 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  validBits_0_34 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  validBits_0_35 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  validBits_0_36 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  validBits_0_37 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  validBits_0_38 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  validBits_0_39 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  validBits_0_40 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  validBits_0_41 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  validBits_0_42 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  validBits_0_43 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  validBits_0_44 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  validBits_0_45 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  validBits_0_46 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  validBits_0_47 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  validBits_0_48 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  validBits_0_49 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  validBits_0_50 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  validBits_0_51 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  validBits_0_52 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  validBits_0_53 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  validBits_0_54 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  validBits_0_55 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  validBits_0_56 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  validBits_0_57 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  validBits_0_58 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  validBits_0_59 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  validBits_0_60 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  validBits_0_61 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  validBits_0_62 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  validBits_0_63 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  validBits_1_0 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  validBits_1_1 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  validBits_1_2 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  validBits_1_3 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  validBits_1_4 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  validBits_1_5 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  validBits_1_6 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  validBits_1_7 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  validBits_1_8 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  validBits_1_9 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  validBits_1_10 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  validBits_1_11 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  validBits_1_12 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  validBits_1_13 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  validBits_1_14 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  validBits_1_15 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  validBits_1_16 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  validBits_1_17 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  validBits_1_18 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  validBits_1_19 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  validBits_1_20 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  validBits_1_21 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  validBits_1_22 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  validBits_1_23 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  validBits_1_24 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  validBits_1_25 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  validBits_1_26 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  validBits_1_27 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  validBits_1_28 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  validBits_1_29 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  validBits_1_30 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  validBits_1_31 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  validBits_1_32 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  validBits_1_33 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  validBits_1_34 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  validBits_1_35 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  validBits_1_36 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  validBits_1_37 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  validBits_1_38 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  validBits_1_39 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  validBits_1_40 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  validBits_1_41 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  validBits_1_42 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  validBits_1_43 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  validBits_1_44 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  validBits_1_45 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  validBits_1_46 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  validBits_1_47 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  validBits_1_48 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  validBits_1_49 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  validBits_1_50 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  validBits_1_51 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  validBits_1_52 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  validBits_1_53 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  validBits_1_54 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  validBits_1_55 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  validBits_1_56 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  validBits_1_57 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  validBits_1_58 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  validBits_1_59 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  validBits_1_60 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  validBits_1_61 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  validBits_1_62 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  validBits_1_63 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  doForward = _RAND_140[0:0];
  _RAND_141 = {2{`RANDOM}};
  readOut_0_data_REG = _RAND_141[63:0];
  _RAND_142 = {1{`RANDOM}};
  readOut_0_valid_REG = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  doForward_1 = _RAND_143[0:0];
  _RAND_144 = {2{`RANDOM}};
  readOut_1_data_REG = _RAND_144[63:0];
  _RAND_145 = {1{`RANDOM}};
  readOut_1_valid_REG = _RAND_145[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module missHandler(
  input         clock,
  input         reset,
  output        replayOut_query_valid,
  output [31:0] replayOut_query_address,
  output [31:0] replayOut_query_instruction,
  output [3:0]  replayOut_query_branchMask,
  output [3:0]  replayOut_query_robAddr,
  output [5:0]  replayOut_query_prfDest,
  output [63:0] replayOut_data,
  output        replayingQuries,
  input         branchOps_valid,
  input  [3:0]  branchOps_branchMask,
  input         branchOps_passed,
  input         cachePipelineEmpty,
  input         missedRequest_query_valid,
  input  [31:0] missedRequest_query_address,
  input  [31:0] missedRequest_query_instruction,
  input  [3:0]  missedRequest_query_branchMask,
  input  [3:0]  missedRequest_query_robAddr,
  input  [5:0]  missedRequest_query_prfDest,
  input  [63:0] missedRequest_data,
  output        pushToCache_ready,
  input         pushToCache_fired,
  output [63:0] pushToCache_cacheWriteOut_data,
  output [8:0]  pushToCache_cacheWriteOut_address,
  output [1:0]  pushToCache_cacheWriteOut_setSelVector,
  output [31:0] axi_ARADDR,
  output        axi_ARVALID,
  input         axi_ARREADY,
  input  [31:0] axi_RDATA,
  input         axi_RLAST,
  input         axi_RVALID,
  output        axi_RREADY,
  output        dependencyCheck_requset_valid,
  output [31:0] dependencyCheck_requset_address,
  input         dependencyCheck_free,
  output        rlastToCache,
  output [1:0]  setInvalidateVector,
  input  [1:0]  setFillStatus,
  output        handlerBusy,
  output        handlerSaturated,
  output        clean,
  output        nonSaturatedReplay
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
`endif // RANDOMIZE_REG_INIT
  reg  saturatedReplayVector_0_query_valid; // @[missHandler.scala 75:38]
  reg [31:0] saturatedReplayVector_0_query_address; // @[missHandler.scala 75:38]
  reg [31:0] saturatedReplayVector_0_query_instruction; // @[missHandler.scala 75:38]
  reg [3:0] saturatedReplayVector_0_query_branchMask; // @[missHandler.scala 75:38]
  reg [3:0] saturatedReplayVector_0_query_robAddr; // @[missHandler.scala 75:38]
  reg [5:0] saturatedReplayVector_0_query_prfDest; // @[missHandler.scala 75:38]
  reg [63:0] saturatedReplayVector_0_data; // @[missHandler.scala 75:38]
  reg  saturatedReplayVector_1_query_valid; // @[missHandler.scala 75:38]
  reg [31:0] saturatedReplayVector_1_query_address; // @[missHandler.scala 75:38]
  reg [31:0] saturatedReplayVector_1_query_instruction; // @[missHandler.scala 75:38]
  reg [3:0] saturatedReplayVector_1_query_branchMask; // @[missHandler.scala 75:38]
  reg [3:0] saturatedReplayVector_1_query_robAddr; // @[missHandler.scala 75:38]
  reg [5:0] saturatedReplayVector_1_query_prfDest; // @[missHandler.scala 75:38]
  reg [63:0] saturatedReplayVector_1_data; // @[missHandler.scala 75:38]
  reg  saturatedReplayVector_2_query_valid; // @[missHandler.scala 75:38]
  reg [31:0] saturatedReplayVector_2_query_address; // @[missHandler.scala 75:38]
  reg [31:0] saturatedReplayVector_2_query_instruction; // @[missHandler.scala 75:38]
  reg [3:0] saturatedReplayVector_2_query_branchMask; // @[missHandler.scala 75:38]
  reg [3:0] saturatedReplayVector_2_query_robAddr; // @[missHandler.scala 75:38]
  reg [5:0] saturatedReplayVector_2_query_prfDest; // @[missHandler.scala 75:38]
  reg [63:0] saturatedReplayVector_2_data; // @[missHandler.scala 75:38]
  reg  saturatedReplayVector_3_query_valid; // @[missHandler.scala 75:38]
  reg [31:0] saturatedReplayVector_3_query_address; // @[missHandler.scala 75:38]
  reg [31:0] saturatedReplayVector_3_query_instruction; // @[missHandler.scala 75:38]
  reg [3:0] saturatedReplayVector_3_query_branchMask; // @[missHandler.scala 75:38]
  reg [3:0] saturatedReplayVector_3_query_robAddr; // @[missHandler.scala 75:38]
  reg [5:0] saturatedReplayVector_3_query_prfDest; // @[missHandler.scala 75:38]
  reg [63:0] saturatedReplayVector_3_data; // @[missHandler.scala 75:38]
  reg  saturatedReplayVector_4_query_valid; // @[missHandler.scala 75:38]
  reg [31:0] saturatedReplayVector_4_query_address; // @[missHandler.scala 75:38]
  reg [31:0] saturatedReplayVector_4_query_instruction; // @[missHandler.scala 75:38]
  reg [3:0] saturatedReplayVector_4_query_branchMask; // @[missHandler.scala 75:38]
  reg [3:0] saturatedReplayVector_4_query_robAddr; // @[missHandler.scala 75:38]
  reg [5:0] saturatedReplayVector_4_query_prfDest; // @[missHandler.scala 75:38]
  reg [63:0] saturatedReplayVector_4_data; // @[missHandler.scala 75:38]
  reg  saturatedCollectVector_0_query_valid; // @[missHandler.scala 81:39]
  reg [31:0] saturatedCollectVector_0_query_address; // @[missHandler.scala 81:39]
  reg [31:0] saturatedCollectVector_0_query_instruction; // @[missHandler.scala 81:39]
  reg [3:0] saturatedCollectVector_0_query_branchMask; // @[missHandler.scala 81:39]
  reg [3:0] saturatedCollectVector_0_query_robAddr; // @[missHandler.scala 81:39]
  reg [5:0] saturatedCollectVector_0_query_prfDest; // @[missHandler.scala 81:39]
  reg [63:0] saturatedCollectVector_0_data; // @[missHandler.scala 81:39]
  reg  saturatedCollectVector_1_query_valid; // @[missHandler.scala 81:39]
  reg [31:0] saturatedCollectVector_1_query_address; // @[missHandler.scala 81:39]
  reg [31:0] saturatedCollectVector_1_query_instruction; // @[missHandler.scala 81:39]
  reg [3:0] saturatedCollectVector_1_query_branchMask; // @[missHandler.scala 81:39]
  reg [3:0] saturatedCollectVector_1_query_robAddr; // @[missHandler.scala 81:39]
  reg [5:0] saturatedCollectVector_1_query_prfDest; // @[missHandler.scala 81:39]
  reg [63:0] saturatedCollectVector_1_data; // @[missHandler.scala 81:39]
  reg  saturatedCollectVector_2_query_valid; // @[missHandler.scala 81:39]
  reg [31:0] saturatedCollectVector_2_query_address; // @[missHandler.scala 81:39]
  reg [31:0] saturatedCollectVector_2_query_instruction; // @[missHandler.scala 81:39]
  reg [3:0] saturatedCollectVector_2_query_branchMask; // @[missHandler.scala 81:39]
  reg [3:0] saturatedCollectVector_2_query_robAddr; // @[missHandler.scala 81:39]
  reg [5:0] saturatedCollectVector_2_query_prfDest; // @[missHandler.scala 81:39]
  reg [63:0] saturatedCollectVector_2_data; // @[missHandler.scala 81:39]
  reg  saturatedCollectVector_3_query_valid; // @[missHandler.scala 81:39]
  reg [31:0] saturatedCollectVector_3_query_address; // @[missHandler.scala 81:39]
  reg [31:0] saturatedCollectVector_3_query_instruction; // @[missHandler.scala 81:39]
  reg [3:0] saturatedCollectVector_3_query_branchMask; // @[missHandler.scala 81:39]
  reg [3:0] saturatedCollectVector_3_query_robAddr; // @[missHandler.scala 81:39]
  reg [5:0] saturatedCollectVector_3_query_prfDest; // @[missHandler.scala 81:39]
  reg [63:0] saturatedCollectVector_3_data; // @[missHandler.scala 81:39]
  reg  saturatedCollectVector_4_query_valid; // @[missHandler.scala 81:39]
  reg [31:0] saturatedCollectVector_4_query_address; // @[missHandler.scala 81:39]
  reg [31:0] saturatedCollectVector_4_query_instruction; // @[missHandler.scala 81:39]
  reg [3:0] saturatedCollectVector_4_query_branchMask; // @[missHandler.scala 81:39]
  reg [3:0] saturatedCollectVector_4_query_robAddr; // @[missHandler.scala 81:39]
  reg [5:0] saturatedCollectVector_4_query_prfDest; // @[missHandler.scala 81:39]
  reg [63:0] saturatedCollectVector_4_data; // @[missHandler.scala 81:39]
  reg  nonSaturatedMisses_0_query_valid; // @[missHandler.scala 83:35]
  reg [31:0] nonSaturatedMisses_0_query_address; // @[missHandler.scala 83:35]
  reg [31:0] nonSaturatedMisses_0_query_instruction; // @[missHandler.scala 83:35]
  reg [3:0] nonSaturatedMisses_0_query_branchMask; // @[missHandler.scala 83:35]
  reg [3:0] nonSaturatedMisses_0_query_robAddr; // @[missHandler.scala 83:35]
  reg [5:0] nonSaturatedMisses_0_query_prfDest; // @[missHandler.scala 83:35]
  reg [63:0] nonSaturatedMisses_0_data; // @[missHandler.scala 83:35]
  reg  nonSaturatedMisses_1_query_valid; // @[missHandler.scala 83:35]
  reg [31:0] nonSaturatedMisses_1_query_address; // @[missHandler.scala 83:35]
  reg [31:0] nonSaturatedMisses_1_query_instruction; // @[missHandler.scala 83:35]
  reg [3:0] nonSaturatedMisses_1_query_branchMask; // @[missHandler.scala 83:35]
  reg [3:0] nonSaturatedMisses_1_query_robAddr; // @[missHandler.scala 83:35]
  reg [5:0] nonSaturatedMisses_1_query_prfDest; // @[missHandler.scala 83:35]
  reg [63:0] nonSaturatedMisses_1_data; // @[missHandler.scala 83:35]
  reg  nonSaturatedMisses_2_query_valid; // @[missHandler.scala 83:35]
  reg [31:0] nonSaturatedMisses_2_query_address; // @[missHandler.scala 83:35]
  reg [31:0] nonSaturatedMisses_2_query_instruction; // @[missHandler.scala 83:35]
  reg [3:0] nonSaturatedMisses_2_query_branchMask; // @[missHandler.scala 83:35]
  reg [3:0] nonSaturatedMisses_2_query_robAddr; // @[missHandler.scala 83:35]
  reg [5:0] nonSaturatedMisses_2_query_prfDest; // @[missHandler.scala 83:35]
  reg [63:0] nonSaturatedMisses_2_data; // @[missHandler.scala 83:35]
  reg  nonSaturatedMisses_3_query_valid; // @[missHandler.scala 83:35]
  reg [31:0] nonSaturatedMisses_3_query_address; // @[missHandler.scala 83:35]
  reg [31:0] nonSaturatedMisses_3_query_instruction; // @[missHandler.scala 83:35]
  reg [3:0] nonSaturatedMisses_3_query_branchMask; // @[missHandler.scala 83:35]
  reg [3:0] nonSaturatedMisses_3_query_robAddr; // @[missHandler.scala 83:35]
  reg [5:0] nonSaturatedMisses_3_query_prfDest; // @[missHandler.scala 83:35]
  reg [63:0] nonSaturatedMisses_3_data; // @[missHandler.scala 83:35]
  reg [1:0] handlerStatus; // @[missHandler.scala 86:30]
  reg  saturated; // @[missHandler.scala 88:32]
  wire  _replayingQuries_T_3 = saturatedReplayVector_0_query_valid | saturatedReplayVector_1_query_valid |
    saturatedReplayVector_2_query_valid | saturatedReplayVector_3_query_valid | saturatedReplayVector_4_query_valid; // @[missHandler.scala 91:72]
  wire  _replayingQuries_T_4 = handlerStatus == 2'h3; // @[missHandler.scala 91:96]
  wire  _replayingQuries_T_6 = handlerStatus == 2'h2; // @[missHandler.scala 91:129]
  wire  _replayOut_T_1_query_valid = _replayingQuries_T_4 ? nonSaturatedMisses_0_query_valid :
    saturatedReplayVector_0_query_valid; // @[missHandler.scala 93:19]
  wire [3:0] _T_1 = branchOps_branchMask & saturatedReplayVector_1_query_branchMask; // @[missHandler.scala 107:52]
  wire  _T_2 = |_T_1; // @[missHandler.scala 107:77]
  wire [3:0] _saturatedReplayVector_0_query_branchMask_T = branchOps_branchMask ^
    saturatedReplayVector_1_query_branchMask; // @[missHandler.scala 107:128]
  wire  _T_3 = ~branchOps_passed; // @[missHandler.scala 108:30]
  wire [3:0] _T_7 = branchOps_branchMask & saturatedReplayVector_2_query_branchMask; // @[missHandler.scala 107:52]
  wire  _T_8 = |_T_7; // @[missHandler.scala 107:77]
  wire [3:0] _saturatedReplayVector_1_query_branchMask_T = branchOps_branchMask ^
    saturatedReplayVector_2_query_branchMask; // @[missHandler.scala 107:128]
  wire [3:0] _T_13 = branchOps_branchMask & saturatedReplayVector_3_query_branchMask; // @[missHandler.scala 107:52]
  wire  _T_14 = |_T_13; // @[missHandler.scala 107:77]
  wire [3:0] _saturatedReplayVector_2_query_branchMask_T = branchOps_branchMask ^
    saturatedReplayVector_3_query_branchMask; // @[missHandler.scala 107:128]
  wire [3:0] _T_19 = branchOps_branchMask & saturatedReplayVector_4_query_branchMask; // @[missHandler.scala 107:52]
  wire  _T_20 = |_T_19; // @[missHandler.scala 107:77]
  wire [3:0] _saturatedReplayVector_3_query_branchMask_T = branchOps_branchMask ^
    saturatedReplayVector_4_query_branchMask; // @[missHandler.scala 107:128]
  wire  _T_28 = nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid | nonSaturatedMisses_2_query_valid
     | nonSaturatedMisses_3_query_valid; // @[missHandler.scala 115:95]
  wire  _T_29 = ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid | nonSaturatedMisses_2_query_valid
     | nonSaturatedMisses_3_query_valid); // @[missHandler.scala 115:47]
  wire  _T_31 = _replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
    nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty; // @[missHandler.scala 115:101]
  wire [3:0] _T_32 = branchOps_branchMask & saturatedCollectVector_0_query_branchMask; // @[missHandler.scala 121:60]
  wire  _T_33 = |_T_32; // @[missHandler.scala 121:85]
  wire [3:0] _saturatedReplayVector_0_query_branchMask_T_1 = branchOps_branchMask ^
    saturatedCollectVector_0_query_branchMask; // @[missHandler.scala 121:136]
  wire [3:0] _T_38 = branchOps_branchMask & saturatedCollectVector_1_query_branchMask; // @[missHandler.scala 121:60]
  wire  _T_39 = |_T_38; // @[missHandler.scala 121:85]
  wire [3:0] _saturatedReplayVector_1_query_branchMask_T_1 = branchOps_branchMask ^
    saturatedCollectVector_1_query_branchMask; // @[missHandler.scala 121:136]
  wire [3:0] _T_44 = branchOps_branchMask & saturatedCollectVector_2_query_branchMask; // @[missHandler.scala 121:60]
  wire  _T_45 = |_T_44; // @[missHandler.scala 121:85]
  wire [3:0] _saturatedReplayVector_2_query_branchMask_T_1 = branchOps_branchMask ^
    saturatedCollectVector_2_query_branchMask; // @[missHandler.scala 121:136]
  wire [3:0] _T_50 = branchOps_branchMask & saturatedCollectVector_3_query_branchMask; // @[missHandler.scala 121:60]
  wire  _T_51 = |_T_50; // @[missHandler.scala 121:85]
  wire [3:0] _saturatedReplayVector_3_query_branchMask_T_1 = branchOps_branchMask ^
    saturatedCollectVector_3_query_branchMask; // @[missHandler.scala 121:136]
  wire [3:0] _T_56 = branchOps_branchMask & saturatedCollectVector_4_query_branchMask; // @[missHandler.scala 121:60]
  wire  _T_57 = |_T_56; // @[missHandler.scala 121:85]
  wire [3:0] _saturatedReplayVector_4_query_branchMask_T = branchOps_branchMask ^
    saturatedCollectVector_4_query_branchMask; // @[missHandler.scala 121:136]
  wire  _GEN_34 = _T_3 & _T_57 ? 1'h0 : saturatedCollectVector_4_query_valid; // @[missHandler.scala 122:{111,129} 119:29]
  wire  _GEN_36 = branchOps_valid ? _GEN_34 : saturatedCollectVector_4_query_valid; // @[missHandler.scala 119:29 120:48]
  wire  _GEN_65 = _replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
    nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty & _GEN_36; // @[missHandler.scala 115:124 112:75]
  reg [31:0] servicingBlock; // @[missHandler.scala 127:33]
  wire  _T_62 = ~saturated; // @[missHandler.scala 131:14]
  wire  _T_63 = handlerStatus != 2'h0; // @[missHandler.scala 134:39]
  wire  _T_64 = handlerStatus != 2'h0 & missedRequest_query_valid; // @[missHandler.scala 134:48]
  wire  _T_68 = nonSaturatedMisses_0_query_valid & nonSaturatedMisses_1_query_valid; // @[missHandler.scala 136:163]
  wire  _T_69 = nonSaturatedMisses_0_query_valid & nonSaturatedMisses_1_query_valid & nonSaturatedMisses_2_query_valid; // @[missHandler.scala 136:163]
  wire  _T_71 = missedRequest_query_address[31:6] != servicingBlock[31:6] | nonSaturatedMisses_0_query_valid &
    nonSaturatedMisses_1_query_valid & nonSaturatedMisses_2_query_valid & nonSaturatedMisses_3_query_valid; // @[missHandler.scala 136:113]
  wire  _T_72 = _T_64 & _T_71; // @[missHandler.scala 135:51]
  wire [3:0] _T_73 = missedRequest_query_branchMask & branchOps_branchMask; // @[missHandler.scala 141:70]
  wire  _T_74 = |_T_73; // @[missHandler.scala 141:94]
  wire [3:0] _saturatedCollectVector_0_query_branchMask_T = missedRequest_query_branchMask ^ branchOps_branchMask; // @[missHandler.scala 141:177]
  wire [3:0] _GEN_72 = |_T_73 ? _saturatedCollectVector_0_query_branchMask_T : missedRequest_query_branchMask; // @[missHandler.scala 141:143 138:51 141:99]
  wire  _GEN_73 = _T_3 & _T_74 ? 1'h0 : missedRequest_query_valid; // @[missHandler.scala 142:{120,160} 138:51]
  wire [3:0] _GEN_74 = branchOps_valid ? _GEN_72 : missedRequest_query_branchMask; // @[missHandler.scala 140:47 138:51]
  wire  _GEN_75 = branchOps_valid ? _GEN_73 : missedRequest_query_valid; // @[missHandler.scala 140:47 138:51]
  wire  _GEN_83 = _T_72 | saturated; // @[missHandler.scala 137:19 139:35 88:32]
  wire [3:0] _T_79 = saturatedCollectVector_0_query_branchMask & branchOps_branchMask; // @[missHandler.scala 150:61]
  wire  _T_80 = |_T_79; // @[missHandler.scala 150:85]
  wire [3:0] _saturatedCollectVectorUpdate_0_query_branchMask_T = saturatedCollectVector_0_query_branchMask ^
    branchOps_branchMask; // @[missHandler.scala 150:140]
  wire  _GEN_85 = _T_3 & _T_80 ? 1'h0 : saturatedCollectVector_0_query_valid; // @[missHandler.scala 151:{111,132} 148:32]
  wire  saturatedCollectVectorUpdate_0_query_valid = branchOps_valid ? _GEN_85 : saturatedCollectVector_0_query_valid; // @[missHandler.scala 148:32 149:47]
  wire [3:0] _T_85 = saturatedCollectVector_1_query_branchMask & branchOps_branchMask; // @[missHandler.scala 150:61]
  wire  _T_86 = |_T_85; // @[missHandler.scala 150:85]
  wire [3:0] _saturatedCollectVectorUpdate_1_query_branchMask_T = saturatedCollectVector_1_query_branchMask ^
    branchOps_branchMask; // @[missHandler.scala 150:140]
  wire  _GEN_89 = _T_3 & _T_86 ? 1'h0 : saturatedCollectVector_1_query_valid; // @[missHandler.scala 151:{111,132} 148:32]
  wire  saturatedCollectVectorUpdate_1_query_valid = branchOps_valid ? _GEN_89 : saturatedCollectVector_1_query_valid; // @[missHandler.scala 148:32 149:47]
  wire [3:0] _T_91 = saturatedCollectVector_2_query_branchMask & branchOps_branchMask; // @[missHandler.scala 150:61]
  wire  _T_92 = |_T_91; // @[missHandler.scala 150:85]
  wire [3:0] _saturatedCollectVectorUpdate_2_query_branchMask_T = saturatedCollectVector_2_query_branchMask ^
    branchOps_branchMask; // @[missHandler.scala 150:140]
  wire  _GEN_93 = _T_3 & _T_92 ? 1'h0 : saturatedCollectVector_2_query_valid; // @[missHandler.scala 151:{111,132} 148:32]
  wire  saturatedCollectVectorUpdate_2_query_valid = branchOps_valid ? _GEN_93 : saturatedCollectVector_2_query_valid; // @[missHandler.scala 148:32 149:47]
  wire [3:0] _T_97 = saturatedCollectVector_3_query_branchMask & branchOps_branchMask; // @[missHandler.scala 150:61]
  wire  _T_98 = |_T_97; // @[missHandler.scala 150:85]
  wire [3:0] _saturatedCollectVectorUpdate_3_query_branchMask_T = saturatedCollectVector_3_query_branchMask ^
    branchOps_branchMask; // @[missHandler.scala 150:140]
  wire  _GEN_97 = _T_3 & _T_98 ? 1'h0 : saturatedCollectVector_3_query_valid; // @[missHandler.scala 151:{111,132} 148:32]
  wire  saturatedCollectVectorUpdate_3_query_valid = branchOps_valid ? _GEN_97 : saturatedCollectVector_3_query_valid; // @[missHandler.scala 148:32 149:47]
  wire [3:0] _T_103 = saturatedCollectVector_4_query_branchMask & branchOps_branchMask; // @[missHandler.scala 150:61]
  wire  _T_104 = |_T_103; // @[missHandler.scala 150:85]
  wire [3:0] _saturatedCollectVectorUpdate_4_query_branchMask_T = saturatedCollectVector_4_query_branchMask ^
    branchOps_branchMask; // @[missHandler.scala 150:140]
  wire  _GEN_101 = _T_3 & _T_104 ? 1'h0 : saturatedCollectVector_4_query_valid; // @[missHandler.scala 151:{111,132} 148:32]
  wire  saturatedCollectVectorUpdate_4_query_valid = branchOps_valid ? _GEN_101 : saturatedCollectVector_4_query_valid; // @[missHandler.scala 148:32 149:47]
  wire  _T_116 = saturatedCollectVector_0_query_valid & saturatedCollectVector_1_query_valid; // @[missHandler.scala 156:79]
  wire  _T_117 = saturatedCollectVector_0_query_valid & saturatedCollectVector_1_query_valid &
    saturatedCollectVector_2_query_valid; // @[missHandler.scala 156:79]
  wire  _T_118 = saturatedCollectVector_0_query_valid & saturatedCollectVector_1_query_valid &
    saturatedCollectVector_2_query_valid & saturatedCollectVector_3_query_valid; // @[missHandler.scala 156:79]
  reg [63:0] cacheWrite_data; // @[missHandler.scala 166:33]
  reg  cacheWrite_valid; // @[missHandler.scala 166:33]
  reg [8:0] cacheWrite_address; // @[missHandler.scala 166:33]
  reg [1:0] cacheWrite_setSelVector; // @[missHandler.scala 166:33]
  reg [31:0] fetched_0_rdata; // @[missHandler.scala 173:30]
  reg  fetched_0_valid; // @[missHandler.scala 173:30]
  reg [31:0] fetched_1_rdata; // @[missHandler.scala 173:30]
  reg  fetched_1_valid; // @[missHandler.scala 173:30]
  wire  _T_143 = pushToCache_fired | ~cacheWrite_valid; // @[missHandler.scala 185:32]
  wire [63:0] _cacheWrite_data_T = {fetched_1_rdata,fetched_0_rdata}; // @[Cat.scala 33:92]
  wire  _cacheWrite_valid_T = fetched_0_valid & fetched_1_valid; // @[missHandler.scala 187:67]
  wire  _T_144 = 2'h0 == handlerStatus; // @[missHandler.scala 190:31]
  wire [9:0] _cacheWrite_address_T_1 = {missedRequest_query_address[12:6],3'h0}; // @[Cat.scala 33:92]
  wire [9:0] _GEN_187 = missedRequest_query_valid ? _cacheWrite_address_T_1 : {{1'd0}, cacheWrite_address}; // @[missHandler.scala 166:33 192:57 193:52]
  wire  _T_145 = 2'h1 == handlerStatus; // @[missHandler.scala 190:31]
  wire [8:0] _cacheWrite_address_T_3 = cacheWrite_address + 9'h1; // @[missHandler.scala 198:74]
  wire [8:0] _GEN_188 = pushToCache_fired ? _cacheWrite_address_T_3 : cacheWrite_address; // @[missHandler.scala 166:33 197:49 198:52]
  wire [8:0] _GEN_189 = 2'h1 == handlerStatus ? _GEN_188 : cacheWrite_address; // @[missHandler.scala 190:31 166:33]
  wire [9:0] _GEN_190 = 2'h0 == handlerStatus ? _GEN_187 : {{1'd0}, _GEN_189}; // @[missHandler.scala 190:31]
  wire  _T_150 = _T_143 & _cacheWrite_valid_T; // @[missHandler.scala 206:63]
  wire  _GEN_192 = ~fetched_0_valid | fetched_0_valid; // @[missHandler.scala 173:30 210:46 212:42]
  wire  _GEN_197 = _T_143 & _cacheWrite_valid_T | _GEN_192; // @[missHandler.scala 206:103 209:42]
  reg  clearToFetch; // @[missHandler.scala 224:35]
  wire  _dependencyCheck_requset_valid_T = handlerStatus == 2'h1; // @[missHandler.scala 234:57]
  reg  requested; // @[missHandler.scala 237:32]
  wire  _T_156 = ~requested; // @[missHandler.scala 239:14]
  wire  _requested_T = axi_ARVALID & axi_ARREADY; // @[missHandler.scala 239:53]
  reg  arvalid; // @[missHandler.scala 246:38]
  reg  rready; // @[missHandler.scala 246:38]
  wire  _GEN_215 = _T_144 ? _GEN_75 : nonSaturatedMisses_0_query_valid; // @[missHandler.scala 256:31 83:35]
  wire [31:0] _GEN_216 = _T_144 ? missedRequest_query_address : nonSaturatedMisses_0_query_address; // @[missHandler.scala 256:31 258:47 83:35]
  wire [31:0] _GEN_217 = _T_144 ? missedRequest_query_instruction : nonSaturatedMisses_0_query_instruction; // @[missHandler.scala 256:31 258:47 83:35]
  wire [3:0] _GEN_218 = _T_144 ? _GEN_74 : nonSaturatedMisses_0_query_branchMask; // @[missHandler.scala 256:31 83:35]
  wire [3:0] _GEN_219 = _T_144 ? missedRequest_query_robAddr : nonSaturatedMisses_0_query_robAddr; // @[missHandler.scala 256:31 258:47 83:35]
  wire [5:0] _GEN_220 = _T_144 ? missedRequest_query_prfDest : nonSaturatedMisses_0_query_prfDest; // @[missHandler.scala 256:31 258:47 83:35]
  wire [63:0] _GEN_221 = _T_144 ? missedRequest_data : nonSaturatedMisses_0_data; // @[missHandler.scala 256:31 258:47 83:35]
  wire [3:0] _T_170 = nonSaturatedMisses_0_query_branchMask & branchOps_branchMask; // @[missHandler.scala 287:61]
  wire  _T_171 = |_T_170; // @[missHandler.scala 287:85]
  wire [3:0] _nonSaturatedMissesUpdate_0_query_branchMask_T = nonSaturatedMisses_0_query_branchMask ^
    branchOps_branchMask; // @[missHandler.scala 287:140]
  wire [3:0] _GEN_222 = |_T_170 ? _nonSaturatedMissesUpdate_0_query_branchMask_T : nonSaturatedMisses_0_query_branchMask
    ; // @[missHandler.scala 287:115 285:32 287:90]
  wire  _GEN_223 = _T_3 & _T_171 ? 1'h0 : nonSaturatedMisses_0_query_valid; // @[missHandler.scala 288:{111,132} 285:32]
  wire [3:0] nonSaturatedMissesUpdate_0_query_branchMask = branchOps_valid ? _GEN_222 :
    nonSaturatedMisses_0_query_branchMask; // @[missHandler.scala 285:32 286:47]
  wire  nonSaturatedMissesUpdate_0_query_valid = branchOps_valid ? _GEN_223 : nonSaturatedMisses_0_query_valid; // @[missHandler.scala 285:32 286:47]
  wire [3:0] _T_176 = nonSaturatedMisses_1_query_branchMask & branchOps_branchMask; // @[missHandler.scala 287:61]
  wire  _T_177 = |_T_176; // @[missHandler.scala 287:85]
  wire [3:0] _nonSaturatedMissesUpdate_1_query_branchMask_T = nonSaturatedMisses_1_query_branchMask ^
    branchOps_branchMask; // @[missHandler.scala 287:140]
  wire [3:0] _GEN_226 = |_T_176 ? _nonSaturatedMissesUpdate_1_query_branchMask_T : nonSaturatedMisses_1_query_branchMask
    ; // @[missHandler.scala 287:115 285:32 287:90]
  wire  _GEN_227 = _T_3 & _T_177 ? 1'h0 : nonSaturatedMisses_1_query_valid; // @[missHandler.scala 288:{111,132} 285:32]
  wire [3:0] nonSaturatedMissesUpdate_1_query_branchMask = branchOps_valid ? _GEN_226 :
    nonSaturatedMisses_1_query_branchMask; // @[missHandler.scala 285:32 286:47]
  wire  nonSaturatedMissesUpdate_1_query_valid = branchOps_valid ? _GEN_227 : nonSaturatedMisses_1_query_valid; // @[missHandler.scala 285:32 286:47]
  wire [3:0] _T_182 = nonSaturatedMisses_2_query_branchMask & branchOps_branchMask; // @[missHandler.scala 287:61]
  wire  _T_183 = |_T_182; // @[missHandler.scala 287:85]
  wire [3:0] _nonSaturatedMissesUpdate_2_query_branchMask_T = nonSaturatedMisses_2_query_branchMask ^
    branchOps_branchMask; // @[missHandler.scala 287:140]
  wire [3:0] _GEN_230 = |_T_182 ? _nonSaturatedMissesUpdate_2_query_branchMask_T : nonSaturatedMisses_2_query_branchMask
    ; // @[missHandler.scala 287:115 285:32 287:90]
  wire  _GEN_231 = _T_3 & _T_183 ? 1'h0 : nonSaturatedMisses_2_query_valid; // @[missHandler.scala 288:{111,132} 285:32]
  wire [3:0] nonSaturatedMissesUpdate_2_query_branchMask = branchOps_valid ? _GEN_230 :
    nonSaturatedMisses_2_query_branchMask; // @[missHandler.scala 285:32 286:47]
  wire  nonSaturatedMissesUpdate_2_query_valid = branchOps_valid ? _GEN_231 : nonSaturatedMisses_2_query_valid; // @[missHandler.scala 285:32 286:47]
  wire [3:0] _T_188 = nonSaturatedMisses_3_query_branchMask & branchOps_branchMask; // @[missHandler.scala 287:61]
  wire  _T_189 = |_T_188; // @[missHandler.scala 287:85]
  wire [3:0] _nonSaturatedMissesUpdate_3_query_branchMask_T = nonSaturatedMisses_3_query_branchMask ^
    branchOps_branchMask; // @[missHandler.scala 287:140]
  wire [3:0] _GEN_234 = |_T_188 ? _nonSaturatedMissesUpdate_3_query_branchMask_T : nonSaturatedMisses_3_query_branchMask
    ; // @[missHandler.scala 287:115 285:32 287:90]
  wire  _GEN_235 = _T_3 & _T_189 ? 1'h0 : nonSaturatedMisses_3_query_valid; // @[missHandler.scala 288:{111,132} 285:32]
  wire [3:0] nonSaturatedMissesUpdate_3_query_branchMask = branchOps_valid ? _GEN_234 :
    nonSaturatedMisses_3_query_branchMask; // @[missHandler.scala 285:32 286:47]
  wire  nonSaturatedMissesUpdate_3_query_valid = branchOps_valid ? _GEN_235 : nonSaturatedMisses_3_query_valid; // @[missHandler.scala 285:32 286:47]
  wire  nonSaturatedMissesUpdate_4_query_valid = missedRequest_query_valid & _T_62 & ~_T_71; // @[missHandler.scala 291:132]
  wire  _GEN_242 = ~nonSaturatedMisses_0_query_valid ? nonSaturatedMissesUpdate_1_query_valid :
    nonSaturatedMissesUpdate_0_query_valid; // @[missHandler.scala 297:{119,125,151}]
  wire [31:0] _GEN_243 = ~nonSaturatedMisses_0_query_valid ? nonSaturatedMisses_1_query_address :
    nonSaturatedMisses_0_query_address; // @[missHandler.scala 297:{119,125,151}]
  wire [31:0] _GEN_244 = ~nonSaturatedMisses_0_query_valid ? nonSaturatedMisses_1_query_instruction :
    nonSaturatedMisses_0_query_instruction; // @[missHandler.scala 297:{119,125,151}]
  wire [3:0] _GEN_245 = ~nonSaturatedMisses_0_query_valid ? nonSaturatedMissesUpdate_1_query_branchMask :
    nonSaturatedMissesUpdate_0_query_branchMask; // @[missHandler.scala 297:{119,125,151}]
  wire [3:0] _GEN_246 = ~nonSaturatedMisses_0_query_valid ? nonSaturatedMisses_1_query_robAddr :
    nonSaturatedMisses_0_query_robAddr; // @[missHandler.scala 297:{119,125,151}]
  wire [5:0] _GEN_247 = ~nonSaturatedMisses_0_query_valid ? nonSaturatedMisses_1_query_prfDest :
    nonSaturatedMisses_0_query_prfDest; // @[missHandler.scala 297:{119,125,151}]
  wire [63:0] _GEN_248 = ~nonSaturatedMisses_0_query_valid ? nonSaturatedMisses_1_data : nonSaturatedMisses_0_data; // @[missHandler.scala 297:{119,125,151}]
  wire  _GEN_249 = ~nonSaturatedMisses_0_query_valid | ~nonSaturatedMisses_1_query_valid ?
    nonSaturatedMissesUpdate_2_query_valid : nonSaturatedMissesUpdate_1_query_valid; // @[missHandler.scala 297:{119,125,151}]
  wire [31:0] _GEN_250 = ~nonSaturatedMisses_0_query_valid | ~nonSaturatedMisses_1_query_valid ?
    nonSaturatedMisses_2_query_address : nonSaturatedMisses_1_query_address; // @[missHandler.scala 297:{119,125,151}]
  wire [31:0] _GEN_251 = ~nonSaturatedMisses_0_query_valid | ~nonSaturatedMisses_1_query_valid ?
    nonSaturatedMisses_2_query_instruction : nonSaturatedMisses_1_query_instruction; // @[missHandler.scala 297:{119,125,151}]
  wire [3:0] _GEN_252 = ~nonSaturatedMisses_0_query_valid | ~nonSaturatedMisses_1_query_valid ?
    nonSaturatedMissesUpdate_2_query_branchMask : nonSaturatedMissesUpdate_1_query_branchMask; // @[missHandler.scala 297:{119,125,151}]
  wire [3:0] _GEN_253 = ~nonSaturatedMisses_0_query_valid | ~nonSaturatedMisses_1_query_valid ?
    nonSaturatedMisses_2_query_robAddr : nonSaturatedMisses_1_query_robAddr; // @[missHandler.scala 297:{119,125,151}]
  wire [5:0] _GEN_254 = ~nonSaturatedMisses_0_query_valid | ~nonSaturatedMisses_1_query_valid ?
    nonSaturatedMisses_2_query_prfDest : nonSaturatedMisses_1_query_prfDest; // @[missHandler.scala 297:{119,125,151}]
  wire [63:0] _GEN_255 = ~nonSaturatedMisses_0_query_valid | ~nonSaturatedMisses_1_query_valid ?
    nonSaturatedMisses_2_data : nonSaturatedMisses_1_data; // @[missHandler.scala 297:{119,125,151}]
  wire  _GEN_256 = ~_T_68 | ~nonSaturatedMisses_2_query_valid ? nonSaturatedMissesUpdate_3_query_valid :
    nonSaturatedMissesUpdate_2_query_valid; // @[missHandler.scala 297:{119,125,151}]
  wire [31:0] _GEN_257 = ~_T_68 | ~nonSaturatedMisses_2_query_valid ? nonSaturatedMisses_3_query_address :
    nonSaturatedMisses_2_query_address; // @[missHandler.scala 297:{119,125,151}]
  wire [31:0] _GEN_258 = ~_T_68 | ~nonSaturatedMisses_2_query_valid ? nonSaturatedMisses_3_query_instruction :
    nonSaturatedMisses_2_query_instruction; // @[missHandler.scala 297:{119,125,151}]
  wire [3:0] _GEN_259 = ~_T_68 | ~nonSaturatedMisses_2_query_valid ? nonSaturatedMissesUpdate_3_query_branchMask :
    nonSaturatedMissesUpdate_2_query_branchMask; // @[missHandler.scala 297:{119,125,151}]
  wire [3:0] _GEN_260 = ~_T_68 | ~nonSaturatedMisses_2_query_valid ? nonSaturatedMisses_3_query_robAddr :
    nonSaturatedMisses_2_query_robAddr; // @[missHandler.scala 297:{119,125,151}]
  wire [5:0] _GEN_261 = ~_T_68 | ~nonSaturatedMisses_2_query_valid ? nonSaturatedMisses_3_query_prfDest :
    nonSaturatedMisses_2_query_prfDest; // @[missHandler.scala 297:{119,125,151}]
  wire [63:0] _GEN_262 = ~_T_68 | ~nonSaturatedMisses_2_query_valid ? nonSaturatedMisses_3_data :
    nonSaturatedMisses_2_data; // @[missHandler.scala 297:{119,125,151}]
  wire  _GEN_263 = ~_T_69 | ~nonSaturatedMisses_3_query_valid ? nonSaturatedMissesUpdate_4_query_valid :
    nonSaturatedMissesUpdate_3_query_valid; // @[missHandler.scala 297:{119,125,151}]
  wire  _GEN_270 = _T_63 ? _GEN_242 : _GEN_215; // @[missHandler.scala 282:38]
  wire [31:0] _GEN_271 = _T_63 ? _GEN_243 : _GEN_216; // @[missHandler.scala 282:38]
  wire [31:0] _GEN_272 = _T_63 ? _GEN_244 : _GEN_217; // @[missHandler.scala 282:38]
  wire [3:0] _GEN_273 = _T_63 ? _GEN_245 : _GEN_218; // @[missHandler.scala 282:38]
  wire [3:0] _GEN_274 = _T_63 ? _GEN_246 : _GEN_219; // @[missHandler.scala 282:38]
  wire [5:0] _GEN_275 = _T_63 ? _GEN_247 : _GEN_220; // @[missHandler.scala 282:38]
  wire [63:0] _GEN_276 = _T_63 ? _GEN_248 : _GEN_221; // @[missHandler.scala 282:38]
  wire  _GEN_277 = _T_63 ? _GEN_249 : nonSaturatedMisses_1_query_valid; // @[missHandler.scala 282:38 83:35]
  wire [31:0] _GEN_278 = _T_63 ? _GEN_250 : nonSaturatedMisses_1_query_address; // @[missHandler.scala 282:38 83:35]
  wire [31:0] _GEN_279 = _T_63 ? _GEN_251 : nonSaturatedMisses_1_query_instruction; // @[missHandler.scala 282:38 83:35]
  wire [3:0] _GEN_280 = _T_63 ? _GEN_252 : nonSaturatedMisses_1_query_branchMask; // @[missHandler.scala 282:38 83:35]
  wire [3:0] _GEN_281 = _T_63 ? _GEN_253 : nonSaturatedMisses_1_query_robAddr; // @[missHandler.scala 282:38 83:35]
  wire [5:0] _GEN_282 = _T_63 ? _GEN_254 : nonSaturatedMisses_1_query_prfDest; // @[missHandler.scala 282:38 83:35]
  wire [63:0] _GEN_283 = _T_63 ? _GEN_255 : nonSaturatedMisses_1_data; // @[missHandler.scala 282:38 83:35]
  wire  _GEN_284 = _T_63 ? _GEN_256 : nonSaturatedMisses_2_query_valid; // @[missHandler.scala 282:38 83:35]
  wire [31:0] _GEN_285 = _T_63 ? _GEN_257 : nonSaturatedMisses_2_query_address; // @[missHandler.scala 282:38 83:35]
  wire [31:0] _GEN_286 = _T_63 ? _GEN_258 : nonSaturatedMisses_2_query_instruction; // @[missHandler.scala 282:38 83:35]
  wire [3:0] _GEN_287 = _T_63 ? _GEN_259 : nonSaturatedMisses_2_query_branchMask; // @[missHandler.scala 282:38 83:35]
  wire [3:0] _GEN_288 = _T_63 ? _GEN_260 : nonSaturatedMisses_2_query_robAddr; // @[missHandler.scala 282:38 83:35]
  wire [5:0] _GEN_289 = _T_63 ? _GEN_261 : nonSaturatedMisses_2_query_prfDest; // @[missHandler.scala 282:38 83:35]
  wire [63:0] _GEN_290 = _T_63 ? _GEN_262 : nonSaturatedMisses_2_data; // @[missHandler.scala 282:38 83:35]
  wire  _GEN_291 = _T_63 ? _GEN_263 : nonSaturatedMisses_3_query_valid; // @[missHandler.scala 282:38 83:35]
  reg [1:0] nextSet; // @[missHandler.scala 300:26]
  reg [1:0] randSelect; // @[missHandler.scala 304:33]
  wire  _rlastToCache_T_1 = &cacheWrite_address[2:0]; // @[missHandler.scala 309:62]
  wire  _setInvalidateVector_T = &setFillStatus; // @[missHandler.scala 317:31]
  wire  _setInvalidateVector_T_3 = ~setFillStatus[0]; // @[missHandler.scala 319:84]
  wire  _setInvalidateVector_T_6 = ~setFillStatus[1]; // @[missHandler.scala 319:84]
  wire [1:0] _setInvalidateVector_T_7 = _setInvalidateVector_T_6 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _setInvalidateVector_T_8 = _setInvalidateVector_T_3 ? 2'h1 : _setInvalidateVector_T_7; // @[Mux.scala 101:16]
  wire [31:0] _servicingBlock_T_1 = {missedRequest_query_address[31:6],6'h0}; // @[Cat.scala 33:92]
  wire [1:0] _GEN_303 = cachePipelineEmpty ? 2'h3 : handlerStatus; // @[missHandler.scala 351:{51,67} 86:30]
  wire [1:0] _GEN_304 = _T_29 & cachePipelineEmpty ? 2'h0 : handlerStatus; // @[missHandler.scala 354:108 355:47 86:30]
  wire [1:0] _GEN_305 = 2'h3 == handlerStatus ? _GEN_304 : handlerStatus; // @[missHandler.scala 340:31 86:30]
  wire  _GEN_306 = 2'h3 == handlerStatus ? nonSaturatedMisses_1_query_valid : _GEN_270; // @[missHandler.scala 340:31 358:107]
  wire  _GEN_313 = 2'h3 == handlerStatus ? nonSaturatedMisses_2_query_valid : _GEN_277; // @[missHandler.scala 340:31 358:107]
  wire  _GEN_320 = 2'h3 == handlerStatus ? nonSaturatedMisses_3_query_valid : _GEN_284; // @[missHandler.scala 340:31 358:107]
  wire  _GEN_327 = 2'h3 == handlerStatus ? 1'h0 : _GEN_291; // @[missHandler.scala 340:31 359:85]
  assign replayOut_query_valid = _replayingQuries_T_6 ? 1'h0 : _replayOut_T_1_query_valid; // @[missHandler.scala 93:13 94:46 95:39]
  assign replayOut_query_address = _replayingQuries_T_4 ? nonSaturatedMisses_0_query_address :
    saturatedReplayVector_0_query_address; // @[missHandler.scala 93:19]
  assign replayOut_query_instruction = _replayingQuries_T_4 ? nonSaturatedMisses_0_query_instruction :
    saturatedReplayVector_0_query_instruction; // @[missHandler.scala 93:19]
  assign replayOut_query_branchMask = _replayingQuries_T_4 ? nonSaturatedMisses_0_query_branchMask :
    saturatedReplayVector_0_query_branchMask; // @[missHandler.scala 93:19]
  assign replayOut_query_robAddr = _replayingQuries_T_4 ? nonSaturatedMisses_0_query_robAddr :
    saturatedReplayVector_0_query_robAddr; // @[missHandler.scala 93:19]
  assign replayOut_query_prfDest = _replayingQuries_T_4 ? nonSaturatedMisses_0_query_prfDest :
    saturatedReplayVector_0_query_prfDest; // @[missHandler.scala 93:19]
  assign replayOut_data = _replayingQuries_T_4 ? nonSaturatedMisses_0_data : saturatedReplayVector_0_data; // @[missHandler.scala 93:19]
  assign replayingQuries = saturatedReplayVector_0_query_valid | saturatedReplayVector_1_query_valid |
    saturatedReplayVector_2_query_valid | saturatedReplayVector_3_query_valid | saturatedReplayVector_4_query_valid |
    handlerStatus == 2'h3 | handlerStatus == 2'h2; // @[missHandler.scala 91:111]
  assign pushToCache_ready = cacheWrite_valid & (cachePipelineEmpty | ~rlastToCache); // @[missHandler.scala 365:47]
  assign pushToCache_cacheWriteOut_data = cacheWrite_data; // @[missHandler.scala 182:35]
  assign pushToCache_cacheWriteOut_address = cacheWrite_address; // @[missHandler.scala 182:35]
  assign pushToCache_cacheWriteOut_setSelVector = cacheWrite_setSelVector; // @[missHandler.scala 182:35]
  assign axi_ARADDR = servicingBlock; // @[missHandler.scala 367:20]
  assign axi_ARVALID = arvalid; // @[missHandler.scala 376:15]
  assign axi_RREADY = rready & (~_cacheWrite_valid_T | pushToCache_fired); // @[missHandler.scala 378:24]
  assign dependencyCheck_requset_valid = handlerStatus == 2'h1; // @[missHandler.scala 234:57]
  assign dependencyCheck_requset_address = servicingBlock; // @[missHandler.scala 233:41]
  assign rlastToCache = &cacheWrite_address[2:0]; // @[missHandler.scala 309:62]
  assign setInvalidateVector = _setInvalidateVector_T ? randSelect : _setInvalidateVector_T_8; // @[missHandler.scala 316:35]
  assign handlerBusy = handlerStatus != 2'h0; // @[missHandler.scala 334:38]
  assign handlerSaturated = saturated; // @[missHandler.scala 337:26]
  assign clean = ~(_T_28 | (saturatedCollectVector_0_query_valid | saturatedCollectVector_1_query_valid |
    saturatedCollectVector_2_query_valid | saturatedCollectVector_3_query_valid | saturatedCollectVector_4_query_valid)
     | _replayingQuries_T_3); // @[missHandler.scala 399:18]
  assign nonSaturatedReplay = handlerStatus == 2'h3; // @[missHandler.scala 402:46]
  always @(posedge clock) begin
    if (reset) begin // @[missHandler.scala 75:38]
      saturatedReplayVector_0_query_valid <= 1'h0; // @[missHandler.scala 75:38]
    end else if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      if (branchOps_valid) begin // @[missHandler.scala 120:48]
        if (_T_3 & _T_33) begin // @[missHandler.scala 122:111]
          saturatedReplayVector_0_query_valid <= 1'h0; // @[missHandler.scala 122:129]
        end else begin
          saturatedReplayVector_0_query_valid <= saturatedCollectVector_0_query_valid; // @[missHandler.scala 119:29]
        end
      end else begin
        saturatedReplayVector_0_query_valid <= saturatedCollectVector_0_query_valid; // @[missHandler.scala 119:29]
      end
    end else if (branchOps_valid) begin // @[missHandler.scala 106:40]
      if (~branchOps_passed & _T_2) begin // @[missHandler.scala 108:103]
        saturatedReplayVector_0_query_valid <= 1'h0; // @[missHandler.scala 108:121]
      end else begin
        saturatedReplayVector_0_query_valid <= saturatedReplayVector_1_query_valid; // @[missHandler.scala 105:21]
      end
    end else begin
      saturatedReplayVector_0_query_valid <= saturatedReplayVector_1_query_valid; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_0_query_address <= saturatedCollectVector_0_query_address; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_0_query_address <= saturatedReplayVector_1_query_address; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_0_query_instruction <= saturatedCollectVector_0_query_instruction; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_0_query_instruction <= saturatedReplayVector_1_query_instruction; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      if (branchOps_valid) begin // @[missHandler.scala 120:48]
        if (|_T_32) begin // @[missHandler.scala 121:90]
          saturatedReplayVector_0_query_branchMask <= _saturatedReplayVector_0_query_branchMask_T_1; // @[missHandler.scala 121:112]
        end else begin
          saturatedReplayVector_0_query_branchMask <= saturatedCollectVector_0_query_branchMask; // @[missHandler.scala 119:29]
        end
      end else begin
        saturatedReplayVector_0_query_branchMask <= saturatedCollectVector_0_query_branchMask; // @[missHandler.scala 119:29]
      end
    end else if (branchOps_valid) begin // @[missHandler.scala 106:40]
      if (|_T_1) begin // @[missHandler.scala 107:82]
        saturatedReplayVector_0_query_branchMask <= _saturatedReplayVector_0_query_branchMask_T; // @[missHandler.scala 107:104]
      end else begin
        saturatedReplayVector_0_query_branchMask <= saturatedReplayVector_1_query_branchMask; // @[missHandler.scala 105:21]
      end
    end else begin
      saturatedReplayVector_0_query_branchMask <= saturatedReplayVector_1_query_branchMask; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_0_query_robAddr <= saturatedCollectVector_0_query_robAddr; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_0_query_robAddr <= saturatedReplayVector_1_query_robAddr; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_0_query_prfDest <= saturatedCollectVector_0_query_prfDest; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_0_query_prfDest <= saturatedReplayVector_1_query_prfDest; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_0_data <= saturatedCollectVector_0_data; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_0_data <= saturatedReplayVector_1_data; // @[missHandler.scala 105:21]
    end
    if (reset) begin // @[missHandler.scala 75:38]
      saturatedReplayVector_1_query_valid <= 1'h0; // @[missHandler.scala 75:38]
    end else if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      if (branchOps_valid) begin // @[missHandler.scala 120:48]
        if (_T_3 & _T_39) begin // @[missHandler.scala 122:111]
          saturatedReplayVector_1_query_valid <= 1'h0; // @[missHandler.scala 122:129]
        end else begin
          saturatedReplayVector_1_query_valid <= saturatedCollectVector_1_query_valid; // @[missHandler.scala 119:29]
        end
      end else begin
        saturatedReplayVector_1_query_valid <= saturatedCollectVector_1_query_valid; // @[missHandler.scala 119:29]
      end
    end else if (branchOps_valid) begin // @[missHandler.scala 106:40]
      if (~branchOps_passed & _T_8) begin // @[missHandler.scala 108:103]
        saturatedReplayVector_1_query_valid <= 1'h0; // @[missHandler.scala 108:121]
      end else begin
        saturatedReplayVector_1_query_valid <= saturatedReplayVector_2_query_valid; // @[missHandler.scala 105:21]
      end
    end else begin
      saturatedReplayVector_1_query_valid <= saturatedReplayVector_2_query_valid; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_1_query_address <= saturatedCollectVector_1_query_address; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_1_query_address <= saturatedReplayVector_2_query_address; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_1_query_instruction <= saturatedCollectVector_1_query_instruction; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_1_query_instruction <= saturatedReplayVector_2_query_instruction; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      if (branchOps_valid) begin // @[missHandler.scala 120:48]
        if (|_T_38) begin // @[missHandler.scala 121:90]
          saturatedReplayVector_1_query_branchMask <= _saturatedReplayVector_1_query_branchMask_T_1; // @[missHandler.scala 121:112]
        end else begin
          saturatedReplayVector_1_query_branchMask <= saturatedCollectVector_1_query_branchMask; // @[missHandler.scala 119:29]
        end
      end else begin
        saturatedReplayVector_1_query_branchMask <= saturatedCollectVector_1_query_branchMask; // @[missHandler.scala 119:29]
      end
    end else if (branchOps_valid) begin // @[missHandler.scala 106:40]
      if (|_T_7) begin // @[missHandler.scala 107:82]
        saturatedReplayVector_1_query_branchMask <= _saturatedReplayVector_1_query_branchMask_T; // @[missHandler.scala 107:104]
      end else begin
        saturatedReplayVector_1_query_branchMask <= saturatedReplayVector_2_query_branchMask; // @[missHandler.scala 105:21]
      end
    end else begin
      saturatedReplayVector_1_query_branchMask <= saturatedReplayVector_2_query_branchMask; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_1_query_robAddr <= saturatedCollectVector_1_query_robAddr; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_1_query_robAddr <= saturatedReplayVector_2_query_robAddr; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_1_query_prfDest <= saturatedCollectVector_1_query_prfDest; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_1_query_prfDest <= saturatedReplayVector_2_query_prfDest; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_1_data <= saturatedCollectVector_1_data; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_1_data <= saturatedReplayVector_2_data; // @[missHandler.scala 105:21]
    end
    if (reset) begin // @[missHandler.scala 75:38]
      saturatedReplayVector_2_query_valid <= 1'h0; // @[missHandler.scala 75:38]
    end else if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      if (branchOps_valid) begin // @[missHandler.scala 120:48]
        if (_T_3 & _T_45) begin // @[missHandler.scala 122:111]
          saturatedReplayVector_2_query_valid <= 1'h0; // @[missHandler.scala 122:129]
        end else begin
          saturatedReplayVector_2_query_valid <= saturatedCollectVector_2_query_valid; // @[missHandler.scala 119:29]
        end
      end else begin
        saturatedReplayVector_2_query_valid <= saturatedCollectVector_2_query_valid; // @[missHandler.scala 119:29]
      end
    end else if (branchOps_valid) begin // @[missHandler.scala 106:40]
      if (~branchOps_passed & _T_14) begin // @[missHandler.scala 108:103]
        saturatedReplayVector_2_query_valid <= 1'h0; // @[missHandler.scala 108:121]
      end else begin
        saturatedReplayVector_2_query_valid <= saturatedReplayVector_3_query_valid; // @[missHandler.scala 105:21]
      end
    end else begin
      saturatedReplayVector_2_query_valid <= saturatedReplayVector_3_query_valid; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_2_query_address <= saturatedCollectVector_2_query_address; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_2_query_address <= saturatedReplayVector_3_query_address; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_2_query_instruction <= saturatedCollectVector_2_query_instruction; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_2_query_instruction <= saturatedReplayVector_3_query_instruction; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      if (branchOps_valid) begin // @[missHandler.scala 120:48]
        if (|_T_44) begin // @[missHandler.scala 121:90]
          saturatedReplayVector_2_query_branchMask <= _saturatedReplayVector_2_query_branchMask_T_1; // @[missHandler.scala 121:112]
        end else begin
          saturatedReplayVector_2_query_branchMask <= saturatedCollectVector_2_query_branchMask; // @[missHandler.scala 119:29]
        end
      end else begin
        saturatedReplayVector_2_query_branchMask <= saturatedCollectVector_2_query_branchMask; // @[missHandler.scala 119:29]
      end
    end else if (branchOps_valid) begin // @[missHandler.scala 106:40]
      if (|_T_13) begin // @[missHandler.scala 107:82]
        saturatedReplayVector_2_query_branchMask <= _saturatedReplayVector_2_query_branchMask_T; // @[missHandler.scala 107:104]
      end else begin
        saturatedReplayVector_2_query_branchMask <= saturatedReplayVector_3_query_branchMask; // @[missHandler.scala 105:21]
      end
    end else begin
      saturatedReplayVector_2_query_branchMask <= saturatedReplayVector_3_query_branchMask; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_2_query_robAddr <= saturatedCollectVector_2_query_robAddr; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_2_query_robAddr <= saturatedReplayVector_3_query_robAddr; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_2_query_prfDest <= saturatedCollectVector_2_query_prfDest; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_2_query_prfDest <= saturatedReplayVector_3_query_prfDest; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_2_data <= saturatedCollectVector_2_data; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_2_data <= saturatedReplayVector_3_data; // @[missHandler.scala 105:21]
    end
    if (reset) begin // @[missHandler.scala 75:38]
      saturatedReplayVector_3_query_valid <= 1'h0; // @[missHandler.scala 75:38]
    end else if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      if (branchOps_valid) begin // @[missHandler.scala 120:48]
        if (_T_3 & _T_51) begin // @[missHandler.scala 122:111]
          saturatedReplayVector_3_query_valid <= 1'h0; // @[missHandler.scala 122:129]
        end else begin
          saturatedReplayVector_3_query_valid <= saturatedCollectVector_3_query_valid; // @[missHandler.scala 119:29]
        end
      end else begin
        saturatedReplayVector_3_query_valid <= saturatedCollectVector_3_query_valid; // @[missHandler.scala 119:29]
      end
    end else if (branchOps_valid) begin // @[missHandler.scala 106:40]
      if (~branchOps_passed & _T_20) begin // @[missHandler.scala 108:103]
        saturatedReplayVector_3_query_valid <= 1'h0; // @[missHandler.scala 108:121]
      end else begin
        saturatedReplayVector_3_query_valid <= saturatedReplayVector_4_query_valid; // @[missHandler.scala 105:21]
      end
    end else begin
      saturatedReplayVector_3_query_valid <= saturatedReplayVector_4_query_valid; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_3_query_address <= saturatedCollectVector_3_query_address; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_3_query_address <= saturatedReplayVector_4_query_address; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_3_query_instruction <= saturatedCollectVector_3_query_instruction; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_3_query_instruction <= saturatedReplayVector_4_query_instruction; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      if (branchOps_valid) begin // @[missHandler.scala 120:48]
        if (|_T_50) begin // @[missHandler.scala 121:90]
          saturatedReplayVector_3_query_branchMask <= _saturatedReplayVector_3_query_branchMask_T_1; // @[missHandler.scala 121:112]
        end else begin
          saturatedReplayVector_3_query_branchMask <= saturatedCollectVector_3_query_branchMask; // @[missHandler.scala 119:29]
        end
      end else begin
        saturatedReplayVector_3_query_branchMask <= saturatedCollectVector_3_query_branchMask; // @[missHandler.scala 119:29]
      end
    end else if (branchOps_valid) begin // @[missHandler.scala 106:40]
      if (|_T_19) begin // @[missHandler.scala 107:82]
        saturatedReplayVector_3_query_branchMask <= _saturatedReplayVector_3_query_branchMask_T; // @[missHandler.scala 107:104]
      end else begin
        saturatedReplayVector_3_query_branchMask <= saturatedReplayVector_4_query_branchMask; // @[missHandler.scala 105:21]
      end
    end else begin
      saturatedReplayVector_3_query_branchMask <= saturatedReplayVector_4_query_branchMask; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_3_query_robAddr <= saturatedCollectVector_3_query_robAddr; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_3_query_robAddr <= saturatedReplayVector_4_query_robAddr; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_3_query_prfDest <= saturatedCollectVector_3_query_prfDest; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_3_query_prfDest <= saturatedReplayVector_4_query_prfDest; // @[missHandler.scala 105:21]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_3_data <= saturatedCollectVector_3_data; // @[missHandler.scala 119:29]
    end else begin
      saturatedReplayVector_3_data <= saturatedReplayVector_4_data; // @[missHandler.scala 105:21]
    end
    if (reset) begin // @[missHandler.scala 75:38]
      saturatedReplayVector_4_query_valid <= 1'h0; // @[missHandler.scala 75:38]
    end else begin
      saturatedReplayVector_4_query_valid <= _GEN_65;
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_4_query_address <= saturatedCollectVector_4_query_address; // @[missHandler.scala 119:29]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_4_query_instruction <= saturatedCollectVector_4_query_instruction; // @[missHandler.scala 119:29]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      if (branchOps_valid) begin // @[missHandler.scala 120:48]
        if (|_T_56) begin // @[missHandler.scala 121:90]
          saturatedReplayVector_4_query_branchMask <= _saturatedReplayVector_4_query_branchMask_T; // @[missHandler.scala 121:112]
        end else begin
          saturatedReplayVector_4_query_branchMask <= saturatedCollectVector_4_query_branchMask; // @[missHandler.scala 119:29]
        end
      end else begin
        saturatedReplayVector_4_query_branchMask <= saturatedCollectVector_4_query_branchMask; // @[missHandler.scala 119:29]
      end
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_4_query_robAddr <= saturatedCollectVector_4_query_robAddr; // @[missHandler.scala 119:29]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_4_query_prfDest <= saturatedCollectVector_4_query_prfDest; // @[missHandler.scala 119:29]
    end
    if (_replayingQuries_T_4 & ~(nonSaturatedMisses_0_query_valid | nonSaturatedMisses_1_query_valid |
      nonSaturatedMisses_2_query_valid | nonSaturatedMisses_3_query_valid) & cachePipelineEmpty) begin // @[missHandler.scala 115:124]
      saturatedReplayVector_4_data <= saturatedCollectVector_4_data; // @[missHandler.scala 119:29]
    end
    if (reset) begin // @[missHandler.scala 81:39]
      saturatedCollectVector_0_query_valid <= 1'h0; // @[missHandler.scala 81:39]
    end else if (~saturated) begin // @[missHandler.scala 131:26]
      if (_T_72) begin // @[missHandler.scala 137:19]
        if (branchOps_valid) begin // @[missHandler.scala 140:47]
          saturatedCollectVector_0_query_valid <= _GEN_73;
        end else begin
          saturatedCollectVector_0_query_valid <= missedRequest_query_valid; // @[missHandler.scala 138:51]
        end
      end
    end else if (_T_31) begin // @[missHandler.scala 160:132]
      saturatedCollectVector_0_query_valid <= 1'h0; // @[missHandler.scala 161:70]
    end else if (~saturatedCollectVector_0_query_valid) begin // @[missHandler.scala 158:117]
      saturatedCollectVector_0_query_valid <= saturatedCollectVectorUpdate_1_query_valid; // @[missHandler.scala 158:123]
    end else begin
      saturatedCollectVector_0_query_valid <= saturatedCollectVectorUpdate_0_query_valid; // @[missHandler.scala 158:149]
    end
    if (~saturated) begin // @[missHandler.scala 131:26]
      if (_T_72) begin // @[missHandler.scala 137:19]
        saturatedCollectVector_0_query_address <= missedRequest_query_address; // @[missHandler.scala 138:51]
      end
    end else if (~saturatedCollectVector_0_query_valid) begin // @[missHandler.scala 158:117]
      saturatedCollectVector_0_query_address <= saturatedCollectVector_1_query_address; // @[missHandler.scala 158:123]
    end
    if (~saturated) begin // @[missHandler.scala 131:26]
      if (_T_72) begin // @[missHandler.scala 137:19]
        saturatedCollectVector_0_query_instruction <= missedRequest_query_instruction; // @[missHandler.scala 138:51]
      end
    end else if (~saturatedCollectVector_0_query_valid) begin // @[missHandler.scala 158:117]
      saturatedCollectVector_0_query_instruction <= saturatedCollectVector_1_query_instruction; // @[missHandler.scala 158:123]
    end
    if (~saturated) begin // @[missHandler.scala 131:26]
      if (_T_72) begin // @[missHandler.scala 137:19]
        if (branchOps_valid) begin // @[missHandler.scala 140:47]
          if (|_T_73) begin // @[missHandler.scala 141:99]
            saturatedCollectVector_0_query_branchMask <= _saturatedCollectVector_0_query_branchMask_T; // @[missHandler.scala 141:143]
          end else begin
            saturatedCollectVector_0_query_branchMask <= missedRequest_query_branchMask; // @[missHandler.scala 138:51]
          end
        end else begin
          saturatedCollectVector_0_query_branchMask <= missedRequest_query_branchMask; // @[missHandler.scala 138:51]
        end
      end
    end else if (~saturatedCollectVector_0_query_valid) begin // @[missHandler.scala 158:117]
      if (branchOps_valid) begin // @[missHandler.scala 149:47]
        if (|_T_85) begin // @[missHandler.scala 150:90]
          saturatedCollectVector_0_query_branchMask <= _saturatedCollectVectorUpdate_1_query_branchMask_T; // @[missHandler.scala 150:115]
        end else begin
          saturatedCollectVector_0_query_branchMask <= saturatedCollectVector_1_query_branchMask; // @[missHandler.scala 148:32]
        end
      end else begin
        saturatedCollectVector_0_query_branchMask <= saturatedCollectVector_1_query_branchMask; // @[missHandler.scala 148:32]
      end
    end else if (branchOps_valid) begin // @[missHandler.scala 149:47]
      if (|_T_79) begin // @[missHandler.scala 150:90]
        saturatedCollectVector_0_query_branchMask <= _saturatedCollectVectorUpdate_0_query_branchMask_T; // @[missHandler.scala 150:115]
      end
    end
    if (~saturated) begin // @[missHandler.scala 131:26]
      if (_T_72) begin // @[missHandler.scala 137:19]
        saturatedCollectVector_0_query_robAddr <= missedRequest_query_robAddr; // @[missHandler.scala 138:51]
      end
    end else if (~saturatedCollectVector_0_query_valid) begin // @[missHandler.scala 158:117]
      saturatedCollectVector_0_query_robAddr <= saturatedCollectVector_1_query_robAddr; // @[missHandler.scala 158:123]
    end
    if (~saturated) begin // @[missHandler.scala 131:26]
      if (_T_72) begin // @[missHandler.scala 137:19]
        saturatedCollectVector_0_query_prfDest <= missedRequest_query_prfDest; // @[missHandler.scala 138:51]
      end
    end else if (~saturatedCollectVector_0_query_valid) begin // @[missHandler.scala 158:117]
      saturatedCollectVector_0_query_prfDest <= saturatedCollectVector_1_query_prfDest; // @[missHandler.scala 158:123]
    end
    if (~saturated) begin // @[missHandler.scala 131:26]
      if (_T_72) begin // @[missHandler.scala 137:19]
        saturatedCollectVector_0_data <= missedRequest_data; // @[missHandler.scala 138:51]
      end
    end else if (~saturatedCollectVector_0_query_valid) begin // @[missHandler.scala 158:117]
      saturatedCollectVector_0_data <= saturatedCollectVector_1_data; // @[missHandler.scala 158:123]
    end
    if (reset) begin // @[missHandler.scala 81:39]
      saturatedCollectVector_1_query_valid <= 1'h0; // @[missHandler.scala 81:39]
    end else if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (_T_31) begin // @[missHandler.scala 160:132]
        saturatedCollectVector_1_query_valid <= 1'h0; // @[missHandler.scala 161:70]
      end else if (~saturatedCollectVector_0_query_valid | ~saturatedCollectVector_1_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_1_query_valid <= saturatedCollectVectorUpdate_2_query_valid; // @[missHandler.scala 158:123]
      end else begin
        saturatedCollectVector_1_query_valid <= saturatedCollectVectorUpdate_1_query_valid; // @[missHandler.scala 158:149]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~saturatedCollectVector_0_query_valid | ~saturatedCollectVector_1_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_1_query_address <= saturatedCollectVector_2_query_address; // @[missHandler.scala 158:123]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~saturatedCollectVector_0_query_valid | ~saturatedCollectVector_1_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_1_query_instruction <= saturatedCollectVector_2_query_instruction; // @[missHandler.scala 158:123]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~saturatedCollectVector_0_query_valid | ~saturatedCollectVector_1_query_valid) begin // @[missHandler.scala 158:117]
        if (branchOps_valid) begin // @[missHandler.scala 149:47]
          if (|_T_91) begin // @[missHandler.scala 150:90]
            saturatedCollectVector_1_query_branchMask <= _saturatedCollectVectorUpdate_2_query_branchMask_T; // @[missHandler.scala 150:115]
          end else begin
            saturatedCollectVector_1_query_branchMask <= saturatedCollectVector_2_query_branchMask; // @[missHandler.scala 148:32]
          end
        end else begin
          saturatedCollectVector_1_query_branchMask <= saturatedCollectVector_2_query_branchMask; // @[missHandler.scala 148:32]
        end
      end else if (branchOps_valid) begin // @[missHandler.scala 149:47]
        if (|_T_85) begin // @[missHandler.scala 150:90]
          saturatedCollectVector_1_query_branchMask <= _saturatedCollectVectorUpdate_1_query_branchMask_T; // @[missHandler.scala 150:115]
        end
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~saturatedCollectVector_0_query_valid | ~saturatedCollectVector_1_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_1_query_robAddr <= saturatedCollectVector_2_query_robAddr; // @[missHandler.scala 158:123]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~saturatedCollectVector_0_query_valid | ~saturatedCollectVector_1_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_1_query_prfDest <= saturatedCollectVector_2_query_prfDest; // @[missHandler.scala 158:123]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~saturatedCollectVector_0_query_valid | ~saturatedCollectVector_1_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_1_data <= saturatedCollectVector_2_data; // @[missHandler.scala 158:123]
      end
    end
    if (reset) begin // @[missHandler.scala 81:39]
      saturatedCollectVector_2_query_valid <= 1'h0; // @[missHandler.scala 81:39]
    end else if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (_T_31) begin // @[missHandler.scala 160:132]
        saturatedCollectVector_2_query_valid <= 1'h0; // @[missHandler.scala 161:70]
      end else if (~_T_116 | ~saturatedCollectVector_2_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_2_query_valid <= saturatedCollectVectorUpdate_3_query_valid; // @[missHandler.scala 158:123]
      end else begin
        saturatedCollectVector_2_query_valid <= saturatedCollectVectorUpdate_2_query_valid; // @[missHandler.scala 158:149]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~_T_116 | ~saturatedCollectVector_2_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_2_query_address <= saturatedCollectVector_3_query_address; // @[missHandler.scala 158:123]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~_T_116 | ~saturatedCollectVector_2_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_2_query_instruction <= saturatedCollectVector_3_query_instruction; // @[missHandler.scala 158:123]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~_T_116 | ~saturatedCollectVector_2_query_valid) begin // @[missHandler.scala 158:117]
        if (branchOps_valid) begin // @[missHandler.scala 149:47]
          if (|_T_97) begin // @[missHandler.scala 150:90]
            saturatedCollectVector_2_query_branchMask <= _saturatedCollectVectorUpdate_3_query_branchMask_T; // @[missHandler.scala 150:115]
          end else begin
            saturatedCollectVector_2_query_branchMask <= saturatedCollectVector_3_query_branchMask; // @[missHandler.scala 148:32]
          end
        end else begin
          saturatedCollectVector_2_query_branchMask <= saturatedCollectVector_3_query_branchMask; // @[missHandler.scala 148:32]
        end
      end else if (branchOps_valid) begin // @[missHandler.scala 149:47]
        if (|_T_91) begin // @[missHandler.scala 150:90]
          saturatedCollectVector_2_query_branchMask <= _saturatedCollectVectorUpdate_2_query_branchMask_T; // @[missHandler.scala 150:115]
        end
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~_T_116 | ~saturatedCollectVector_2_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_2_query_robAddr <= saturatedCollectVector_3_query_robAddr; // @[missHandler.scala 158:123]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~_T_116 | ~saturatedCollectVector_2_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_2_query_prfDest <= saturatedCollectVector_3_query_prfDest; // @[missHandler.scala 158:123]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~_T_116 | ~saturatedCollectVector_2_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_2_data <= saturatedCollectVector_3_data; // @[missHandler.scala 158:123]
      end
    end
    if (reset) begin // @[missHandler.scala 81:39]
      saturatedCollectVector_3_query_valid <= 1'h0; // @[missHandler.scala 81:39]
    end else if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (_T_31) begin // @[missHandler.scala 160:132]
        saturatedCollectVector_3_query_valid <= 1'h0; // @[missHandler.scala 161:70]
      end else if (~_T_117 | ~saturatedCollectVector_3_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_3_query_valid <= saturatedCollectVectorUpdate_4_query_valid; // @[missHandler.scala 158:123]
      end else begin
        saturatedCollectVector_3_query_valid <= saturatedCollectVectorUpdate_3_query_valid; // @[missHandler.scala 158:149]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~_T_117 | ~saturatedCollectVector_3_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_3_query_address <= saturatedCollectVector_4_query_address; // @[missHandler.scala 158:123]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~_T_117 | ~saturatedCollectVector_3_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_3_query_instruction <= saturatedCollectVector_4_query_instruction; // @[missHandler.scala 158:123]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~_T_117 | ~saturatedCollectVector_3_query_valid) begin // @[missHandler.scala 158:117]
        if (branchOps_valid) begin // @[missHandler.scala 149:47]
          if (|_T_103) begin // @[missHandler.scala 150:90]
            saturatedCollectVector_3_query_branchMask <= _saturatedCollectVectorUpdate_4_query_branchMask_T; // @[missHandler.scala 150:115]
          end else begin
            saturatedCollectVector_3_query_branchMask <= saturatedCollectVector_4_query_branchMask; // @[missHandler.scala 148:32]
          end
        end else begin
          saturatedCollectVector_3_query_branchMask <= saturatedCollectVector_4_query_branchMask; // @[missHandler.scala 148:32]
        end
      end else if (branchOps_valid) begin // @[missHandler.scala 149:47]
        if (|_T_97) begin // @[missHandler.scala 150:90]
          saturatedCollectVector_3_query_branchMask <= _saturatedCollectVectorUpdate_3_query_branchMask_T; // @[missHandler.scala 150:115]
        end
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~_T_117 | ~saturatedCollectVector_3_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_3_query_robAddr <= saturatedCollectVector_4_query_robAddr; // @[missHandler.scala 158:123]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~_T_117 | ~saturatedCollectVector_3_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_3_query_prfDest <= saturatedCollectVector_4_query_prfDest; // @[missHandler.scala 158:123]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~_T_117 | ~saturatedCollectVector_3_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_3_data <= saturatedCollectVector_4_data; // @[missHandler.scala 158:123]
      end
    end
    if (reset) begin // @[missHandler.scala 81:39]
      saturatedCollectVector_4_query_valid <= 1'h0; // @[missHandler.scala 81:39]
    end else if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (_T_31) begin // @[missHandler.scala 160:132]
        saturatedCollectVector_4_query_valid <= 1'h0; // @[missHandler.scala 161:70]
      end else if (~_T_118 | ~saturatedCollectVector_4_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_4_query_valid <= _GEN_75; // @[missHandler.scala 158:123]
      end else begin
        saturatedCollectVector_4_query_valid <= saturatedCollectVectorUpdate_4_query_valid; // @[missHandler.scala 158:149]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~_T_118 | ~saturatedCollectVector_4_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_4_query_address <= missedRequest_query_address; // @[missHandler.scala 158:123]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~_T_118 | ~saturatedCollectVector_4_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_4_query_instruction <= missedRequest_query_instruction; // @[missHandler.scala 158:123]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~_T_118 | ~saturatedCollectVector_4_query_valid) begin // @[missHandler.scala 158:117]
        if (branchOps_valid) begin // @[missHandler.scala 140:47]
          if (|_T_73) begin // @[missHandler.scala 141:99]
            saturatedCollectVector_4_query_branchMask <= _saturatedCollectVector_0_query_branchMask_T; // @[missHandler.scala 141:143]
          end else begin
            saturatedCollectVector_4_query_branchMask <= missedRequest_query_branchMask; // @[missHandler.scala 138:51]
          end
        end else begin
          saturatedCollectVector_4_query_branchMask <= missedRequest_query_branchMask; // @[missHandler.scala 138:51]
        end
      end else if (branchOps_valid) begin // @[missHandler.scala 149:47]
        if (|_T_103) begin // @[missHandler.scala 150:90]
          saturatedCollectVector_4_query_branchMask <= _saturatedCollectVectorUpdate_4_query_branchMask_T; // @[missHandler.scala 150:115]
        end
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~_T_118 | ~saturatedCollectVector_4_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_4_query_robAddr <= missedRequest_query_robAddr; // @[missHandler.scala 158:123]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~_T_118 | ~saturatedCollectVector_4_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_4_query_prfDest <= missedRequest_query_prfDest; // @[missHandler.scala 158:123]
      end
    end
    if (!(~saturated)) begin // @[missHandler.scala 131:26]
      if (~_T_118 | ~saturatedCollectVector_4_query_valid) begin // @[missHandler.scala 158:117]
        saturatedCollectVector_4_data <= missedRequest_data; // @[missHandler.scala 158:123]
      end
    end
    if (reset) begin // @[missHandler.scala 83:35]
      nonSaturatedMisses_0_query_valid <= 1'h0; // @[missHandler.scala 83:35]
    end else if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_valid <= _GEN_270;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_valid <= _GEN_270;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_valid <= _GEN_270;
    end else begin
      nonSaturatedMisses_0_query_valid <= _GEN_306;
    end
    if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_address <= _GEN_271;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_address <= _GEN_271;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_address <= _GEN_271;
    end else if (2'h3 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_address <= nonSaturatedMisses_1_query_address; // @[missHandler.scala 358:107]
    end else begin
      nonSaturatedMisses_0_query_address <= _GEN_271;
    end
    if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_instruction <= _GEN_272;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_instruction <= _GEN_272;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_instruction <= _GEN_272;
    end else if (2'h3 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_instruction <= nonSaturatedMisses_1_query_instruction; // @[missHandler.scala 358:107]
    end else begin
      nonSaturatedMisses_0_query_instruction <= _GEN_272;
    end
    if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_branchMask <= _GEN_273;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_branchMask <= _GEN_273;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_branchMask <= _GEN_273;
    end else if (2'h3 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_branchMask <= nonSaturatedMisses_1_query_branchMask; // @[missHandler.scala 358:107]
    end else begin
      nonSaturatedMisses_0_query_branchMask <= _GEN_273;
    end
    if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_robAddr <= _GEN_274;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_robAddr <= _GEN_274;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_robAddr <= _GEN_274;
    end else if (2'h3 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_robAddr <= nonSaturatedMisses_1_query_robAddr; // @[missHandler.scala 358:107]
    end else begin
      nonSaturatedMisses_0_query_robAddr <= _GEN_274;
    end
    if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_prfDest <= _GEN_275;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_prfDest <= _GEN_275;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_prfDest <= _GEN_275;
    end else if (2'h3 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_query_prfDest <= nonSaturatedMisses_1_query_prfDest; // @[missHandler.scala 358:107]
    end else begin
      nonSaturatedMisses_0_query_prfDest <= _GEN_275;
    end
    if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_data <= _GEN_276;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_data <= _GEN_276;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_data <= _GEN_276;
    end else if (2'h3 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_0_data <= nonSaturatedMisses_1_data; // @[missHandler.scala 358:107]
    end else begin
      nonSaturatedMisses_0_data <= _GEN_276;
    end
    if (reset) begin // @[missHandler.scala 83:35]
      nonSaturatedMisses_1_query_valid <= 1'h0; // @[missHandler.scala 83:35]
    end else if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_valid <= _GEN_277;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_valid <= _GEN_277;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_valid <= _GEN_277;
    end else begin
      nonSaturatedMisses_1_query_valid <= _GEN_313;
    end
    if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_address <= _GEN_278;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_address <= _GEN_278;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_address <= _GEN_278;
    end else if (2'h3 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_address <= nonSaturatedMisses_2_query_address; // @[missHandler.scala 358:107]
    end else begin
      nonSaturatedMisses_1_query_address <= _GEN_278;
    end
    if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_instruction <= _GEN_279;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_instruction <= _GEN_279;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_instruction <= _GEN_279;
    end else if (2'h3 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_instruction <= nonSaturatedMisses_2_query_instruction; // @[missHandler.scala 358:107]
    end else begin
      nonSaturatedMisses_1_query_instruction <= _GEN_279;
    end
    if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_branchMask <= _GEN_280;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_branchMask <= _GEN_280;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_branchMask <= _GEN_280;
    end else if (2'h3 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_branchMask <= nonSaturatedMisses_2_query_branchMask; // @[missHandler.scala 358:107]
    end else begin
      nonSaturatedMisses_1_query_branchMask <= _GEN_280;
    end
    if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_robAddr <= _GEN_281;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_robAddr <= _GEN_281;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_robAddr <= _GEN_281;
    end else if (2'h3 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_robAddr <= nonSaturatedMisses_2_query_robAddr; // @[missHandler.scala 358:107]
    end else begin
      nonSaturatedMisses_1_query_robAddr <= _GEN_281;
    end
    if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_prfDest <= _GEN_282;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_prfDest <= _GEN_282;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_prfDest <= _GEN_282;
    end else if (2'h3 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_query_prfDest <= nonSaturatedMisses_2_query_prfDest; // @[missHandler.scala 358:107]
    end else begin
      nonSaturatedMisses_1_query_prfDest <= _GEN_282;
    end
    if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_data <= _GEN_283;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_data <= _GEN_283;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_data <= _GEN_283;
    end else if (2'h3 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_1_data <= nonSaturatedMisses_2_data; // @[missHandler.scala 358:107]
    end else begin
      nonSaturatedMisses_1_data <= _GEN_283;
    end
    if (reset) begin // @[missHandler.scala 83:35]
      nonSaturatedMisses_2_query_valid <= 1'h0; // @[missHandler.scala 83:35]
    end else if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_valid <= _GEN_284;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_valid <= _GEN_284;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_valid <= _GEN_284;
    end else begin
      nonSaturatedMisses_2_query_valid <= _GEN_320;
    end
    if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_address <= _GEN_285;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_address <= _GEN_285;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_address <= _GEN_285;
    end else if (2'h3 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_address <= nonSaturatedMisses_3_query_address; // @[missHandler.scala 358:107]
    end else begin
      nonSaturatedMisses_2_query_address <= _GEN_285;
    end
    if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_instruction <= _GEN_286;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_instruction <= _GEN_286;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_instruction <= _GEN_286;
    end else if (2'h3 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_instruction <= nonSaturatedMisses_3_query_instruction; // @[missHandler.scala 358:107]
    end else begin
      nonSaturatedMisses_2_query_instruction <= _GEN_286;
    end
    if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_branchMask <= _GEN_287;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_branchMask <= _GEN_287;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_branchMask <= _GEN_287;
    end else if (2'h3 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_branchMask <= nonSaturatedMisses_3_query_branchMask; // @[missHandler.scala 358:107]
    end else begin
      nonSaturatedMisses_2_query_branchMask <= _GEN_287;
    end
    if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_robAddr <= _GEN_288;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_robAddr <= _GEN_288;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_robAddr <= _GEN_288;
    end else if (2'h3 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_robAddr <= nonSaturatedMisses_3_query_robAddr; // @[missHandler.scala 358:107]
    end else begin
      nonSaturatedMisses_2_query_robAddr <= _GEN_288;
    end
    if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_prfDest <= _GEN_289;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_prfDest <= _GEN_289;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_prfDest <= _GEN_289;
    end else if (2'h3 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_query_prfDest <= nonSaturatedMisses_3_query_prfDest; // @[missHandler.scala 358:107]
    end else begin
      nonSaturatedMisses_2_query_prfDest <= _GEN_289;
    end
    if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_data <= _GEN_290;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_data <= _GEN_290;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_data <= _GEN_290;
    end else if (2'h3 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_2_data <= nonSaturatedMisses_3_data; // @[missHandler.scala 358:107]
    end else begin
      nonSaturatedMisses_2_data <= _GEN_290;
    end
    if (reset) begin // @[missHandler.scala 83:35]
      nonSaturatedMisses_3_query_valid <= 1'h0; // @[missHandler.scala 83:35]
    end else if (_T_144) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_3_query_valid <= _GEN_291;
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_3_query_valid <= _GEN_291;
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      nonSaturatedMisses_3_query_valid <= _GEN_291;
    end else begin
      nonSaturatedMisses_3_query_valid <= _GEN_327;
    end
    if (_T_63) begin // @[missHandler.scala 282:38]
      if (~_T_69 | ~nonSaturatedMisses_3_query_valid) begin // @[missHandler.scala 297:119]
        nonSaturatedMisses_3_query_address <= missedRequest_query_address; // @[missHandler.scala 297:125]
      end
    end
    if (_T_63) begin // @[missHandler.scala 282:38]
      if (~_T_69 | ~nonSaturatedMisses_3_query_valid) begin // @[missHandler.scala 297:119]
        nonSaturatedMisses_3_query_instruction <= missedRequest_query_instruction; // @[missHandler.scala 297:125]
      end
    end
    if (_T_63) begin // @[missHandler.scala 282:38]
      if (~_T_69 | ~nonSaturatedMisses_3_query_valid) begin // @[missHandler.scala 297:119]
        if (branchOps_valid) begin // @[missHandler.scala 140:47]
          if (|_T_73) begin // @[missHandler.scala 141:99]
            nonSaturatedMisses_3_query_branchMask <= _saturatedCollectVector_0_query_branchMask_T; // @[missHandler.scala 141:143]
          end else begin
            nonSaturatedMisses_3_query_branchMask <= missedRequest_query_branchMask; // @[missHandler.scala 138:51]
          end
        end else begin
          nonSaturatedMisses_3_query_branchMask <= missedRequest_query_branchMask; // @[missHandler.scala 138:51]
        end
      end else if (branchOps_valid) begin // @[missHandler.scala 286:47]
        if (|_T_188) begin // @[missHandler.scala 287:90]
          nonSaturatedMisses_3_query_branchMask <= _nonSaturatedMissesUpdate_3_query_branchMask_T; // @[missHandler.scala 287:115]
        end
      end
    end
    if (_T_63) begin // @[missHandler.scala 282:38]
      if (~_T_69 | ~nonSaturatedMisses_3_query_valid) begin // @[missHandler.scala 297:119]
        nonSaturatedMisses_3_query_robAddr <= missedRequest_query_robAddr; // @[missHandler.scala 297:125]
      end
    end
    if (_T_63) begin // @[missHandler.scala 282:38]
      if (~_T_69 | ~nonSaturatedMisses_3_query_valid) begin // @[missHandler.scala 297:119]
        nonSaturatedMisses_3_query_prfDest <= missedRequest_query_prfDest; // @[missHandler.scala 297:125]
      end
    end
    if (_T_63) begin // @[missHandler.scala 282:38]
      if (~_T_69 | ~nonSaturatedMisses_3_query_valid) begin // @[missHandler.scala 297:119]
        nonSaturatedMisses_3_data <= missedRequest_data; // @[missHandler.scala 297:125]
      end
    end
    if (reset) begin // @[missHandler.scala 86:30]
      handlerStatus <= 2'h0; // @[missHandler.scala 86:30]
    end else if (_T_144) begin // @[missHandler.scala 340:31]
      if (missedRequest_query_valid) begin // @[missHandler.scala 342:57]
        handlerStatus <= 2'h1; // @[missHandler.scala 343:47]
      end
    end else if (_T_145) begin // @[missHandler.scala 340:31]
      if (_rlastToCache_T_1 & pushToCache_fired) begin // @[missHandler.scala 348:94]
        handlerStatus <= 2'h2; // @[missHandler.scala 348:110]
      end
    end else if (2'h2 == handlerStatus) begin // @[missHandler.scala 340:31]
      handlerStatus <= _GEN_303;
    end else begin
      handlerStatus <= _GEN_305;
    end
    if (reset) begin // @[missHandler.scala 88:32]
      saturated <= 1'h0; // @[missHandler.scala 88:32]
    end else if (~saturated) begin // @[missHandler.scala 131:26]
      saturated <= _GEN_83;
    end else if (_T_31) begin // @[missHandler.scala 160:132]
      saturated <= 1'h0; // @[missHandler.scala 162:35]
    end
    if (_T_144) begin // @[missHandler.scala 340:31]
      if (missedRequest_query_valid) begin // @[missHandler.scala 342:57]
        servicingBlock <= _servicingBlock_T_1; // @[missHandler.scala 344:48]
      end
    end
    if (pushToCache_fired | ~cacheWrite_valid) begin // @[missHandler.scala 185:54]
      cacheWrite_data <= _cacheWrite_data_T; // @[missHandler.scala 186:33]
    end
    if (reset) begin // @[missHandler.scala 166:33]
      cacheWrite_valid <= 1'h0; // @[missHandler.scala 166:33]
    end else if (pushToCache_fired | ~cacheWrite_valid) begin // @[missHandler.scala 185:54]
      cacheWrite_valid <= fetched_0_valid & fetched_1_valid; // @[missHandler.scala 187:34]
    end
    cacheWrite_address <= _GEN_190[8:0];
    cacheWrite_setSelVector <= nextSet; // @[missHandler.scala 301:33]
    if (axi_RREADY & axi_RVALID) begin // @[missHandler.scala 205:40]
      if (_T_143 & _cacheWrite_valid_T) begin // @[missHandler.scala 206:103]
        fetched_0_rdata <= axi_RDATA; // @[missHandler.scala 208:42]
      end else if (~fetched_0_valid) begin // @[missHandler.scala 210:46]
        fetched_0_rdata <= axi_RDATA; // @[missHandler.scala 211:42]
      end
    end
    if (reset) begin // @[missHandler.scala 173:30]
      fetched_0_valid <= 1'h0; // @[missHandler.scala 173:30]
    end else if (axi_RREADY & axi_RVALID) begin // @[missHandler.scala 205:40]
      fetched_0_valid <= _GEN_197;
    end else if (_T_150) begin // @[missHandler.scala 217:101]
      fetched_0_valid <= 1'h0; // @[missHandler.scala 218:34]
    end
    if (axi_RREADY & axi_RVALID) begin // @[missHandler.scala 205:40]
      if (!(_T_143 & _cacheWrite_valid_T)) begin // @[missHandler.scala 206:103]
        if (!(~fetched_0_valid)) begin // @[missHandler.scala 210:46]
          fetched_1_rdata <= axi_RDATA; // @[missHandler.scala 214:42]
        end
      end
    end
    if (reset) begin // @[missHandler.scala 173:30]
      fetched_1_valid <= 1'h0; // @[missHandler.scala 173:30]
    end else if (axi_RREADY & axi_RVALID) begin // @[missHandler.scala 205:40]
      if (_T_143 & _cacheWrite_valid_T) begin // @[missHandler.scala 206:103]
        fetched_1_valid <= 1'h0; // @[missHandler.scala 207:42]
      end else if (!(~fetched_0_valid)) begin // @[missHandler.scala 210:46]
        fetched_1_valid <= 1'h1; // @[missHandler.scala 215:42]
      end
    end else if (_T_150) begin // @[missHandler.scala 217:101]
      fetched_1_valid <= 1'h0; // @[missHandler.scala 219:34]
    end
    if (reset) begin // @[missHandler.scala 224:35]
      clearToFetch <= 1'h0; // @[missHandler.scala 224:35]
    end else if (~clearToFetch) begin // @[missHandler.scala 242:29]
      if (_dependencyCheck_requset_valid_T) begin // @[missHandler.scala 243:51]
        clearToFetch <= dependencyCheck_free | clearToFetch;
      end
    end else begin
      clearToFetch <= _T_63; // @[missHandler.scala 244:36]
    end
    if (reset) begin // @[missHandler.scala 237:32]
      requested <= 1'h0; // @[missHandler.scala 237:32]
    end else if (~requested) begin // @[missHandler.scala 239:26]
      requested <= axi_ARVALID & axi_ARREADY; // @[missHandler.scala 239:38]
    end else begin
      requested <= _T_63; // @[missHandler.scala 240:32]
    end
    if (reset) begin // @[missHandler.scala 246:38]
      arvalid <= 1'h0; // @[missHandler.scala 246:38]
    end else if (~arvalid) begin // @[missHandler.scala 247:25]
      arvalid <= _T_156 & clearToFetch; // @[missHandler.scala 247:35]
    end else begin
      arvalid <= ~_requested_T; // @[missHandler.scala 248:30]
    end
    if (reset) begin // @[missHandler.scala 246:38]
      rready <= 1'h0; // @[missHandler.scala 246:38]
    end else if (~rready) begin // @[missHandler.scala 250:24]
      rready <= _requested_T; // @[missHandler.scala 250:33]
    end else begin
      rready <= ~(axi_RVALID & axi_RREADY & axi_RLAST); // @[missHandler.scala 251:29]
    end
    if (handlerStatus == 2'h0) begin // @[missHandler.scala 322:38]
      if (missedRequest_query_valid) begin // @[missHandler.scala 323:50]
        if (_setInvalidateVector_T) begin // @[missHandler.scala 316:35]
          nextSet <= randSelect;
        end else if (_setInvalidateVector_T_3) begin // @[Mux.scala 101:16]
          nextSet <= 2'h1;
        end else begin
          nextSet <= _setInvalidateVector_T_7;
        end
      end
    end
    if (reset) begin // @[missHandler.scala 304:33]
      randSelect <= 2'h1; // @[missHandler.scala 304:33]
    end else if (randSelect[0]) begin // @[missHandler.scala 305:26]
      randSelect <= 2'h2;
    end else begin
      randSelect <= {{1'd0}, randSelect[1]};
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  saturatedReplayVector_0_query_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  saturatedReplayVector_0_query_address = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  saturatedReplayVector_0_query_instruction = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  saturatedReplayVector_0_query_branchMask = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  saturatedReplayVector_0_query_robAddr = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  saturatedReplayVector_0_query_prfDest = _RAND_5[5:0];
  _RAND_6 = {2{`RANDOM}};
  saturatedReplayVector_0_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  saturatedReplayVector_1_query_valid = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  saturatedReplayVector_1_query_address = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  saturatedReplayVector_1_query_instruction = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  saturatedReplayVector_1_query_branchMask = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  saturatedReplayVector_1_query_robAddr = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  saturatedReplayVector_1_query_prfDest = _RAND_12[5:0];
  _RAND_13 = {2{`RANDOM}};
  saturatedReplayVector_1_data = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  saturatedReplayVector_2_query_valid = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  saturatedReplayVector_2_query_address = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  saturatedReplayVector_2_query_instruction = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  saturatedReplayVector_2_query_branchMask = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  saturatedReplayVector_2_query_robAddr = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  saturatedReplayVector_2_query_prfDest = _RAND_19[5:0];
  _RAND_20 = {2{`RANDOM}};
  saturatedReplayVector_2_data = _RAND_20[63:0];
  _RAND_21 = {1{`RANDOM}};
  saturatedReplayVector_3_query_valid = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  saturatedReplayVector_3_query_address = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  saturatedReplayVector_3_query_instruction = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  saturatedReplayVector_3_query_branchMask = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  saturatedReplayVector_3_query_robAddr = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  saturatedReplayVector_3_query_prfDest = _RAND_26[5:0];
  _RAND_27 = {2{`RANDOM}};
  saturatedReplayVector_3_data = _RAND_27[63:0];
  _RAND_28 = {1{`RANDOM}};
  saturatedReplayVector_4_query_valid = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  saturatedReplayVector_4_query_address = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  saturatedReplayVector_4_query_instruction = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  saturatedReplayVector_4_query_branchMask = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  saturatedReplayVector_4_query_robAddr = _RAND_32[3:0];
  _RAND_33 = {1{`RANDOM}};
  saturatedReplayVector_4_query_prfDest = _RAND_33[5:0];
  _RAND_34 = {2{`RANDOM}};
  saturatedReplayVector_4_data = _RAND_34[63:0];
  _RAND_35 = {1{`RANDOM}};
  saturatedCollectVector_0_query_valid = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  saturatedCollectVector_0_query_address = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  saturatedCollectVector_0_query_instruction = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  saturatedCollectVector_0_query_branchMask = _RAND_38[3:0];
  _RAND_39 = {1{`RANDOM}};
  saturatedCollectVector_0_query_robAddr = _RAND_39[3:0];
  _RAND_40 = {1{`RANDOM}};
  saturatedCollectVector_0_query_prfDest = _RAND_40[5:0];
  _RAND_41 = {2{`RANDOM}};
  saturatedCollectVector_0_data = _RAND_41[63:0];
  _RAND_42 = {1{`RANDOM}};
  saturatedCollectVector_1_query_valid = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  saturatedCollectVector_1_query_address = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  saturatedCollectVector_1_query_instruction = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  saturatedCollectVector_1_query_branchMask = _RAND_45[3:0];
  _RAND_46 = {1{`RANDOM}};
  saturatedCollectVector_1_query_robAddr = _RAND_46[3:0];
  _RAND_47 = {1{`RANDOM}};
  saturatedCollectVector_1_query_prfDest = _RAND_47[5:0];
  _RAND_48 = {2{`RANDOM}};
  saturatedCollectVector_1_data = _RAND_48[63:0];
  _RAND_49 = {1{`RANDOM}};
  saturatedCollectVector_2_query_valid = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  saturatedCollectVector_2_query_address = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  saturatedCollectVector_2_query_instruction = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  saturatedCollectVector_2_query_branchMask = _RAND_52[3:0];
  _RAND_53 = {1{`RANDOM}};
  saturatedCollectVector_2_query_robAddr = _RAND_53[3:0];
  _RAND_54 = {1{`RANDOM}};
  saturatedCollectVector_2_query_prfDest = _RAND_54[5:0];
  _RAND_55 = {2{`RANDOM}};
  saturatedCollectVector_2_data = _RAND_55[63:0];
  _RAND_56 = {1{`RANDOM}};
  saturatedCollectVector_3_query_valid = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  saturatedCollectVector_3_query_address = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  saturatedCollectVector_3_query_instruction = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  saturatedCollectVector_3_query_branchMask = _RAND_59[3:0];
  _RAND_60 = {1{`RANDOM}};
  saturatedCollectVector_3_query_robAddr = _RAND_60[3:0];
  _RAND_61 = {1{`RANDOM}};
  saturatedCollectVector_3_query_prfDest = _RAND_61[5:0];
  _RAND_62 = {2{`RANDOM}};
  saturatedCollectVector_3_data = _RAND_62[63:0];
  _RAND_63 = {1{`RANDOM}};
  saturatedCollectVector_4_query_valid = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  saturatedCollectVector_4_query_address = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  saturatedCollectVector_4_query_instruction = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  saturatedCollectVector_4_query_branchMask = _RAND_66[3:0];
  _RAND_67 = {1{`RANDOM}};
  saturatedCollectVector_4_query_robAddr = _RAND_67[3:0];
  _RAND_68 = {1{`RANDOM}};
  saturatedCollectVector_4_query_prfDest = _RAND_68[5:0];
  _RAND_69 = {2{`RANDOM}};
  saturatedCollectVector_4_data = _RAND_69[63:0];
  _RAND_70 = {1{`RANDOM}};
  nonSaturatedMisses_0_query_valid = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  nonSaturatedMisses_0_query_address = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  nonSaturatedMisses_0_query_instruction = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  nonSaturatedMisses_0_query_branchMask = _RAND_73[3:0];
  _RAND_74 = {1{`RANDOM}};
  nonSaturatedMisses_0_query_robAddr = _RAND_74[3:0];
  _RAND_75 = {1{`RANDOM}};
  nonSaturatedMisses_0_query_prfDest = _RAND_75[5:0];
  _RAND_76 = {2{`RANDOM}};
  nonSaturatedMisses_0_data = _RAND_76[63:0];
  _RAND_77 = {1{`RANDOM}};
  nonSaturatedMisses_1_query_valid = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  nonSaturatedMisses_1_query_address = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  nonSaturatedMisses_1_query_instruction = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  nonSaturatedMisses_1_query_branchMask = _RAND_80[3:0];
  _RAND_81 = {1{`RANDOM}};
  nonSaturatedMisses_1_query_robAddr = _RAND_81[3:0];
  _RAND_82 = {1{`RANDOM}};
  nonSaturatedMisses_1_query_prfDest = _RAND_82[5:0];
  _RAND_83 = {2{`RANDOM}};
  nonSaturatedMisses_1_data = _RAND_83[63:0];
  _RAND_84 = {1{`RANDOM}};
  nonSaturatedMisses_2_query_valid = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  nonSaturatedMisses_2_query_address = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  nonSaturatedMisses_2_query_instruction = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  nonSaturatedMisses_2_query_branchMask = _RAND_87[3:0];
  _RAND_88 = {1{`RANDOM}};
  nonSaturatedMisses_2_query_robAddr = _RAND_88[3:0];
  _RAND_89 = {1{`RANDOM}};
  nonSaturatedMisses_2_query_prfDest = _RAND_89[5:0];
  _RAND_90 = {2{`RANDOM}};
  nonSaturatedMisses_2_data = _RAND_90[63:0];
  _RAND_91 = {1{`RANDOM}};
  nonSaturatedMisses_3_query_valid = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  nonSaturatedMisses_3_query_address = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  nonSaturatedMisses_3_query_instruction = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  nonSaturatedMisses_3_query_branchMask = _RAND_94[3:0];
  _RAND_95 = {1{`RANDOM}};
  nonSaturatedMisses_3_query_robAddr = _RAND_95[3:0];
  _RAND_96 = {1{`RANDOM}};
  nonSaturatedMisses_3_query_prfDest = _RAND_96[5:0];
  _RAND_97 = {2{`RANDOM}};
  nonSaturatedMisses_3_data = _RAND_97[63:0];
  _RAND_98 = {1{`RANDOM}};
  handlerStatus = _RAND_98[1:0];
  _RAND_99 = {1{`RANDOM}};
  saturated = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  servicingBlock = _RAND_100[31:0];
  _RAND_101 = {2{`RANDOM}};
  cacheWrite_data = _RAND_101[63:0];
  _RAND_102 = {1{`RANDOM}};
  cacheWrite_valid = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  cacheWrite_address = _RAND_103[8:0];
  _RAND_104 = {1{`RANDOM}};
  cacheWrite_setSelVector = _RAND_104[1:0];
  _RAND_105 = {1{`RANDOM}};
  fetched_0_rdata = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  fetched_0_valid = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  fetched_1_rdata = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  fetched_1_valid = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  clearToFetch = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  requested = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  arvalid = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  rready = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  nextSet = _RAND_113[1:0];
  _RAND_114 = {1{`RANDOM}};
  randSelect = _RAND_114[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module writeHandler(
  input         clock,
  input         reset,
  input         itWasPeripheral,
  output        writeCommit_ready,
  input         writeCommit_fired,
  output [31:0] axi_AWADDR,
  output [7:0]  axi_AWLEN,
  output [2:0]  axi_AWSIZE,
  output        axi_AWVALID,
  input         axi_AWREADY,
  output [31:0] axi_WDATA,
  output [3:0]  axi_WSTRB,
  output        axi_WLAST,
  output        axi_WVALID,
  input         axi_WREADY,
  input         axi_BVALID,
  output        axi_BREADY,
  input         request_valid,
  input  [31:0] request_address,
  input  [31:0] request_instruction,
  input  [63:0] request_alignedData,
  input  [7:0]  request_mask,
  input         dependencyCheck_requset_valid,
  input  [31:0] dependencyCheck_requset_address,
  output        dependencyCheck_free,
  output        clean
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] addressQueue_0_status; // @[writeHandler.scala 17:29]
  reg [31:0] addressQueue_0_address; // @[writeHandler.scala 17:29]
  reg  addressQueue_0_len; // @[writeHandler.scala 17:29]
  reg [2:0] addressQueue_0_size; // @[writeHandler.scala 17:29]
  reg  addressQueue_0_becausePeripheral; // @[writeHandler.scala 17:29]
  reg [1:0] addressQueue_1_status; // @[writeHandler.scala 17:29]
  reg [31:0] addressQueue_1_address; // @[writeHandler.scala 17:29]
  reg  addressQueue_1_len; // @[writeHandler.scala 17:29]
  reg [2:0] addressQueue_1_size; // @[writeHandler.scala 17:29]
  reg  addressQueue_1_becausePeripheral; // @[writeHandler.scala 17:29]
  reg [1:0] addressQueue_2_status; // @[writeHandler.scala 17:29]
  reg [31:0] addressQueue_2_address; // @[writeHandler.scala 17:29]
  reg  addressQueue_2_len; // @[writeHandler.scala 17:29]
  reg [2:0] addressQueue_2_size; // @[writeHandler.scala 17:29]
  reg  addressQueue_2_becausePeripheral; // @[writeHandler.scala 17:29]
  reg [1:0] addressQueue_3_status; // @[writeHandler.scala 17:29]
  reg [31:0] addressQueue_3_address; // @[writeHandler.scala 17:29]
  reg  addressQueue_3_len; // @[writeHandler.scala 17:29]
  reg [2:0] addressQueue_3_size; // @[writeHandler.scala 17:29]
  reg  addressQueue_3_becausePeripheral; // @[writeHandler.scala 17:29]
  reg [1:0] allocatePointer; // @[writeHandler.scala 29:91]
  reg [1:0] queryInsertPointer; // @[writeHandler.scala 29:91]
  reg [1:0] queryIniatePointer; // @[writeHandler.scala 29:91]
  reg [1:0] deallocatePointer; // @[writeHandler.scala 29:91]
  wire [1:0] _GEN_1 = 2'h1 == allocatePointer ? addressQueue_1_status : addressQueue_0_status; // @[writeHandler.scala 32:{62,62}]
  wire [1:0] _GEN_2 = 2'h2 == allocatePointer ? addressQueue_2_status : _GEN_1; // @[writeHandler.scala 32:{62,62}]
  wire [1:0] _GEN_3 = 2'h3 == allocatePointer ? addressQueue_3_status : _GEN_2; // @[writeHandler.scala 32:{62,62}]
  wire [1:0] _GEN_4 = 2'h0 == allocatePointer ? 2'h1 : addressQueue_0_status; // @[writeHandler.scala 17:29 35:{42,42}]
  wire [1:0] _GEN_5 = 2'h1 == allocatePointer ? 2'h1 : addressQueue_1_status; // @[writeHandler.scala 17:29 35:{42,42}]
  wire [1:0] _GEN_6 = 2'h2 == allocatePointer ? 2'h1 : addressQueue_2_status; // @[writeHandler.scala 17:29 35:{42,42}]
  wire [1:0] _GEN_7 = 2'h3 == allocatePointer ? 2'h1 : addressQueue_3_status; // @[writeHandler.scala 17:29 35:{42,42}]
  wire [1:0] _T_1 = allocatePointer + 2'h1; // @[writeHandler.scala 36:34]
  wire  _GEN_8 = 2'h0 == _T_1 ? 1'h0 : addressQueue_0_becausePeripheral; // @[writeHandler.scala 17:29 36:{59,59}]
  wire  _GEN_9 = 2'h1 == _T_1 ? 1'h0 : addressQueue_1_becausePeripheral; // @[writeHandler.scala 17:29 36:{59,59}]
  wire  _GEN_10 = 2'h2 == _T_1 ? 1'h0 : addressQueue_2_becausePeripheral; // @[writeHandler.scala 17:29 36:{59,59}]
  wire  _GEN_11 = 2'h3 == _T_1 ? 1'h0 : addressQueue_3_becausePeripheral; // @[writeHandler.scala 17:29 36:{59,59}]
  wire [1:0] _GEN_12 = writeCommit_fired ? _GEN_4 : addressQueue_0_status; // @[writeHandler.scala 34:27 17:29]
  wire [1:0] _GEN_13 = writeCommit_fired ? _GEN_5 : addressQueue_1_status; // @[writeHandler.scala 34:27 17:29]
  wire [1:0] _GEN_14 = writeCommit_fired ? _GEN_6 : addressQueue_2_status; // @[writeHandler.scala 34:27 17:29]
  wire [1:0] _GEN_15 = writeCommit_fired ? _GEN_7 : addressQueue_3_status; // @[writeHandler.scala 34:27 17:29]
  wire  _GEN_16 = writeCommit_fired ? _GEN_8 : addressQueue_0_becausePeripheral; // @[writeHandler.scala 34:27 17:29]
  wire  _GEN_17 = writeCommit_fired ? _GEN_9 : addressQueue_1_becausePeripheral; // @[writeHandler.scala 34:27 17:29]
  wire  _GEN_18 = writeCommit_fired ? _GEN_10 : addressQueue_2_becausePeripheral; // @[writeHandler.scala 34:27 17:29]
  wire  _GEN_19 = writeCommit_fired ? _GEN_11 : addressQueue_3_becausePeripheral; // @[writeHandler.scala 34:27 17:29]
  wire [1:0] _GEN_21 = 2'h0 == queryInsertPointer ? 2'h2 : _GEN_12; // @[writeHandler.scala 48:{45,45}]
  wire [1:0] _GEN_22 = 2'h1 == queryInsertPointer ? 2'h2 : _GEN_13; // @[writeHandler.scala 48:{45,45}]
  wire [1:0] _GEN_23 = 2'h2 == queryInsertPointer ? 2'h2 : _GEN_14; // @[writeHandler.scala 48:{45,45}]
  wire [1:0] _GEN_24 = 2'h3 == queryInsertPointer ? 2'h2 : _GEN_15; // @[writeHandler.scala 48:{45,45}]
  wire  _addressQueue_len_T_1 = request_instruction[13:12] == 2'h3; // @[writeHandler.scala 50:74]
  wire [1:0] _queryInsertPointer_T_1 = queryInsertPointer + 2'h1; // @[writeHandler.scala 52:46]
  wire [1:0] _GEN_37 = request_valid ? _GEN_21 : _GEN_12; // @[writeHandler.scala 47:23]
  wire [1:0] _GEN_38 = request_valid ? _GEN_22 : _GEN_13; // @[writeHandler.scala 47:23]
  wire [1:0] _GEN_39 = request_valid ? _GEN_23 : _GEN_14; // @[writeHandler.scala 47:23]
  wire [1:0] _GEN_40 = request_valid ? _GEN_24 : _GEN_15; // @[writeHandler.scala 47:23]
  wire [1:0] _GEN_54 = 2'h0 == queryInsertPointer ? 2'h0 : _GEN_37; // @[writeHandler.scala 55:{45,45}]
  wire [1:0] _GEN_55 = 2'h1 == queryInsertPointer ? 2'h0 : _GEN_38; // @[writeHandler.scala 55:{45,45}]
  wire [1:0] _GEN_56 = 2'h2 == queryInsertPointer ? 2'h0 : _GEN_39; // @[writeHandler.scala 55:{45,45}]
  wire [1:0] _GEN_57 = 2'h3 == queryInsertPointer ? 2'h0 : _GEN_40; // @[writeHandler.scala 55:{45,45}]
  wire  _GEN_58 = 2'h0 == queryInsertPointer | _GEN_16; // @[writeHandler.scala 56:{56,56}]
  wire  _GEN_59 = 2'h1 == queryInsertPointer | _GEN_17; // @[writeHandler.scala 56:{56,56}]
  wire  _GEN_60 = 2'h2 == queryInsertPointer | _GEN_18; // @[writeHandler.scala 56:{56,56}]
  wire  _GEN_61 = 2'h3 == queryInsertPointer | _GEN_19; // @[writeHandler.scala 56:{56,56}]
  wire [1:0] _GEN_62 = itWasPeripheral ? _GEN_54 : _GEN_37; // @[writeHandler.scala 54:25]
  wire [1:0] _GEN_63 = itWasPeripheral ? _GEN_55 : _GEN_38; // @[writeHandler.scala 54:25]
  wire [1:0] _GEN_64 = itWasPeripheral ? _GEN_56 : _GEN_39; // @[writeHandler.scala 54:25]
  wire [1:0] _GEN_65 = itWasPeripheral ? _GEN_57 : _GEN_40; // @[writeHandler.scala 54:25]
  wire [1:0] _GEN_71 = 2'h0 == queryIniatePointer ? 2'h3 : _GEN_62; // @[writeHandler.scala 61:{45,45}]
  wire [1:0] _GEN_72 = 2'h1 == queryIniatePointer ? 2'h3 : _GEN_63; // @[writeHandler.scala 61:{45,45}]
  wire [1:0] _GEN_73 = 2'h2 == queryIniatePointer ? 2'h3 : _GEN_64; // @[writeHandler.scala 61:{45,45}]
  wire [1:0] _GEN_74 = 2'h3 == queryIniatePointer ? 2'h3 : _GEN_65; // @[writeHandler.scala 61:{45,45}]
  wire [1:0] _queryIniatePointer_T_1 = queryIniatePointer + 2'h1; // @[writeHandler.scala 62:46]
  wire [1:0] _GEN_75 = axi_AWVALID & axi_AWREADY ? _GEN_71 : _GEN_62; // @[writeHandler.scala 60:36]
  wire [1:0] _GEN_76 = axi_AWVALID & axi_AWREADY ? _GEN_72 : _GEN_63; // @[writeHandler.scala 60:36]
  wire [1:0] _GEN_77 = axi_AWVALID & axi_AWREADY ? _GEN_73 : _GEN_64; // @[writeHandler.scala 60:36]
  wire [1:0] _GEN_78 = axi_AWVALID & axi_AWREADY ? _GEN_74 : _GEN_65; // @[writeHandler.scala 60:36]
  wire [1:0] _GEN_81 = 2'h1 == queryIniatePointer ? addressQueue_1_status : addressQueue_0_status; // @[writeHandler.scala 64:{49,49}]
  wire [1:0] _GEN_82 = 2'h2 == queryIniatePointer ? addressQueue_2_status : _GEN_81; // @[writeHandler.scala 64:{49,49}]
  wire [1:0] _GEN_83 = 2'h3 == queryIniatePointer ? addressQueue_3_status : _GEN_82; // @[writeHandler.scala 64:{49,49}]
  wire  _GEN_85 = 2'h1 == queryIniatePointer ? addressQueue_1_becausePeripheral : addressQueue_0_becausePeripheral; // @[writeHandler.scala 64:{67,67}]
  wire  _GEN_86 = 2'h2 == queryIniatePointer ? addressQueue_2_becausePeripheral : _GEN_85; // @[writeHandler.scala 64:{67,67}]
  wire  _GEN_87 = 2'h3 == queryIniatePointer ? addressQueue_3_becausePeripheral : _GEN_86; // @[writeHandler.scala 64:{67,67}]
  wire [1:0] _deallocatePointer_T_1 = deallocatePointer + 2'h1; // @[writeHandler.scala 70:44]
  wire [1:0] _GEN_99 = 2'h1 == deallocatePointer ? addressQueue_1_status : addressQueue_0_status; // @[writeHandler.scala 72:{48,48}]
  wire [1:0] _GEN_100 = 2'h2 == deallocatePointer ? addressQueue_2_status : _GEN_99; // @[writeHandler.scala 72:{48,48}]
  wire [1:0] _GEN_101 = 2'h3 == deallocatePointer ? addressQueue_3_status : _GEN_100; // @[writeHandler.scala 72:{48,48}]
  wire  _GEN_103 = 2'h1 == deallocatePointer ? addressQueue_1_becausePeripheral : addressQueue_0_becausePeripheral; // @[writeHandler.scala 72:{66,66}]
  wire  _GEN_104 = 2'h2 == deallocatePointer ? addressQueue_2_becausePeripheral : _GEN_103; // @[writeHandler.scala 72:{66,66}]
  wire  _GEN_105 = 2'h3 == deallocatePointer ? addressQueue_3_becausePeripheral : _GEN_104; // @[writeHandler.scala 72:{66,66}]
  reg  dataQueue_0_wvalid; // @[writeHandler.scala 76:26]
  reg  dataQueue_0_wlast; // @[writeHandler.scala 76:26]
  reg [31:0] dataQueue_0_wdata; // @[writeHandler.scala 76:26]
  reg [3:0] dataQueue_0_wstrb; // @[writeHandler.scala 76:26]
  reg  dataQueue_1_wvalid; // @[writeHandler.scala 76:26]
  reg  dataQueue_1_wlast; // @[writeHandler.scala 76:26]
  reg [31:0] dataQueue_1_wdata; // @[writeHandler.scala 76:26]
  reg [3:0] dataQueue_1_wstrb; // @[writeHandler.scala 76:26]
  reg  dataQueue_2_wvalid; // @[writeHandler.scala 76:26]
  reg  dataQueue_2_wlast; // @[writeHandler.scala 76:26]
  reg [31:0] dataQueue_2_wdata; // @[writeHandler.scala 76:26]
  reg [3:0] dataQueue_2_wstrb; // @[writeHandler.scala 76:26]
  reg  dataQueue_3_wvalid; // @[writeHandler.scala 76:26]
  reg  dataQueue_3_wlast; // @[writeHandler.scala 76:26]
  reg [31:0] dataQueue_3_wdata; // @[writeHandler.scala 76:26]
  reg [3:0] dataQueue_3_wstrb; // @[writeHandler.scala 76:26]
  reg  dataQueue_4_wvalid; // @[writeHandler.scala 76:26]
  reg  dataQueue_4_wlast; // @[writeHandler.scala 76:26]
  reg [31:0] dataQueue_4_wdata; // @[writeHandler.scala 76:26]
  reg [3:0] dataQueue_4_wstrb; // @[writeHandler.scala 76:26]
  reg  dataQueue_5_wvalid; // @[writeHandler.scala 76:26]
  reg  dataQueue_5_wlast; // @[writeHandler.scala 76:26]
  reg [31:0] dataQueue_5_wdata; // @[writeHandler.scala 76:26]
  reg [3:0] dataQueue_5_wstrb; // @[writeHandler.scala 76:26]
  reg  dataQueue_6_wvalid; // @[writeHandler.scala 76:26]
  reg  dataQueue_6_wlast; // @[writeHandler.scala 76:26]
  reg [31:0] dataQueue_6_wdata; // @[writeHandler.scala 76:26]
  reg [3:0] dataQueue_6_wstrb; // @[writeHandler.scala 76:26]
  reg  dataQueue_7_wvalid; // @[writeHandler.scala 76:26]
  reg  dataQueue_7_wlast; // @[writeHandler.scala 76:26]
  reg [31:0] dataQueue_7_wdata; // @[writeHandler.scala 76:26]
  reg [3:0] dataQueue_7_wstrb; // @[writeHandler.scala 76:26]
  reg [2:0] dataAllocatePointer; // @[writeHandler.scala 83:59]
  reg [2:0] dataDeallocatePointer; // @[writeHandler.scala 83:59]
  wire [31:0] _GEN_107 = 3'h0 == dataAllocatePointer ? request_alignedData[31:0] : dataQueue_0_wdata; // @[writeHandler.scala 76:26 87:{44,44}]
  wire [31:0] _GEN_108 = 3'h1 == dataAllocatePointer ? request_alignedData[31:0] : dataQueue_1_wdata; // @[writeHandler.scala 76:26 87:{44,44}]
  wire [31:0] _GEN_109 = 3'h2 == dataAllocatePointer ? request_alignedData[31:0] : dataQueue_2_wdata; // @[writeHandler.scala 76:26 87:{44,44}]
  wire [31:0] _GEN_110 = 3'h3 == dataAllocatePointer ? request_alignedData[31:0] : dataQueue_3_wdata; // @[writeHandler.scala 76:26 87:{44,44}]
  wire [31:0] _GEN_111 = 3'h4 == dataAllocatePointer ? request_alignedData[31:0] : dataQueue_4_wdata; // @[writeHandler.scala 76:26 87:{44,44}]
  wire [31:0] _GEN_112 = 3'h5 == dataAllocatePointer ? request_alignedData[31:0] : dataQueue_5_wdata; // @[writeHandler.scala 76:26 87:{44,44}]
  wire [31:0] _GEN_113 = 3'h6 == dataAllocatePointer ? request_alignedData[31:0] : dataQueue_6_wdata; // @[writeHandler.scala 76:26 87:{44,44}]
  wire [31:0] _GEN_114 = 3'h7 == dataAllocatePointer ? request_alignedData[31:0] : dataQueue_7_wdata; // @[writeHandler.scala 76:26 87:{44,44}]
  wire  _GEN_115 = 3'h0 == dataAllocatePointer ? 1'h0 : dataQueue_0_wlast; // @[writeHandler.scala 76:26 88:{44,44}]
  wire  _GEN_116 = 3'h1 == dataAllocatePointer ? 1'h0 : dataQueue_1_wlast; // @[writeHandler.scala 76:26 88:{44,44}]
  wire  _GEN_117 = 3'h2 == dataAllocatePointer ? 1'h0 : dataQueue_2_wlast; // @[writeHandler.scala 76:26 88:{44,44}]
  wire  _GEN_118 = 3'h3 == dataAllocatePointer ? 1'h0 : dataQueue_3_wlast; // @[writeHandler.scala 76:26 88:{44,44}]
  wire  _GEN_119 = 3'h4 == dataAllocatePointer ? 1'h0 : dataQueue_4_wlast; // @[writeHandler.scala 76:26 88:{44,44}]
  wire  _GEN_120 = 3'h5 == dataAllocatePointer ? 1'h0 : dataQueue_5_wlast; // @[writeHandler.scala 76:26 88:{44,44}]
  wire  _GEN_121 = 3'h6 == dataAllocatePointer ? 1'h0 : dataQueue_6_wlast; // @[writeHandler.scala 76:26 88:{44,44}]
  wire  _GEN_122 = 3'h7 == dataAllocatePointer ? 1'h0 : dataQueue_7_wlast; // @[writeHandler.scala 76:26 88:{44,44}]
  wire  _GEN_366 = 3'h0 == dataAllocatePointer; // @[writeHandler.scala 76:26 90:{45,45}]
  wire  _GEN_131 = 3'h0 == dataAllocatePointer | dataQueue_0_wvalid; // @[writeHandler.scala 76:26 90:{45,45}]
  wire  _GEN_367 = 3'h1 == dataAllocatePointer; // @[writeHandler.scala 76:26 90:{45,45}]
  wire  _GEN_132 = 3'h1 == dataAllocatePointer | dataQueue_1_wvalid; // @[writeHandler.scala 76:26 90:{45,45}]
  wire  _GEN_368 = 3'h2 == dataAllocatePointer; // @[writeHandler.scala 76:26 90:{45,45}]
  wire  _GEN_133 = 3'h2 == dataAllocatePointer | dataQueue_2_wvalid; // @[writeHandler.scala 76:26 90:{45,45}]
  wire  _GEN_369 = 3'h3 == dataAllocatePointer; // @[writeHandler.scala 76:26 90:{45,45}]
  wire  _GEN_134 = 3'h3 == dataAllocatePointer | dataQueue_3_wvalid; // @[writeHandler.scala 76:26 90:{45,45}]
  wire  _GEN_370 = 3'h4 == dataAllocatePointer; // @[writeHandler.scala 76:26 90:{45,45}]
  wire  _GEN_135 = 3'h4 == dataAllocatePointer | dataQueue_4_wvalid; // @[writeHandler.scala 76:26 90:{45,45}]
  wire  _GEN_371 = 3'h5 == dataAllocatePointer; // @[writeHandler.scala 76:26 90:{45,45}]
  wire  _GEN_136 = 3'h5 == dataAllocatePointer | dataQueue_5_wvalid; // @[writeHandler.scala 76:26 90:{45,45}]
  wire  _GEN_372 = 3'h6 == dataAllocatePointer; // @[writeHandler.scala 76:26 90:{45,45}]
  wire  _GEN_137 = 3'h6 == dataAllocatePointer | dataQueue_6_wvalid; // @[writeHandler.scala 76:26 90:{45,45}]
  wire  _GEN_373 = 3'h7 == dataAllocatePointer; // @[writeHandler.scala 76:26 90:{45,45}]
  wire  _GEN_138 = 3'h7 == dataAllocatePointer | dataQueue_7_wvalid; // @[writeHandler.scala 76:26 90:{45,45}]
  wire [2:0] _T_11 = dataAllocatePointer + 3'h1; // @[writeHandler.scala 91:36]
  wire  _GEN_374 = 3'h0 == _T_11; // @[writeHandler.scala 92:{48,48}]
  wire  _GEN_147 = 3'h0 == _T_11 | _GEN_115; // @[writeHandler.scala 92:{48,48}]
  wire  _GEN_375 = 3'h1 == _T_11; // @[writeHandler.scala 92:{48,48}]
  wire  _GEN_148 = 3'h1 == _T_11 | _GEN_116; // @[writeHandler.scala 92:{48,48}]
  wire  _GEN_376 = 3'h2 == _T_11; // @[writeHandler.scala 92:{48,48}]
  wire  _GEN_149 = 3'h2 == _T_11 | _GEN_117; // @[writeHandler.scala 92:{48,48}]
  wire  _GEN_377 = 3'h3 == _T_11; // @[writeHandler.scala 92:{48,48}]
  wire  _GEN_150 = 3'h3 == _T_11 | _GEN_118; // @[writeHandler.scala 92:{48,48}]
  wire  _GEN_378 = 3'h4 == _T_11; // @[writeHandler.scala 92:{48,48}]
  wire  _GEN_151 = 3'h4 == _T_11 | _GEN_119; // @[writeHandler.scala 92:{48,48}]
  wire  _GEN_379 = 3'h5 == _T_11; // @[writeHandler.scala 92:{48,48}]
  wire  _GEN_152 = 3'h5 == _T_11 | _GEN_120; // @[writeHandler.scala 92:{48,48}]
  wire  _GEN_380 = 3'h6 == _T_11; // @[writeHandler.scala 92:{48,48}]
  wire  _GEN_153 = 3'h6 == _T_11 | _GEN_121; // @[writeHandler.scala 92:{48,48}]
  wire  _GEN_381 = 3'h7 == _T_11; // @[writeHandler.scala 92:{48,48}]
  wire  _GEN_154 = 3'h7 == _T_11 | _GEN_122; // @[writeHandler.scala 92:{48,48}]
  wire  _GEN_163 = _GEN_374 | _GEN_131; // @[writeHandler.scala 94:{49,49}]
  wire  _GEN_164 = _GEN_375 | _GEN_132; // @[writeHandler.scala 94:{49,49}]
  wire  _GEN_165 = _GEN_376 | _GEN_133; // @[writeHandler.scala 94:{49,49}]
  wire  _GEN_166 = _GEN_377 | _GEN_134; // @[writeHandler.scala 94:{49,49}]
  wire  _GEN_167 = _GEN_378 | _GEN_135; // @[writeHandler.scala 94:{49,49}]
  wire  _GEN_168 = _GEN_379 | _GEN_136; // @[writeHandler.scala 94:{49,49}]
  wire  _GEN_169 = _GEN_380 | _GEN_137; // @[writeHandler.scala 94:{49,49}]
  wire  _GEN_170 = _GEN_381 | _GEN_138; // @[writeHandler.scala 94:{49,49}]
  wire [2:0] _dataAllocatePointer_T_1 = dataAllocatePointer + 3'h2; // @[writeHandler.scala 95:50]
  wire  _GEN_171 = _GEN_366 | dataQueue_0_wlast; // @[writeHandler.scala 76:26 97:{44,44}]
  wire  _GEN_172 = _GEN_367 | dataQueue_1_wlast; // @[writeHandler.scala 76:26 97:{44,44}]
  wire  _GEN_173 = _GEN_368 | dataQueue_2_wlast; // @[writeHandler.scala 76:26 97:{44,44}]
  wire  _GEN_174 = _GEN_369 | dataQueue_3_wlast; // @[writeHandler.scala 76:26 97:{44,44}]
  wire  _GEN_175 = _GEN_370 | dataQueue_4_wlast; // @[writeHandler.scala 76:26 97:{44,44}]
  wire  _GEN_176 = _GEN_371 | dataQueue_5_wlast; // @[writeHandler.scala 76:26 97:{44,44}]
  wire  _GEN_177 = _GEN_372 | dataQueue_6_wlast; // @[writeHandler.scala 76:26 97:{44,44}]
  wire  _GEN_178 = _GEN_373 | dataQueue_7_wlast; // @[writeHandler.scala 76:26 97:{44,44}]
  wire  _GEN_259 = _addressQueue_len_T_1 ? _GEN_163 : _GEN_131; // @[writeHandler.scala 86:47]
  wire  _GEN_260 = _addressQueue_len_T_1 ? _GEN_164 : _GEN_132; // @[writeHandler.scala 86:47]
  wire  _GEN_261 = _addressQueue_len_T_1 ? _GEN_165 : _GEN_133; // @[writeHandler.scala 86:47]
  wire  _GEN_262 = _addressQueue_len_T_1 ? _GEN_166 : _GEN_134; // @[writeHandler.scala 86:47]
  wire  _GEN_263 = _addressQueue_len_T_1 ? _GEN_167 : _GEN_135; // @[writeHandler.scala 86:47]
  wire  _GEN_264 = _addressQueue_len_T_1 ? _GEN_168 : _GEN_136; // @[writeHandler.scala 86:47]
  wire  _GEN_265 = _addressQueue_len_T_1 ? _GEN_169 : _GEN_137; // @[writeHandler.scala 86:47]
  wire  _GEN_266 = _addressQueue_len_T_1 ? _GEN_170 : _GEN_138; // @[writeHandler.scala 86:47]
  wire  _GEN_292 = request_valid ? _GEN_259 : dataQueue_0_wvalid; // @[writeHandler.scala 85:23 76:26]
  wire  _GEN_293 = request_valid ? _GEN_260 : dataQueue_1_wvalid; // @[writeHandler.scala 85:23 76:26]
  wire  _GEN_294 = request_valid ? _GEN_261 : dataQueue_2_wvalid; // @[writeHandler.scala 85:23 76:26]
  wire  _GEN_295 = request_valid ? _GEN_262 : dataQueue_3_wvalid; // @[writeHandler.scala 85:23 76:26]
  wire  _GEN_296 = request_valid ? _GEN_263 : dataQueue_4_wvalid; // @[writeHandler.scala 85:23 76:26]
  wire  _GEN_297 = request_valid ? _GEN_264 : dataQueue_5_wvalid; // @[writeHandler.scala 85:23 76:26]
  wire  _GEN_298 = request_valid ? _GEN_265 : dataQueue_6_wvalid; // @[writeHandler.scala 85:23 76:26]
  wire  _GEN_299 = request_valid ? _GEN_266 : dataQueue_7_wvalid; // @[writeHandler.scala 85:23 76:26]
  wire [2:0] _dataDeallocatePointer_T_1 = dataDeallocatePointer + 3'h1; // @[writeHandler.scala 112:52]
  wire  _dependencyCheck_free_T_23 = ~(addressQueue_0_address[31:6] == dependencyCheck_requset_address[31:6] &
    addressQueue_0_status > 2'h1 | addressQueue_1_address[31:6] == dependencyCheck_requset_address[31:6] &
    addressQueue_1_status > 2'h1 | addressQueue_2_address[31:6] == dependencyCheck_requset_address[31:6] &
    addressQueue_2_status > 2'h1 | addressQueue_3_address[31:6] == dependencyCheck_requset_address[31:6] &
    addressQueue_3_status > 2'h1); // @[writeHandler.scala 124:3]
  reg  dependencyCheck_free_REG; // @[writeHandler.scala 123:34]
  wire [31:0] _GEN_319 = 2'h1 == queryIniatePointer ? addressQueue_1_address : addressQueue_0_address; // @[writeHandler.scala 126:{14,14}]
  wire [31:0] _GEN_320 = 2'h2 == queryIniatePointer ? addressQueue_2_address : _GEN_319; // @[writeHandler.scala 126:{14,14}]
  wire  _GEN_323 = 2'h1 == queryIniatePointer ? addressQueue_1_len : addressQueue_0_len; // @[writeHandler.scala 130:{13,13}]
  wire  _GEN_324 = 2'h2 == queryIniatePointer ? addressQueue_2_len : _GEN_323; // @[writeHandler.scala 130:{13,13}]
  wire  _GEN_325 = 2'h3 == queryIniatePointer ? addressQueue_3_len : _GEN_324; // @[writeHandler.scala 130:{13,13}]
  wire [2:0] _GEN_327 = 2'h1 == queryIniatePointer ? addressQueue_1_size : addressQueue_0_size; // @[writeHandler.scala 134:{14,14}]
  wire [2:0] _GEN_328 = 2'h2 == queryIniatePointer ? addressQueue_2_size : _GEN_327; // @[writeHandler.scala 134:{14,14}]
  wire [31:0] _GEN_331 = 3'h1 == dataDeallocatePointer ? dataQueue_1_wdata : dataQueue_0_wdata; // @[writeHandler.scala 137:{13,13}]
  wire [31:0] _GEN_332 = 3'h2 == dataDeallocatePointer ? dataQueue_2_wdata : _GEN_331; // @[writeHandler.scala 137:{13,13}]
  wire [31:0] _GEN_333 = 3'h3 == dataDeallocatePointer ? dataQueue_3_wdata : _GEN_332; // @[writeHandler.scala 137:{13,13}]
  wire [31:0] _GEN_334 = 3'h4 == dataDeallocatePointer ? dataQueue_4_wdata : _GEN_333; // @[writeHandler.scala 137:{13,13}]
  wire [31:0] _GEN_335 = 3'h5 == dataDeallocatePointer ? dataQueue_5_wdata : _GEN_334; // @[writeHandler.scala 137:{13,13}]
  wire [31:0] _GEN_336 = 3'h6 == dataDeallocatePointer ? dataQueue_6_wdata : _GEN_335; // @[writeHandler.scala 137:{13,13}]
  wire  _GEN_339 = 3'h1 == dataDeallocatePointer ? dataQueue_1_wlast : dataQueue_0_wlast; // @[writeHandler.scala 138:{13,13}]
  wire  _GEN_340 = 3'h2 == dataDeallocatePointer ? dataQueue_2_wlast : _GEN_339; // @[writeHandler.scala 138:{13,13}]
  wire  _GEN_341 = 3'h3 == dataDeallocatePointer ? dataQueue_3_wlast : _GEN_340; // @[writeHandler.scala 138:{13,13}]
  wire  _GEN_342 = 3'h4 == dataDeallocatePointer ? dataQueue_4_wlast : _GEN_341; // @[writeHandler.scala 138:{13,13}]
  wire  _GEN_343 = 3'h5 == dataDeallocatePointer ? dataQueue_5_wlast : _GEN_342; // @[writeHandler.scala 138:{13,13}]
  wire  _GEN_344 = 3'h6 == dataDeallocatePointer ? dataQueue_6_wlast : _GEN_343; // @[writeHandler.scala 138:{13,13}]
  wire [3:0] _GEN_347 = 3'h1 == dataDeallocatePointer ? dataQueue_1_wstrb : dataQueue_0_wstrb; // @[writeHandler.scala 139:{13,13}]
  wire [3:0] _GEN_348 = 3'h2 == dataDeallocatePointer ? dataQueue_2_wstrb : _GEN_347; // @[writeHandler.scala 139:{13,13}]
  wire [3:0] _GEN_349 = 3'h3 == dataDeallocatePointer ? dataQueue_3_wstrb : _GEN_348; // @[writeHandler.scala 139:{13,13}]
  wire [3:0] _GEN_350 = 3'h4 == dataDeallocatePointer ? dataQueue_4_wstrb : _GEN_349; // @[writeHandler.scala 139:{13,13}]
  wire [3:0] _GEN_351 = 3'h5 == dataDeallocatePointer ? dataQueue_5_wstrb : _GEN_350; // @[writeHandler.scala 139:{13,13}]
  wire [3:0] _GEN_352 = 3'h6 == dataDeallocatePointer ? dataQueue_6_wstrb : _GEN_351; // @[writeHandler.scala 139:{13,13}]
  wire  _GEN_355 = 3'h1 == dataDeallocatePointer ? dataQueue_1_wvalid : dataQueue_0_wvalid; // @[writeHandler.scala 140:{14,14}]
  wire  _GEN_356 = 3'h2 == dataDeallocatePointer ? dataQueue_2_wvalid : _GEN_355; // @[writeHandler.scala 140:{14,14}]
  wire  _GEN_357 = 3'h3 == dataDeallocatePointer ? dataQueue_3_wvalid : _GEN_356; // @[writeHandler.scala 140:{14,14}]
  wire  _GEN_358 = 3'h4 == dataDeallocatePointer ? dataQueue_4_wvalid : _GEN_357; // @[writeHandler.scala 140:{14,14}]
  wire  _GEN_359 = 3'h5 == dataDeallocatePointer ? dataQueue_5_wvalid : _GEN_358; // @[writeHandler.scala 140:{14,14}]
  wire  _GEN_360 = 3'h6 == dataDeallocatePointer ? dataQueue_6_wvalid : _GEN_359; // @[writeHandler.scala 140:{14,14}]
  assign writeCommit_ready = _GEN_3 == 2'h0; // @[writeHandler.scala 32:62]
  assign axi_AWADDR = 2'h3 == queryIniatePointer ? addressQueue_3_address : _GEN_320; // @[writeHandler.scala 126:{14,14}]
  assign axi_AWLEN = {{7'd0}, _GEN_325}; // @[writeHandler.scala 130:13]
  assign axi_AWSIZE = 2'h3 == queryIniatePointer ? addressQueue_3_size : _GEN_328; // @[writeHandler.scala 134:{14,14}]
  assign axi_AWVALID = _GEN_83 == 2'h2; // @[writeHandler.scala 135:59]
  assign axi_WDATA = 3'h7 == dataDeallocatePointer ? dataQueue_7_wdata : _GEN_336; // @[writeHandler.scala 137:{13,13}]
  assign axi_WSTRB = 3'h7 == dataDeallocatePointer ? dataQueue_7_wstrb : _GEN_352; // @[writeHandler.scala 139:{13,13}]
  assign axi_WLAST = 3'h7 == dataDeallocatePointer ? dataQueue_7_wlast : _GEN_344; // @[writeHandler.scala 138:{13,13}]
  assign axi_WVALID = 3'h7 == dataDeallocatePointer ? dataQueue_7_wvalid : _GEN_360; // @[writeHandler.scala 140:{14,14}]
  assign axi_BREADY = _GEN_101 == 2'h3; // @[writeHandler.scala 142:57]
  assign dependencyCheck_free = dependencyCheck_free_REG; // @[writeHandler.scala 123:24]
  assign clean = addressQueue_0_status == 2'h0 & addressQueue_1_status == 2'h0 & addressQueue_2_status == 2'h0 &
    addressQueue_3_status == 2'h0; // @[writeHandler.scala 160:65]
  always @(posedge clock) begin
    if (reset) begin // @[writeHandler.scala 17:29]
      addressQueue_0_status <= 2'h0; // @[writeHandler.scala 17:29]
    end else if (axi_BVALID & axi_BREADY) begin // @[writeHandler.scala 68:34]
      if (2'h0 == deallocatePointer) begin // @[writeHandler.scala 69:44]
        addressQueue_0_status <= 2'h0; // @[writeHandler.scala 69:44]
      end else begin
        addressQueue_0_status <= _GEN_75;
      end
    end else begin
      addressQueue_0_status <= _GEN_75;
    end
    if (request_valid) begin // @[writeHandler.scala 47:23]
      if (2'h0 == queryInsertPointer) begin // @[writeHandler.scala 49:46]
        addressQueue_0_address <= request_address; // @[writeHandler.scala 49:46]
      end
    end
    if (request_valid) begin // @[writeHandler.scala 47:23]
      if (2'h0 == queryInsertPointer) begin // @[writeHandler.scala 50:42]
        addressQueue_0_len <= request_instruction[13:12] == 2'h3; // @[writeHandler.scala 50:42]
      end
    end
    if (request_valid) begin // @[writeHandler.scala 47:23]
      if (2'h0 == queryInsertPointer) begin // @[writeHandler.scala 51:43]
        if (_addressQueue_len_T_1) begin // @[writeHandler.scala 51:49]
          addressQueue_0_size <= 3'h2;
        end else begin
          addressQueue_0_size <= request_instruction[14:12];
        end
      end
    end
    if (reset) begin // @[writeHandler.scala 17:29]
      addressQueue_0_becausePeripheral <= 1'h0; // @[writeHandler.scala 17:29]
    end else if (itWasPeripheral) begin // @[writeHandler.scala 54:25]
      addressQueue_0_becausePeripheral <= _GEN_58;
    end else if (writeCommit_fired) begin // @[writeHandler.scala 34:27]
      if (2'h0 == _T_1) begin // @[writeHandler.scala 36:59]
        addressQueue_0_becausePeripheral <= 1'h0; // @[writeHandler.scala 36:59]
      end
    end
    if (reset) begin // @[writeHandler.scala 17:29]
      addressQueue_1_status <= 2'h0; // @[writeHandler.scala 17:29]
    end else if (axi_BVALID & axi_BREADY) begin // @[writeHandler.scala 68:34]
      if (2'h1 == deallocatePointer) begin // @[writeHandler.scala 69:44]
        addressQueue_1_status <= 2'h0; // @[writeHandler.scala 69:44]
      end else begin
        addressQueue_1_status <= _GEN_76;
      end
    end else begin
      addressQueue_1_status <= _GEN_76;
    end
    if (request_valid) begin // @[writeHandler.scala 47:23]
      if (2'h1 == queryInsertPointer) begin // @[writeHandler.scala 49:46]
        addressQueue_1_address <= request_address; // @[writeHandler.scala 49:46]
      end
    end
    if (request_valid) begin // @[writeHandler.scala 47:23]
      if (2'h1 == queryInsertPointer) begin // @[writeHandler.scala 50:42]
        addressQueue_1_len <= request_instruction[13:12] == 2'h3; // @[writeHandler.scala 50:42]
      end
    end
    if (request_valid) begin // @[writeHandler.scala 47:23]
      if (2'h1 == queryInsertPointer) begin // @[writeHandler.scala 51:43]
        if (_addressQueue_len_T_1) begin // @[writeHandler.scala 51:49]
          addressQueue_1_size <= 3'h2;
        end else begin
          addressQueue_1_size <= request_instruction[14:12];
        end
      end
    end
    if (reset) begin // @[writeHandler.scala 17:29]
      addressQueue_1_becausePeripheral <= 1'h0; // @[writeHandler.scala 17:29]
    end else if (itWasPeripheral) begin // @[writeHandler.scala 54:25]
      addressQueue_1_becausePeripheral <= _GEN_59;
    end else if (writeCommit_fired) begin // @[writeHandler.scala 34:27]
      if (2'h1 == _T_1) begin // @[writeHandler.scala 36:59]
        addressQueue_1_becausePeripheral <= 1'h0; // @[writeHandler.scala 36:59]
      end
    end
    if (reset) begin // @[writeHandler.scala 17:29]
      addressQueue_2_status <= 2'h0; // @[writeHandler.scala 17:29]
    end else if (axi_BVALID & axi_BREADY) begin // @[writeHandler.scala 68:34]
      if (2'h2 == deallocatePointer) begin // @[writeHandler.scala 69:44]
        addressQueue_2_status <= 2'h0; // @[writeHandler.scala 69:44]
      end else begin
        addressQueue_2_status <= _GEN_77;
      end
    end else begin
      addressQueue_2_status <= _GEN_77;
    end
    if (request_valid) begin // @[writeHandler.scala 47:23]
      if (2'h2 == queryInsertPointer) begin // @[writeHandler.scala 49:46]
        addressQueue_2_address <= request_address; // @[writeHandler.scala 49:46]
      end
    end
    if (request_valid) begin // @[writeHandler.scala 47:23]
      if (2'h2 == queryInsertPointer) begin // @[writeHandler.scala 50:42]
        addressQueue_2_len <= request_instruction[13:12] == 2'h3; // @[writeHandler.scala 50:42]
      end
    end
    if (request_valid) begin // @[writeHandler.scala 47:23]
      if (2'h2 == queryInsertPointer) begin // @[writeHandler.scala 51:43]
        if (_addressQueue_len_T_1) begin // @[writeHandler.scala 51:49]
          addressQueue_2_size <= 3'h2;
        end else begin
          addressQueue_2_size <= request_instruction[14:12];
        end
      end
    end
    if (reset) begin // @[writeHandler.scala 17:29]
      addressQueue_2_becausePeripheral <= 1'h0; // @[writeHandler.scala 17:29]
    end else if (itWasPeripheral) begin // @[writeHandler.scala 54:25]
      addressQueue_2_becausePeripheral <= _GEN_60;
    end else if (writeCommit_fired) begin // @[writeHandler.scala 34:27]
      if (2'h2 == _T_1) begin // @[writeHandler.scala 36:59]
        addressQueue_2_becausePeripheral <= 1'h0; // @[writeHandler.scala 36:59]
      end
    end
    if (reset) begin // @[writeHandler.scala 17:29]
      addressQueue_3_status <= 2'h0; // @[writeHandler.scala 17:29]
    end else if (axi_BVALID & axi_BREADY) begin // @[writeHandler.scala 68:34]
      if (2'h3 == deallocatePointer) begin // @[writeHandler.scala 69:44]
        addressQueue_3_status <= 2'h0; // @[writeHandler.scala 69:44]
      end else begin
        addressQueue_3_status <= _GEN_78;
      end
    end else begin
      addressQueue_3_status <= _GEN_78;
    end
    if (request_valid) begin // @[writeHandler.scala 47:23]
      if (2'h3 == queryInsertPointer) begin // @[writeHandler.scala 49:46]
        addressQueue_3_address <= request_address; // @[writeHandler.scala 49:46]
      end
    end
    if (request_valid) begin // @[writeHandler.scala 47:23]
      if (2'h3 == queryInsertPointer) begin // @[writeHandler.scala 50:42]
        addressQueue_3_len <= request_instruction[13:12] == 2'h3; // @[writeHandler.scala 50:42]
      end
    end
    if (request_valid) begin // @[writeHandler.scala 47:23]
      if (2'h3 == queryInsertPointer) begin // @[writeHandler.scala 51:43]
        if (_addressQueue_len_T_1) begin // @[writeHandler.scala 51:49]
          addressQueue_3_size <= 3'h2;
        end else begin
          addressQueue_3_size <= request_instruction[14:12];
        end
      end
    end
    if (reset) begin // @[writeHandler.scala 17:29]
      addressQueue_3_becausePeripheral <= 1'h0; // @[writeHandler.scala 17:29]
    end else if (itWasPeripheral) begin // @[writeHandler.scala 54:25]
      addressQueue_3_becausePeripheral <= _GEN_61;
    end else if (writeCommit_fired) begin // @[writeHandler.scala 34:27]
      if (2'h3 == _T_1) begin // @[writeHandler.scala 36:59]
        addressQueue_3_becausePeripheral <= 1'h0; // @[writeHandler.scala 36:59]
      end
    end
    if (reset) begin // @[writeHandler.scala 29:91]
      allocatePointer <= 2'h0; // @[writeHandler.scala 29:91]
    end else if (writeCommit_fired) begin // @[writeHandler.scala 34:27]
      allocatePointer <= _T_1; // @[writeHandler.scala 37:21]
    end
    if (reset) begin // @[writeHandler.scala 29:91]
      queryInsertPointer <= 2'h0; // @[writeHandler.scala 29:91]
    end else if (itWasPeripheral) begin // @[writeHandler.scala 54:25]
      queryInsertPointer <= _queryInsertPointer_T_1; // @[writeHandler.scala 57:24]
    end else if (request_valid) begin // @[writeHandler.scala 47:23]
      queryInsertPointer <= _queryInsertPointer_T_1; // @[writeHandler.scala 52:24]
    end
    if (reset) begin // @[writeHandler.scala 29:91]
      queryIniatePointer <= 2'h0; // @[writeHandler.scala 29:91]
    end else if (_GEN_83 == 2'h0 & _GEN_87) begin // @[writeHandler.scala 64:124]
      queryIniatePointer <= _queryIniatePointer_T_1; // @[writeHandler.scala 65:24]
    end else if (axi_AWVALID & axi_AWREADY) begin // @[writeHandler.scala 60:36]
      queryIniatePointer <= _queryIniatePointer_T_1; // @[writeHandler.scala 62:24]
    end
    if (reset) begin // @[writeHandler.scala 29:91]
      deallocatePointer <= 2'h0; // @[writeHandler.scala 29:91]
    end else if (_GEN_101 == 2'h0 & _GEN_105) begin // @[writeHandler.scala 72:122]
      deallocatePointer <= _deallocatePointer_T_1; // @[writeHandler.scala 73:23]
    end else if (axi_BVALID & axi_BREADY) begin // @[writeHandler.scala 68:34]
      deallocatePointer <= _deallocatePointer_T_1; // @[writeHandler.scala 70:23]
    end
    if (reset) begin // @[writeHandler.scala 76:26]
      dataQueue_0_wvalid <= 1'h0; // @[writeHandler.scala 76:26]
    end else if (axi_WVALID & axi_WREADY) begin // @[writeHandler.scala 110:34]
      if (3'h0 == dataDeallocatePointer) begin // @[writeHandler.scala 111:45]
        dataQueue_0_wvalid <= 1'h0; // @[writeHandler.scala 111:45]
      end else begin
        dataQueue_0_wvalid <= _GEN_292;
      end
    end else begin
      dataQueue_0_wvalid <= _GEN_292;
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        dataQueue_0_wlast <= _GEN_147;
      end else begin
        dataQueue_0_wlast <= _GEN_171;
      end
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        if (3'h0 == _T_11) begin // @[writeHandler.scala 91:48]
          dataQueue_0_wdata <= request_alignedData[63:32]; // @[writeHandler.scala 91:48]
        end else begin
          dataQueue_0_wdata <= _GEN_107;
        end
      end else if (|request_mask[3:0]) begin // @[writeHandler.scala 100:36]
        dataQueue_0_wdata <= _GEN_107;
      end else if (3'h0 == dataAllocatePointer) begin // @[writeHandler.scala 104:46]
        dataQueue_0_wdata <= request_alignedData[63:32]; // @[writeHandler.scala 104:46]
      end
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        if (3'h0 == _T_11) begin // @[writeHandler.scala 93:48]
          dataQueue_0_wstrb <= 4'hf; // @[writeHandler.scala 93:48]
        end else if (3'h0 == dataAllocatePointer) begin // @[writeHandler.scala 89:44]
          dataQueue_0_wstrb <= 4'hf; // @[writeHandler.scala 89:44]
        end
      end else if (|request_mask[3:0]) begin // @[writeHandler.scala 100:36]
        if (3'h0 == dataAllocatePointer) begin // @[writeHandler.scala 102:46]
          dataQueue_0_wstrb <= request_mask[3:0]; // @[writeHandler.scala 102:46]
        end
      end else if (3'h0 == dataAllocatePointer) begin // @[writeHandler.scala 105:46]
        dataQueue_0_wstrb <= request_mask[7:4]; // @[writeHandler.scala 105:46]
      end
    end
    if (reset) begin // @[writeHandler.scala 76:26]
      dataQueue_1_wvalid <= 1'h0; // @[writeHandler.scala 76:26]
    end else if (axi_WVALID & axi_WREADY) begin // @[writeHandler.scala 110:34]
      if (3'h1 == dataDeallocatePointer) begin // @[writeHandler.scala 111:45]
        dataQueue_1_wvalid <= 1'h0; // @[writeHandler.scala 111:45]
      end else begin
        dataQueue_1_wvalid <= _GEN_293;
      end
    end else begin
      dataQueue_1_wvalid <= _GEN_293;
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        dataQueue_1_wlast <= _GEN_148;
      end else begin
        dataQueue_1_wlast <= _GEN_172;
      end
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        if (3'h1 == _T_11) begin // @[writeHandler.scala 91:48]
          dataQueue_1_wdata <= request_alignedData[63:32]; // @[writeHandler.scala 91:48]
        end else begin
          dataQueue_1_wdata <= _GEN_108;
        end
      end else if (|request_mask[3:0]) begin // @[writeHandler.scala 100:36]
        dataQueue_1_wdata <= _GEN_108;
      end else if (3'h1 == dataAllocatePointer) begin // @[writeHandler.scala 104:46]
        dataQueue_1_wdata <= request_alignedData[63:32]; // @[writeHandler.scala 104:46]
      end
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        if (3'h1 == _T_11) begin // @[writeHandler.scala 93:48]
          dataQueue_1_wstrb <= 4'hf; // @[writeHandler.scala 93:48]
        end else if (3'h1 == dataAllocatePointer) begin // @[writeHandler.scala 89:44]
          dataQueue_1_wstrb <= 4'hf; // @[writeHandler.scala 89:44]
        end
      end else if (|request_mask[3:0]) begin // @[writeHandler.scala 100:36]
        if (3'h1 == dataAllocatePointer) begin // @[writeHandler.scala 102:46]
          dataQueue_1_wstrb <= request_mask[3:0]; // @[writeHandler.scala 102:46]
        end
      end else if (3'h1 == dataAllocatePointer) begin // @[writeHandler.scala 105:46]
        dataQueue_1_wstrb <= request_mask[7:4]; // @[writeHandler.scala 105:46]
      end
    end
    if (reset) begin // @[writeHandler.scala 76:26]
      dataQueue_2_wvalid <= 1'h0; // @[writeHandler.scala 76:26]
    end else if (axi_WVALID & axi_WREADY) begin // @[writeHandler.scala 110:34]
      if (3'h2 == dataDeallocatePointer) begin // @[writeHandler.scala 111:45]
        dataQueue_2_wvalid <= 1'h0; // @[writeHandler.scala 111:45]
      end else begin
        dataQueue_2_wvalid <= _GEN_294;
      end
    end else begin
      dataQueue_2_wvalid <= _GEN_294;
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        dataQueue_2_wlast <= _GEN_149;
      end else begin
        dataQueue_2_wlast <= _GEN_173;
      end
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        if (3'h2 == _T_11) begin // @[writeHandler.scala 91:48]
          dataQueue_2_wdata <= request_alignedData[63:32]; // @[writeHandler.scala 91:48]
        end else begin
          dataQueue_2_wdata <= _GEN_109;
        end
      end else if (|request_mask[3:0]) begin // @[writeHandler.scala 100:36]
        dataQueue_2_wdata <= _GEN_109;
      end else if (3'h2 == dataAllocatePointer) begin // @[writeHandler.scala 104:46]
        dataQueue_2_wdata <= request_alignedData[63:32]; // @[writeHandler.scala 104:46]
      end
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        if (3'h2 == _T_11) begin // @[writeHandler.scala 93:48]
          dataQueue_2_wstrb <= 4'hf; // @[writeHandler.scala 93:48]
        end else if (3'h2 == dataAllocatePointer) begin // @[writeHandler.scala 89:44]
          dataQueue_2_wstrb <= 4'hf; // @[writeHandler.scala 89:44]
        end
      end else if (|request_mask[3:0]) begin // @[writeHandler.scala 100:36]
        if (3'h2 == dataAllocatePointer) begin // @[writeHandler.scala 102:46]
          dataQueue_2_wstrb <= request_mask[3:0]; // @[writeHandler.scala 102:46]
        end
      end else if (3'h2 == dataAllocatePointer) begin // @[writeHandler.scala 105:46]
        dataQueue_2_wstrb <= request_mask[7:4]; // @[writeHandler.scala 105:46]
      end
    end
    if (reset) begin // @[writeHandler.scala 76:26]
      dataQueue_3_wvalid <= 1'h0; // @[writeHandler.scala 76:26]
    end else if (axi_WVALID & axi_WREADY) begin // @[writeHandler.scala 110:34]
      if (3'h3 == dataDeallocatePointer) begin // @[writeHandler.scala 111:45]
        dataQueue_3_wvalid <= 1'h0; // @[writeHandler.scala 111:45]
      end else begin
        dataQueue_3_wvalid <= _GEN_295;
      end
    end else begin
      dataQueue_3_wvalid <= _GEN_295;
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        dataQueue_3_wlast <= _GEN_150;
      end else begin
        dataQueue_3_wlast <= _GEN_174;
      end
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        if (3'h3 == _T_11) begin // @[writeHandler.scala 91:48]
          dataQueue_3_wdata <= request_alignedData[63:32]; // @[writeHandler.scala 91:48]
        end else begin
          dataQueue_3_wdata <= _GEN_110;
        end
      end else if (|request_mask[3:0]) begin // @[writeHandler.scala 100:36]
        dataQueue_3_wdata <= _GEN_110;
      end else if (3'h3 == dataAllocatePointer) begin // @[writeHandler.scala 104:46]
        dataQueue_3_wdata <= request_alignedData[63:32]; // @[writeHandler.scala 104:46]
      end
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        if (3'h3 == _T_11) begin // @[writeHandler.scala 93:48]
          dataQueue_3_wstrb <= 4'hf; // @[writeHandler.scala 93:48]
        end else if (3'h3 == dataAllocatePointer) begin // @[writeHandler.scala 89:44]
          dataQueue_3_wstrb <= 4'hf; // @[writeHandler.scala 89:44]
        end
      end else if (|request_mask[3:0]) begin // @[writeHandler.scala 100:36]
        if (3'h3 == dataAllocatePointer) begin // @[writeHandler.scala 102:46]
          dataQueue_3_wstrb <= request_mask[3:0]; // @[writeHandler.scala 102:46]
        end
      end else if (3'h3 == dataAllocatePointer) begin // @[writeHandler.scala 105:46]
        dataQueue_3_wstrb <= request_mask[7:4]; // @[writeHandler.scala 105:46]
      end
    end
    if (reset) begin // @[writeHandler.scala 76:26]
      dataQueue_4_wvalid <= 1'h0; // @[writeHandler.scala 76:26]
    end else if (axi_WVALID & axi_WREADY) begin // @[writeHandler.scala 110:34]
      if (3'h4 == dataDeallocatePointer) begin // @[writeHandler.scala 111:45]
        dataQueue_4_wvalid <= 1'h0; // @[writeHandler.scala 111:45]
      end else begin
        dataQueue_4_wvalid <= _GEN_296;
      end
    end else begin
      dataQueue_4_wvalid <= _GEN_296;
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        dataQueue_4_wlast <= _GEN_151;
      end else begin
        dataQueue_4_wlast <= _GEN_175;
      end
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        if (3'h4 == _T_11) begin // @[writeHandler.scala 91:48]
          dataQueue_4_wdata <= request_alignedData[63:32]; // @[writeHandler.scala 91:48]
        end else begin
          dataQueue_4_wdata <= _GEN_111;
        end
      end else if (|request_mask[3:0]) begin // @[writeHandler.scala 100:36]
        dataQueue_4_wdata <= _GEN_111;
      end else if (3'h4 == dataAllocatePointer) begin // @[writeHandler.scala 104:46]
        dataQueue_4_wdata <= request_alignedData[63:32]; // @[writeHandler.scala 104:46]
      end
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        if (3'h4 == _T_11) begin // @[writeHandler.scala 93:48]
          dataQueue_4_wstrb <= 4'hf; // @[writeHandler.scala 93:48]
        end else if (3'h4 == dataAllocatePointer) begin // @[writeHandler.scala 89:44]
          dataQueue_4_wstrb <= 4'hf; // @[writeHandler.scala 89:44]
        end
      end else if (|request_mask[3:0]) begin // @[writeHandler.scala 100:36]
        if (3'h4 == dataAllocatePointer) begin // @[writeHandler.scala 102:46]
          dataQueue_4_wstrb <= request_mask[3:0]; // @[writeHandler.scala 102:46]
        end
      end else if (3'h4 == dataAllocatePointer) begin // @[writeHandler.scala 105:46]
        dataQueue_4_wstrb <= request_mask[7:4]; // @[writeHandler.scala 105:46]
      end
    end
    if (reset) begin // @[writeHandler.scala 76:26]
      dataQueue_5_wvalid <= 1'h0; // @[writeHandler.scala 76:26]
    end else if (axi_WVALID & axi_WREADY) begin // @[writeHandler.scala 110:34]
      if (3'h5 == dataDeallocatePointer) begin // @[writeHandler.scala 111:45]
        dataQueue_5_wvalid <= 1'h0; // @[writeHandler.scala 111:45]
      end else begin
        dataQueue_5_wvalid <= _GEN_297;
      end
    end else begin
      dataQueue_5_wvalid <= _GEN_297;
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        dataQueue_5_wlast <= _GEN_152;
      end else begin
        dataQueue_5_wlast <= _GEN_176;
      end
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        if (3'h5 == _T_11) begin // @[writeHandler.scala 91:48]
          dataQueue_5_wdata <= request_alignedData[63:32]; // @[writeHandler.scala 91:48]
        end else begin
          dataQueue_5_wdata <= _GEN_112;
        end
      end else if (|request_mask[3:0]) begin // @[writeHandler.scala 100:36]
        dataQueue_5_wdata <= _GEN_112;
      end else if (3'h5 == dataAllocatePointer) begin // @[writeHandler.scala 104:46]
        dataQueue_5_wdata <= request_alignedData[63:32]; // @[writeHandler.scala 104:46]
      end
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        if (3'h5 == _T_11) begin // @[writeHandler.scala 93:48]
          dataQueue_5_wstrb <= 4'hf; // @[writeHandler.scala 93:48]
        end else if (3'h5 == dataAllocatePointer) begin // @[writeHandler.scala 89:44]
          dataQueue_5_wstrb <= 4'hf; // @[writeHandler.scala 89:44]
        end
      end else if (|request_mask[3:0]) begin // @[writeHandler.scala 100:36]
        if (3'h5 == dataAllocatePointer) begin // @[writeHandler.scala 102:46]
          dataQueue_5_wstrb <= request_mask[3:0]; // @[writeHandler.scala 102:46]
        end
      end else if (3'h5 == dataAllocatePointer) begin // @[writeHandler.scala 105:46]
        dataQueue_5_wstrb <= request_mask[7:4]; // @[writeHandler.scala 105:46]
      end
    end
    if (reset) begin // @[writeHandler.scala 76:26]
      dataQueue_6_wvalid <= 1'h0; // @[writeHandler.scala 76:26]
    end else if (axi_WVALID & axi_WREADY) begin // @[writeHandler.scala 110:34]
      if (3'h6 == dataDeallocatePointer) begin // @[writeHandler.scala 111:45]
        dataQueue_6_wvalid <= 1'h0; // @[writeHandler.scala 111:45]
      end else begin
        dataQueue_6_wvalid <= _GEN_298;
      end
    end else begin
      dataQueue_6_wvalid <= _GEN_298;
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        dataQueue_6_wlast <= _GEN_153;
      end else begin
        dataQueue_6_wlast <= _GEN_177;
      end
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        if (3'h6 == _T_11) begin // @[writeHandler.scala 91:48]
          dataQueue_6_wdata <= request_alignedData[63:32]; // @[writeHandler.scala 91:48]
        end else begin
          dataQueue_6_wdata <= _GEN_113;
        end
      end else if (|request_mask[3:0]) begin // @[writeHandler.scala 100:36]
        dataQueue_6_wdata <= _GEN_113;
      end else if (3'h6 == dataAllocatePointer) begin // @[writeHandler.scala 104:46]
        dataQueue_6_wdata <= request_alignedData[63:32]; // @[writeHandler.scala 104:46]
      end
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        if (3'h6 == _T_11) begin // @[writeHandler.scala 93:48]
          dataQueue_6_wstrb <= 4'hf; // @[writeHandler.scala 93:48]
        end else if (3'h6 == dataAllocatePointer) begin // @[writeHandler.scala 89:44]
          dataQueue_6_wstrb <= 4'hf; // @[writeHandler.scala 89:44]
        end
      end else if (|request_mask[3:0]) begin // @[writeHandler.scala 100:36]
        if (3'h6 == dataAllocatePointer) begin // @[writeHandler.scala 102:46]
          dataQueue_6_wstrb <= request_mask[3:0]; // @[writeHandler.scala 102:46]
        end
      end else if (3'h6 == dataAllocatePointer) begin // @[writeHandler.scala 105:46]
        dataQueue_6_wstrb <= request_mask[7:4]; // @[writeHandler.scala 105:46]
      end
    end
    if (reset) begin // @[writeHandler.scala 76:26]
      dataQueue_7_wvalid <= 1'h0; // @[writeHandler.scala 76:26]
    end else if (axi_WVALID & axi_WREADY) begin // @[writeHandler.scala 110:34]
      if (3'h7 == dataDeallocatePointer) begin // @[writeHandler.scala 111:45]
        dataQueue_7_wvalid <= 1'h0; // @[writeHandler.scala 111:45]
      end else begin
        dataQueue_7_wvalid <= _GEN_299;
      end
    end else begin
      dataQueue_7_wvalid <= _GEN_299;
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        dataQueue_7_wlast <= _GEN_154;
      end else begin
        dataQueue_7_wlast <= _GEN_178;
      end
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        if (3'h7 == _T_11) begin // @[writeHandler.scala 91:48]
          dataQueue_7_wdata <= request_alignedData[63:32]; // @[writeHandler.scala 91:48]
        end else begin
          dataQueue_7_wdata <= _GEN_114;
        end
      end else if (|request_mask[3:0]) begin // @[writeHandler.scala 100:36]
        dataQueue_7_wdata <= _GEN_114;
      end else if (3'h7 == dataAllocatePointer) begin // @[writeHandler.scala 104:46]
        dataQueue_7_wdata <= request_alignedData[63:32]; // @[writeHandler.scala 104:46]
      end
    end
    if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        if (3'h7 == _T_11) begin // @[writeHandler.scala 93:48]
          dataQueue_7_wstrb <= 4'hf; // @[writeHandler.scala 93:48]
        end else if (3'h7 == dataAllocatePointer) begin // @[writeHandler.scala 89:44]
          dataQueue_7_wstrb <= 4'hf; // @[writeHandler.scala 89:44]
        end
      end else if (|request_mask[3:0]) begin // @[writeHandler.scala 100:36]
        if (3'h7 == dataAllocatePointer) begin // @[writeHandler.scala 102:46]
          dataQueue_7_wstrb <= request_mask[3:0]; // @[writeHandler.scala 102:46]
        end
      end else if (3'h7 == dataAllocatePointer) begin // @[writeHandler.scala 105:46]
        dataQueue_7_wstrb <= request_mask[7:4]; // @[writeHandler.scala 105:46]
      end
    end
    if (reset) begin // @[writeHandler.scala 83:59]
      dataAllocatePointer <= 3'h0; // @[writeHandler.scala 83:59]
    end else if (request_valid) begin // @[writeHandler.scala 85:23]
      if (_addressQueue_len_T_1) begin // @[writeHandler.scala 86:47]
        dataAllocatePointer <= _dataAllocatePointer_T_1; // @[writeHandler.scala 95:27]
      end else begin
        dataAllocatePointer <= _T_11; // @[writeHandler.scala 99:27]
      end
    end
    if (reset) begin // @[writeHandler.scala 83:59]
      dataDeallocatePointer <= 3'h0; // @[writeHandler.scala 83:59]
    end else if (axi_WVALID & axi_WREADY) begin // @[writeHandler.scala 110:34]
      dataDeallocatePointer <= _dataDeallocatePointer_T_1; // @[writeHandler.scala 112:27]
    end
    if (reset) begin // @[writeHandler.scala 123:34]
      dependencyCheck_free_REG <= 1'h0; // @[writeHandler.scala 123:34]
    end else begin
      dependencyCheck_free_REG <= dependencyCheck_requset_valid & _dependencyCheck_free_T_23; // @[writeHandler.scala 123:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addressQueue_0_status = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  addressQueue_0_address = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  addressQueue_0_len = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  addressQueue_0_size = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  addressQueue_0_becausePeripheral = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  addressQueue_1_status = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  addressQueue_1_address = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  addressQueue_1_len = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  addressQueue_1_size = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  addressQueue_1_becausePeripheral = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  addressQueue_2_status = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  addressQueue_2_address = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  addressQueue_2_len = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  addressQueue_2_size = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  addressQueue_2_becausePeripheral = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  addressQueue_3_status = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  addressQueue_3_address = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  addressQueue_3_len = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  addressQueue_3_size = _RAND_18[2:0];
  _RAND_19 = {1{`RANDOM}};
  addressQueue_3_becausePeripheral = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  allocatePointer = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  queryInsertPointer = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  queryIniatePointer = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  deallocatePointer = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  dataQueue_0_wvalid = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  dataQueue_0_wlast = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  dataQueue_0_wdata = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  dataQueue_0_wstrb = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  dataQueue_1_wvalid = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  dataQueue_1_wlast = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  dataQueue_1_wdata = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  dataQueue_1_wstrb = _RAND_31[3:0];
  _RAND_32 = {1{`RANDOM}};
  dataQueue_2_wvalid = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  dataQueue_2_wlast = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  dataQueue_2_wdata = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  dataQueue_2_wstrb = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  dataQueue_3_wvalid = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  dataQueue_3_wlast = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  dataQueue_3_wdata = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  dataQueue_3_wstrb = _RAND_39[3:0];
  _RAND_40 = {1{`RANDOM}};
  dataQueue_4_wvalid = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  dataQueue_4_wlast = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  dataQueue_4_wdata = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  dataQueue_4_wstrb = _RAND_43[3:0];
  _RAND_44 = {1{`RANDOM}};
  dataQueue_5_wvalid = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  dataQueue_5_wlast = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  dataQueue_5_wdata = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  dataQueue_5_wstrb = _RAND_47[3:0];
  _RAND_48 = {1{`RANDOM}};
  dataQueue_6_wvalid = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  dataQueue_6_wlast = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  dataQueue_6_wdata = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  dataQueue_6_wstrb = _RAND_51[3:0];
  _RAND_52 = {1{`RANDOM}};
  dataQueue_7_wvalid = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  dataQueue_7_wlast = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  dataQueue_7_wdata = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  dataQueue_7_wstrb = _RAND_55[3:0];
  _RAND_56 = {1{`RANDOM}};
  dataAllocatePointer = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  dataDeallocatePointer = _RAND_57[2:0];
  _RAND_58 = {1{`RANDOM}};
  dependencyCheck_free_REG = _RAND_58[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module core_Anon_1(
  input         clock,
  input         reset,
  output [31:0] peripheral_AWADDR,
  output [7:0]  peripheral_AWLEN,
  output [2:0]  peripheral_AWSIZE,
  output        peripheral_AWVALID,
  input         peripheral_AWREADY,
  output [31:0] peripheral_WDATA,
  output [3:0]  peripheral_WSTRB,
  output        peripheral_WLAST,
  output        peripheral_WVALID,
  input         peripheral_WREADY,
  input         peripheral_BVALID,
  output        peripheral_BREADY,
  output [31:0] peripheral_ARADDR,
  output [7:0]  peripheral_ARLEN,
  output [2:0]  peripheral_ARSIZE,
  output        peripheral_ARVALID,
  input         peripheral_ARREADY,
  input  [31:0] peripheral_RDATA,
  input         peripheral_RLAST,
  input         peripheral_RVALID,
  output        peripheral_RREADY,
  input         branchOps_valid,
  input  [3:0]  branchOps_branchMask,
  input         branchOps_passed,
  input         writeDataIn_valid,
  input  [63:0] writeDataIn_data,
  output        responseOut_valid,
  output [5:0]  responseOut_prfDest,
  output [3:0]  responseOut_robAddr,
  output [63:0] responseOut_result,
  output [31:0] responseOut_instruction,
  input         request_valid,
  input  [31:0] request_address,
  input  [31:0] request_instruction,
  input  [3:0]  request_branchMask,
  input  [3:0]  request_robAddr,
  input  [5:0]  request_prfDest,
  output [31:0] dPort_AWADDR,
  output [7:0]  dPort_AWLEN,
  output [2:0]  dPort_AWSIZE,
  output        dPort_AWVALID,
  input         dPort_AWREADY,
  output [31:0] dPort_WDATA,
  output [3:0]  dPort_WSTRB,
  output        dPort_WLAST,
  output        dPort_WVALID,
  input         dPort_WREADY,
  input         dPort_BVALID,
  output        dPort_BREADY,
  output [31:0] dPort_ARADDR,
  output        dPort_ARVALID,
  input         dPort_ARREADY,
  input  [31:0] dPort_RDATA,
  input         dPort_RLAST,
  input         dPort_RVALID,
  output        dPort_RREADY,
  output        writeCommit_ready,
  input         writeCommit_fired,
  output        canAllocate,
  input         initiateFence,
  output        fenceInstructions_ready,
  input         fenceInstructions_fired
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
`endif // RANDOMIZE_REG_INIT
  wire  scheduler_clock; // @[memAccess.scala 13:25]
  wire  scheduler_reset; // @[memAccess.scala 13:25]
  wire  scheduler_toCache_queryWithData_query_valid; // @[memAccess.scala 13:25]
  wire [31:0] scheduler_toCache_queryWithData_query_address; // @[memAccess.scala 13:25]
  wire [31:0] scheduler_toCache_queryWithData_query_instruction; // @[memAccess.scala 13:25]
  wire [3:0] scheduler_toCache_queryWithData_query_branchMask; // @[memAccess.scala 13:25]
  wire [3:0] scheduler_toCache_queryWithData_query_robAddr; // @[memAccess.scala 13:25]
  wire [5:0] scheduler_toCache_queryWithData_query_prfDest; // @[memAccess.scala 13:25]
  wire [63:0] scheduler_toCache_queryWithData_data; // @[memAccess.scala 13:25]
  wire  scheduler_toCache_replaying; // @[memAccess.scala 13:25]
  wire  scheduler_storeCommit_ready; // @[memAccess.scala 13:25]
  wire  scheduler_storeCommit_fired; // @[memAccess.scala 13:25]
  wire  scheduler_replaying; // @[memAccess.scala 13:25]
  wire  scheduler_cacheStalled; // @[memAccess.scala 13:25]
  wire  scheduler_replayQueue_query_valid; // @[memAccess.scala 13:25]
  wire [31:0] scheduler_replayQueue_query_address; // @[memAccess.scala 13:25]
  wire [31:0] scheduler_replayQueue_query_instruction; // @[memAccess.scala 13:25]
  wire [3:0] scheduler_replayQueue_query_branchMask; // @[memAccess.scala 13:25]
  wire [3:0] scheduler_replayQueue_query_robAddr; // @[memAccess.scala 13:25]
  wire [5:0] scheduler_replayQueue_query_prfDest; // @[memAccess.scala 13:25]
  wire [63:0] scheduler_replayQueue_data; // @[memAccess.scala 13:25]
  wire  scheduler_branchOps_valid; // @[memAccess.scala 13:25]
  wire [3:0] scheduler_branchOps_branchMask; // @[memAccess.scala 13:25]
  wire  scheduler_branchOps_passed; // @[memAccess.scala 13:25]
  wire  scheduler_peripheral_ready; // @[memAccess.scala 13:25]
  wire  scheduler_peripheral_bits_valid; // @[memAccess.scala 13:25]
  wire [31:0] scheduler_peripheral_bits_address; // @[memAccess.scala 13:25]
  wire [31:0] scheduler_peripheral_bits_instruction; // @[memAccess.scala 13:25]
  wire [3:0] scheduler_peripheral_bits_branchMask; // @[memAccess.scala 13:25]
  wire [3:0] scheduler_peripheral_bits_robAddr; // @[memAccess.scala 13:25]
  wire [5:0] scheduler_peripheral_bits_prfDest; // @[memAccess.scala 13:25]
  wire  scheduler_newInstruction_valid; // @[memAccess.scala 13:25]
  wire [31:0] scheduler_newInstruction_address; // @[memAccess.scala 13:25]
  wire [31:0] scheduler_newInstruction_instruction; // @[memAccess.scala 13:25]
  wire [3:0] scheduler_newInstruction_branchMask; // @[memAccess.scala 13:25]
  wire [3:0] scheduler_newInstruction_robAddr; // @[memAccess.scala 13:25]
  wire [5:0] scheduler_newInstruction_prfDest; // @[memAccess.scala 13:25]
  wire  scheduler_canAllocate; // @[memAccess.scala 13:25]
  wire  scheduler_clean; // @[memAccess.scala 13:25]
  wire  peripheralHandler_clock; // @[memAccess.scala 19:33]
  wire  peripheralHandler_reset; // @[memAccess.scala 19:33]
  wire  peripheralHandler_request_valid; // @[memAccess.scala 19:33]
  wire [31:0] peripheralHandler_request_address; // @[memAccess.scala 19:33]
  wire [31:0] peripheralHandler_request_instruction; // @[memAccess.scala 19:33]
  wire [3:0] peripheralHandler_request_branchMask; // @[memAccess.scala 19:33]
  wire [3:0] peripheralHandler_request_robAddr; // @[memAccess.scala 19:33]
  wire [5:0] peripheralHandler_request_prfDest; // @[memAccess.scala 19:33]
  wire  peripheralHandler_finishedRequest_valid; // @[memAccess.scala 19:33]
  wire [31:0] peripheralHandler_finishedRequest_address; // @[memAccess.scala 19:33]
  wire [31:0] peripheralHandler_finishedRequest_instruction; // @[memAccess.scala 19:33]
  wire [3:0] peripheralHandler_finishedRequest_robAddr; // @[memAccess.scala 19:33]
  wire [5:0] peripheralHandler_finishedRequest_prfDest; // @[memAccess.scala 19:33]
  wire  peripheralHandler_ready; // @[memAccess.scala 19:33]
  wire  peripheralHandler_branchOps_valid; // @[memAccess.scala 19:33]
  wire [3:0] peripheralHandler_branchOps_branchMask; // @[memAccess.scala 19:33]
  wire  peripheralHandler_branchOps_passed; // @[memAccess.scala 19:33]
  wire [31:0] peripheralHandler_axi_AWADDR; // @[memAccess.scala 19:33]
  wire [7:0] peripheralHandler_axi_AWLEN; // @[memAccess.scala 19:33]
  wire [2:0] peripheralHandler_axi_AWSIZE; // @[memAccess.scala 19:33]
  wire  peripheralHandler_axi_AWVALID; // @[memAccess.scala 19:33]
  wire  peripheralHandler_axi_AWREADY; // @[memAccess.scala 19:33]
  wire [31:0] peripheralHandler_axi_WDATA; // @[memAccess.scala 19:33]
  wire [3:0] peripheralHandler_axi_WSTRB; // @[memAccess.scala 19:33]
  wire  peripheralHandler_axi_WLAST; // @[memAccess.scala 19:33]
  wire  peripheralHandler_axi_WVALID; // @[memAccess.scala 19:33]
  wire  peripheralHandler_axi_WREADY; // @[memAccess.scala 19:33]
  wire  peripheralHandler_axi_BVALID; // @[memAccess.scala 19:33]
  wire  peripheralHandler_axi_BREADY; // @[memAccess.scala 19:33]
  wire [31:0] peripheralHandler_axi_ARADDR; // @[memAccess.scala 19:33]
  wire [7:0] peripheralHandler_axi_ARLEN; // @[memAccess.scala 19:33]
  wire [2:0] peripheralHandler_axi_ARSIZE; // @[memAccess.scala 19:33]
  wire  peripheralHandler_axi_ARVALID; // @[memAccess.scala 19:33]
  wire  peripheralHandler_axi_ARREADY; // @[memAccess.scala 19:33]
  wire [31:0] peripheralHandler_axi_RDATA; // @[memAccess.scala 19:33]
  wire  peripheralHandler_axi_RLAST; // @[memAccess.scala 19:33]
  wire  peripheralHandler_axi_RVALID; // @[memAccess.scala 19:33]
  wire  peripheralHandler_axi_RREADY; // @[memAccess.scala 19:33]
  wire  peripheralHandler_readFinished_ready; // @[memAccess.scala 19:33]
  wire  peripheralHandler_readFinished_fired; // @[memAccess.scala 19:33]
  wire [63:0] peripheralHandler_readDataOut; // @[memAccess.scala 19:33]
  wire  peripheralHandler_writeIn_valid; // @[memAccess.scala 19:33]
  wire [63:0] peripheralHandler_writeIn_data; // @[memAccess.scala 19:33]
  wire  cache_clock; // @[memAccess.scala 46:21]
  wire  cache_reset; // @[memAccess.scala 46:21]
  wire [31:0] cache_readAddress; // @[memAccess.scala 46:21]
  wire [63:0] cache_readOut_0_data; // @[memAccess.scala 46:21]
  wire [19:0] cache_readOut_0_tag; // @[memAccess.scala 46:21]
  wire  cache_readOut_0_valid; // @[memAccess.scala 46:21]
  wire [63:0] cache_readOut_1_data; // @[memAccess.scala 46:21]
  wire [19:0] cache_readOut_1_tag; // @[memAccess.scala 46:21]
  wire  cache_readOut_1_valid; // @[memAccess.scala 46:21]
  wire  cache_writePorts_0_enable; // @[memAccess.scala 46:21]
  wire [31:0] cache_writePorts_0_cacheAddress; // @[memAccess.scala 46:21]
  wire [63:0] cache_writePorts_0_data; // @[memAccess.scala 46:21]
  wire  cache_writePorts_1_enable; // @[memAccess.scala 46:21]
  wire [31:0] cache_writePorts_1_cacheAddress; // @[memAccess.scala 46:21]
  wire [63:0] cache_writePorts_1_data; // @[memAccess.scala 46:21]
  wire  cache_invalidateSet_valid; // @[memAccess.scala 46:21]
  wire [5:0] cache_invalidateSet_cacheIndex; // @[memAccess.scala 46:21]
  wire  cache_invalidateSet_invalidateVector_0; // @[memAccess.scala 46:21]
  wire  cache_invalidateSet_invalidateVector_1; // @[memAccess.scala 46:21]
  wire  cache_cacheFillDone_valid; // @[memAccess.scala 46:21]
  wire [5:0] cache_cacheFillDone_cacheIndex; // @[memAccess.scala 46:21]
  wire  cache_cacheFillDone_validateVector_0; // @[memAccess.scala 46:21]
  wire  cache_cacheFillDone_validateVector_1; // @[memAccess.scala 46:21]
  wire [19:0] cache_cacheFillDone_tag; // @[memAccess.scala 46:21]
  wire  missHandler_clock; // @[memAccess.scala 128:27]
  wire  missHandler_reset; // @[memAccess.scala 128:27]
  wire  missHandler_replayOut_query_valid; // @[memAccess.scala 128:27]
  wire [31:0] missHandler_replayOut_query_address; // @[memAccess.scala 128:27]
  wire [31:0] missHandler_replayOut_query_instruction; // @[memAccess.scala 128:27]
  wire [3:0] missHandler_replayOut_query_branchMask; // @[memAccess.scala 128:27]
  wire [3:0] missHandler_replayOut_query_robAddr; // @[memAccess.scala 128:27]
  wire [5:0] missHandler_replayOut_query_prfDest; // @[memAccess.scala 128:27]
  wire [63:0] missHandler_replayOut_data; // @[memAccess.scala 128:27]
  wire  missHandler_replayingQuries; // @[memAccess.scala 128:27]
  wire  missHandler_branchOps_valid; // @[memAccess.scala 128:27]
  wire [3:0] missHandler_branchOps_branchMask; // @[memAccess.scala 128:27]
  wire  missHandler_branchOps_passed; // @[memAccess.scala 128:27]
  wire  missHandler_cachePipelineEmpty; // @[memAccess.scala 128:27]
  wire  missHandler_missedRequest_query_valid; // @[memAccess.scala 128:27]
  wire [31:0] missHandler_missedRequest_query_address; // @[memAccess.scala 128:27]
  wire [31:0] missHandler_missedRequest_query_instruction; // @[memAccess.scala 128:27]
  wire [3:0] missHandler_missedRequest_query_branchMask; // @[memAccess.scala 128:27]
  wire [3:0] missHandler_missedRequest_query_robAddr; // @[memAccess.scala 128:27]
  wire [5:0] missHandler_missedRequest_query_prfDest; // @[memAccess.scala 128:27]
  wire [63:0] missHandler_missedRequest_data; // @[memAccess.scala 128:27]
  wire  missHandler_pushToCache_ready; // @[memAccess.scala 128:27]
  wire  missHandler_pushToCache_fired; // @[memAccess.scala 128:27]
  wire [63:0] missHandler_pushToCache_cacheWriteOut_data; // @[memAccess.scala 128:27]
  wire [8:0] missHandler_pushToCache_cacheWriteOut_address; // @[memAccess.scala 128:27]
  wire [1:0] missHandler_pushToCache_cacheWriteOut_setSelVector; // @[memAccess.scala 128:27]
  wire [31:0] missHandler_axi_ARADDR; // @[memAccess.scala 128:27]
  wire  missHandler_axi_ARVALID; // @[memAccess.scala 128:27]
  wire  missHandler_axi_ARREADY; // @[memAccess.scala 128:27]
  wire [31:0] missHandler_axi_RDATA; // @[memAccess.scala 128:27]
  wire  missHandler_axi_RLAST; // @[memAccess.scala 128:27]
  wire  missHandler_axi_RVALID; // @[memAccess.scala 128:27]
  wire  missHandler_axi_RREADY; // @[memAccess.scala 128:27]
  wire  missHandler_dependencyCheck_requset_valid; // @[memAccess.scala 128:27]
  wire [31:0] missHandler_dependencyCheck_requset_address; // @[memAccess.scala 128:27]
  wire  missHandler_dependencyCheck_free; // @[memAccess.scala 128:27]
  wire  missHandler_rlastToCache; // @[memAccess.scala 128:27]
  wire [1:0] missHandler_setInvalidateVector; // @[memAccess.scala 128:27]
  wire [1:0] missHandler_setFillStatus; // @[memAccess.scala 128:27]
  wire  missHandler_handlerBusy; // @[memAccess.scala 128:27]
  wire  missHandler_handlerSaturated; // @[memAccess.scala 128:27]
  wire  missHandler_clean; // @[memAccess.scala 128:27]
  wire  missHandler_nonSaturatedReplay; // @[memAccess.scala 128:27]
  wire  writeHandler_clock; // @[memAccess.scala 378:28]
  wire  writeHandler_reset; // @[memAccess.scala 378:28]
  wire  writeHandler_itWasPeripheral; // @[memAccess.scala 378:28]
  wire  writeHandler_writeCommit_ready; // @[memAccess.scala 378:28]
  wire  writeHandler_writeCommit_fired; // @[memAccess.scala 378:28]
  wire [31:0] writeHandler_axi_AWADDR; // @[memAccess.scala 378:28]
  wire [7:0] writeHandler_axi_AWLEN; // @[memAccess.scala 378:28]
  wire [2:0] writeHandler_axi_AWSIZE; // @[memAccess.scala 378:28]
  wire  writeHandler_axi_AWVALID; // @[memAccess.scala 378:28]
  wire  writeHandler_axi_AWREADY; // @[memAccess.scala 378:28]
  wire [31:0] writeHandler_axi_WDATA; // @[memAccess.scala 378:28]
  wire [3:0] writeHandler_axi_WSTRB; // @[memAccess.scala 378:28]
  wire  writeHandler_axi_WLAST; // @[memAccess.scala 378:28]
  wire  writeHandler_axi_WVALID; // @[memAccess.scala 378:28]
  wire  writeHandler_axi_WREADY; // @[memAccess.scala 378:28]
  wire  writeHandler_axi_BVALID; // @[memAccess.scala 378:28]
  wire  writeHandler_axi_BREADY; // @[memAccess.scala 378:28]
  wire  writeHandler_request_valid; // @[memAccess.scala 378:28]
  wire [31:0] writeHandler_request_address; // @[memAccess.scala 378:28]
  wire [31:0] writeHandler_request_instruction; // @[memAccess.scala 378:28]
  wire [63:0] writeHandler_request_alignedData; // @[memAccess.scala 378:28]
  wire [7:0] writeHandler_request_mask; // @[memAccess.scala 378:28]
  wire  writeHandler_dependencyCheck_requset_valid; // @[memAccess.scala 378:28]
  wire [31:0] writeHandler_dependencyCheck_requset_address; // @[memAccess.scala 378:28]
  wire  writeHandler_dependencyCheck_free; // @[memAccess.scala 378:28]
  wire  writeHandler_clean; // @[memAccess.scala 378:28]
  reg  reservation_valid; // @[memAccess.scala 33:28]
  reg [31:0] reservation_address; // @[memAccess.scala 33:28]
  reg  reservation64_valid; // @[memAccess.scala 38:30]
  reg [31:0] reservation64_address; // @[memAccess.scala 38:30]
  reg  dataQueue_0_valid; // @[memAccess.scala 52:26]
  reg [63:0] dataQueue_0_data; // @[memAccess.scala 52:26]
  reg  dataQueue_1_valid; // @[memAccess.scala 52:26]
  reg [63:0] dataQueue_1_data; // @[memAccess.scala 52:26]
  reg  dataQueue_2_valid; // @[memAccess.scala 52:26]
  reg [63:0] dataQueue_2_data; // @[memAccess.scala 52:26]
  reg  dataQueue_3_valid; // @[memAccess.scala 52:26]
  reg [63:0] dataQueue_3_data; // @[memAccess.scala 52:26]
  reg [63:0] dataToCache; // @[memAccess.scala 57:24]
  reg  servicing_query_valid; // @[memAccess.scala 61:26]
  reg [31:0] servicing_query_address; // @[memAccess.scala 61:26]
  reg [31:0] servicing_query_instruction; // @[memAccess.scala 61:26]
  reg [3:0] servicing_query_branchMask; // @[memAccess.scala 61:26]
  reg [3:0] servicing_query_robAddr; // @[memAccess.scala 61:26]
  reg [5:0] servicing_query_prfDest; // @[memAccess.scala 61:26]
  reg [63:0] servicing_data; // @[memAccess.scala 61:26]
  wire  _T_2 = scheduler_toCache_queryWithData_query_address >= 32'h80000000; // @[configuration.scala 41:44]
  wire  _GEN_2 = ~_T_2 ? 1'h0 : scheduler_toCache_queryWithData_query_valid; // @[memAccess.scala 63:19 73:68 74:27]
  reg  cacheLookUp_query_valid; // @[memAccess.scala 79:28]
  reg [31:0] cacheLookUp_query_address; // @[memAccess.scala 79:28]
  reg [31:0] cacheLookUp_query_instruction; // @[memAccess.scala 79:28]
  reg [3:0] cacheLookUp_query_branchMask; // @[memAccess.scala 79:28]
  reg [3:0] cacheLookUp_query_robAddr; // @[memAccess.scala 79:28]
  reg [5:0] cacheLookUp_query_prfDest; // @[memAccess.scala 79:28]
  reg [63:0] cacheLookUp_write_dataByteAligned; // @[memAccess.scala 79:28]
  reg [7:0] cacheLookUp_write_aligedMask; // @[memAccess.scala 79:28]
  reg [1:0] cacheLookUp_hitVector; // @[memAccess.scala 79:28]
  reg [1:0] cacheLookUp_setFillVector; // @[memAccess.scala 79:28]
  reg [63:0] cacheLookUp_cacheDouble; // @[memAccess.scala 79:28]
  wire  _cacheLookUp_hitVector_T_2 = cache_readOut_0_valid & cache_readOut_0_tag == servicing_query_address[31:12]; // @[memAccess.scala 90:63]
  wire  _cacheLookUp_hitVector_T_5 = cache_readOut_1_valid & cache_readOut_1_tag == servicing_query_address[31:12]; // @[memAccess.scala 90:63]
  wire [5:0] _GEN_5 = 3'h1 == servicing_query_address[2:0] ? 6'h8 : 6'h0; // @[memAccess.scala 92:{55,55}]
  wire [5:0] _GEN_6 = 3'h2 == servicing_query_address[2:0] ? 6'h10 : _GEN_5; // @[memAccess.scala 92:{55,55}]
  wire [5:0] _GEN_7 = 3'h3 == servicing_query_address[2:0] ? 6'h18 : _GEN_6; // @[memAccess.scala 92:{55,55}]
  wire [5:0] _GEN_8 = 3'h4 == servicing_query_address[2:0] ? 6'h20 : _GEN_7; // @[memAccess.scala 92:{55,55}]
  wire [5:0] _GEN_9 = 3'h5 == servicing_query_address[2:0] ? 6'h28 : _GEN_8; // @[memAccess.scala 92:{55,55}]
  wire [5:0] _GEN_10 = 3'h6 == servicing_query_address[2:0] ? 6'h30 : _GEN_9; // @[memAccess.scala 92:{55,55}]
  wire [5:0] _GEN_11 = 3'h7 == servicing_query_address[2:0] ? 6'h38 : _GEN_10; // @[memAccess.scala 92:{55,55}]
  wire [126:0] _GEN_97 = {{63'd0}, servicing_data}; // @[memAccess.scala 92:55]
  wire [126:0] _cacheLookUp_write_dataByteAligned_T_1 = _GEN_97 << _GEN_11; // @[memAccess.scala 92:55]
  wire [7:0] _GEN_13 = 2'h1 == servicing_query_instruction[13:12] ? 8'h3 : 8'h1; // @[memAccess.scala 93:{103,103}]
  wire [7:0] _GEN_14 = 2'h2 == servicing_query_instruction[13:12] ? 8'hf : _GEN_13; // @[memAccess.scala 93:{103,103}]
  wire [7:0] _GEN_15 = 2'h3 == servicing_query_instruction[13:12] ? 8'hff : _GEN_14; // @[memAccess.scala 93:{103,103}]
  wire [14:0] _GEN_99 = {{7'd0}, _GEN_15}; // @[memAccess.scala 93:103]
  wire [14:0] _cacheLookUp_write_aligedMask_T_2 = _GEN_99 << servicing_query_address[2:0]; // @[memAccess.scala 93:103]
  reg  memoryResponse_query_valid; // @[memAccess.scala 96:31]
  reg [31:0] memoryResponse_query_address; // @[memAccess.scala 96:31]
  reg [31:0] memoryResponse_query_instruction; // @[memAccess.scala 96:31]
  reg [3:0] memoryResponse_query_robAddr; // @[memAccess.scala 96:31]
  reg [5:0] memoryResponse_query_prfDest; // @[memAccess.scala 96:31]
  reg [63:0] memoryResponse_write_dataByteAligned; // @[memAccess.scala 96:31]
  reg [7:0] memoryResponse_write_aligedMask; // @[memAccess.scala 96:31]
  reg  memoryResponse_hit; // @[memAccess.scala 96:31]
  reg [1:0] memoryResponse_hitVector; // @[memAccess.scala 96:31]
  reg [63:0] memoryResponse_readData; // @[memAccess.scala 96:31]
  reg  memoryResponse_invalidate_valid; // @[memAccess.scala 96:31]
  reg [5:0] memoryResponse_invalidate_cacheIndex; // @[memAccess.scala 96:31]
  reg  memoryResponse_invalidate_invalidateVector_0; // @[memAccess.scala 96:31]
  reg  memoryResponse_invalidate_invalidateVector_1; // @[memAccess.scala 96:31]
  reg  memoryResponse_cacheSetFill_valid; // @[memAccess.scala 96:31]
  reg [5:0] memoryResponse_cacheSetFill_cacheIndex; // @[memAccess.scala 96:31]
  reg  memoryResponse_cacheSetFill_validateVector_0; // @[memAccess.scala 96:31]
  reg  memoryResponse_cacheSetFill_validateVector_1; // @[memAccess.scala 96:31]
  reg [19:0] memoryResponse_cacheSetFill_tag; // @[memAccess.scala 96:31]
  reg  memoryResponse_filling; // @[memAccess.scala 96:31]
  wire  _memoryResponseWriteDataByteAligned_semaphore64_T = reservation64_address == cacheLookUp_query_address; // @[memAccess.scala 213:58]
  wire [63:0] _memoryResponseWriteDataByteAligned_semaphore64_T_2 = reservation64_valid & reservation64_address ==
    cacheLookUp_query_address ? cacheLookUp_write_dataByteAligned : cacheLookUp_cacheDouble; // @[memAccess.scala 213:12]
  wire [63:0] _GEN_74 = cacheLookUp_query_instruction[27] ? _memoryResponseWriteDataByteAligned_semaphore64_T_2 :
    cacheLookUp_cacheDouble; // @[memAccess.scala 219:{25,25}]
  wire  _memoryResponseWriteDataByteAligned_atomic64_T_20 = cacheLookUp_cacheDouble < cacheLookUp_write_dataByteAligned; // @[memAccess.scala 227:37]
  wire [63:0] _memoryResponseWriteDataByteAligned_atomic64_T_21 = cacheLookUp_cacheDouble <
    cacheLookUp_write_dataByteAligned ? cacheLookUp_write_dataByteAligned : cacheLookUp_cacheDouble; // @[memAccess.scala 227:12]
  wire [63:0] _memoryResponseWriteDataByteAligned_atomic64_T_19 = _memoryResponseWriteDataByteAligned_atomic64_T_20 ?
    cacheLookUp_cacheDouble : cacheLookUp_write_dataByteAligned; // @[memAccess.scala 226:12]
  wire  _memoryResponseWriteDataByteAligned_atomic64_T_16 = $signed(cacheLookUp_cacheDouble) < $signed(
    cacheLookUp_write_dataByteAligned); // @[memAccess.scala 225:44]
  wire [63:0] _memoryResponseWriteDataByteAligned_atomic64_T_17 = $signed(cacheLookUp_cacheDouble) < $signed(
    cacheLookUp_write_dataByteAligned) ? cacheLookUp_write_dataByteAligned : cacheLookUp_cacheDouble; // @[memAccess.scala 225:12]
  wire [63:0] _memoryResponseWriteDataByteAligned_atomic64_T_13 = _memoryResponseWriteDataByteAligned_atomic64_T_16 ?
    cacheLookUp_cacheDouble : cacheLookUp_write_dataByteAligned; // @[memAccess.scala 224:12]
  wire [63:0] _memoryResponseWriteDataByteAligned_atomic64_T_9 = cacheLookUp_cacheDouble &
    cacheLookUp_write_dataByteAligned; // @[memAccess.scala 223:33]
  wire [63:0] _memoryResponseWriteDataByteAligned_atomic64_T_8 = cacheLookUp_cacheDouble |
    cacheLookUp_write_dataByteAligned; // @[memAccess.scala 222:33]
  wire [63:0] _memoryResponseWriteDataByteAligned_atomic64_T_7 = cacheLookUp_cacheDouble ^
    cacheLookUp_write_dataByteAligned; // @[memAccess.scala 221:33]
  wire [63:0] _memoryResponseWriteDataByteAligned_atomic64_T_5 = cacheLookUp_cacheDouble +
    cacheLookUp_write_dataByteAligned; // @[memAccess.scala 220:114]
  wire [63:0] _memoryResponseWriteDataByteAligned_atomic64_T_6 = cacheLookUp_query_instruction[27] ?
    cacheLookUp_write_dataByteAligned : _memoryResponseWriteDataByteAligned_atomic64_T_5; // @[memAccess.scala 220:12]
  wire [63:0] _GEN_76 = 3'h1 == cacheLookUp_query_instruction[31:29] ? _memoryResponseWriteDataByteAligned_atomic64_T_7
     : _memoryResponseWriteDataByteAligned_atomic64_T_6; // @[memAccess.scala 219:{25,25}]
  wire [63:0] _GEN_77 = 3'h2 == cacheLookUp_query_instruction[31:29] ? _memoryResponseWriteDataByteAligned_atomic64_T_8
     : _GEN_76; // @[memAccess.scala 219:{25,25}]
  wire [63:0] _GEN_78 = 3'h3 == cacheLookUp_query_instruction[31:29] ? _memoryResponseWriteDataByteAligned_atomic64_T_9
     : _GEN_77; // @[memAccess.scala 219:{25,25}]
  wire [63:0] _GEN_79 = 3'h4 == cacheLookUp_query_instruction[31:29] ? _memoryResponseWriteDataByteAligned_atomic64_T_13
     : _GEN_78; // @[memAccess.scala 219:{25,25}]
  wire [63:0] _GEN_80 = 3'h5 == cacheLookUp_query_instruction[31:29] ? _memoryResponseWriteDataByteAligned_atomic64_T_17
     : _GEN_79; // @[memAccess.scala 219:{25,25}]
  wire [63:0] _GEN_81 = 3'h6 == cacheLookUp_query_instruction[31:29] ? _memoryResponseWriteDataByteAligned_atomic64_T_19
     : _GEN_80; // @[memAccess.scala 219:{25,25}]
  wire [63:0] _GEN_82 = 3'h7 == cacheLookUp_query_instruction[31:29] ? _memoryResponseWriteDataByteAligned_atomic64_T_21
     : _GEN_81; // @[memAccess.scala 219:{25,25}]
  wire [63:0] memoryResponseWriteDataByteAligned_atomic64 = cacheLookUp_query_instruction[28] ? _GEN_74 : _GEN_82; // @[memAccess.scala 219:25]
  wire  _memoryResponseWriteDataByteAligned_semaphore32High_T_1 = reservation_address == cacheLookUp_query_address; // @[memAccess.scala 236:30]
  wire  _memoryResponseWriteDataByteAligned_semaphore32High_T_2 = reservation_valid &
    _memoryResponseWriteDataByteAligned_semaphore32High_T_1; // @[memAccess.scala 235:31]
  wire [31:0] _memoryResponseWriteDataByteAligned_semaphore32High_T_5 = reservation_valid &
    _memoryResponseWriteDataByteAligned_semaphore32High_T_1 ? cacheLookUp_write_dataByteAligned[63:32] :
    cacheLookUp_cacheDouble[63:32]; // @[memAccess.scala 235:12]
  wire [31:0] _GEN_84 = cacheLookUp_query_instruction[27] ? _memoryResponseWriteDataByteAligned_semaphore32High_T_5 :
    cacheLookUp_cacheDouble[63:32]; // @[memAccess.scala 250:{28,28}]
  wire [31:0] _memoryResponseWriteDataByteAligned_semaphore32Low_T_5 =
    _memoryResponseWriteDataByteAligned_semaphore32High_T_2 ? cacheLookUp_write_dataByteAligned[31:0] :
    cacheLookUp_cacheDouble[31:0]; // @[memAccess.scala 244:12]
  wire [31:0] _GEN_86 = cacheLookUp_query_instruction[27] ? _memoryResponseWriteDataByteAligned_semaphore32Low_T_5 :
    cacheLookUp_cacheDouble[31:0]; // @[memAccess.scala 250:{28,28}]
  wire [31:0] memoryResponseWriteDataByteAligned_semaphore32 = cacheLookUp_query_address[2] ? _GEN_84 : _GEN_86; // @[memAccess.scala 250:28]
  wire [31:0] memoryResponseWriteDataByteAligned_atomic32Src1 = cacheLookUp_query_address[2] ? cacheLookUp_cacheDouble[
    63:32] : cacheLookUp_cacheDouble[31:0]; // @[memAccess.scala 230:29]
  wire [31:0] memoryResponseWriteDataByteAligned_atomic32Src2 = cacheLookUp_query_address[2] ?
    cacheLookUp_write_dataByteAligned[63:32] : cacheLookUp_write_dataByteAligned[31:0]; // @[memAccess.scala 231:29]
  wire  _memoryResponseWriteDataByteAligned_atomic32_T_20 = memoryResponseWriteDataByteAligned_atomic32Src1 <
    memoryResponseWriteDataByteAligned_atomic32Src2; // @[memAccess.scala 260:26]
  wire [31:0] _memoryResponseWriteDataByteAligned_atomic32_T_21 = memoryResponseWriteDataByteAligned_atomic32Src1 <
    memoryResponseWriteDataByteAligned_atomic32Src2 ? memoryResponseWriteDataByteAligned_atomic32Src2 :
    memoryResponseWriteDataByteAligned_atomic32Src1; // @[memAccess.scala 260:12]
  wire [31:0] _memoryResponseWriteDataByteAligned_atomic32_T_19 = _memoryResponseWriteDataByteAligned_atomic32_T_20 ?
    memoryResponseWriteDataByteAligned_atomic32Src1 : memoryResponseWriteDataByteAligned_atomic32Src2; // @[memAccess.scala 259:12]
  wire [31:0] _memoryResponseWriteDataByteAligned_atomic32_T_14 = cacheLookUp_query_address[2] ? cacheLookUp_cacheDouble
    [63:32] : cacheLookUp_cacheDouble[31:0]; // @[memAccess.scala 258:26]
  wire [31:0] _memoryResponseWriteDataByteAligned_atomic32_T_15 = cacheLookUp_query_address[2] ?
    cacheLookUp_write_dataByteAligned[63:32] : cacheLookUp_write_dataByteAligned[31:0]; // @[memAccess.scala 258:48]
  wire  _memoryResponseWriteDataByteAligned_atomic32_T_16 = $signed(_memoryResponseWriteDataByteAligned_atomic32_T_14)
     < $signed(_memoryResponseWriteDataByteAligned_atomic32_T_15); // @[memAccess.scala 258:33]
  wire [31:0] _memoryResponseWriteDataByteAligned_atomic32_T_17 = $signed(
    _memoryResponseWriteDataByteAligned_atomic32_T_14) < $signed(_memoryResponseWriteDataByteAligned_atomic32_T_15) ?
    memoryResponseWriteDataByteAligned_atomic32Src2 : memoryResponseWriteDataByteAligned_atomic32Src1; // @[memAccess.scala 258:12]
  wire [31:0] _memoryResponseWriteDataByteAligned_atomic32_T_13 = _memoryResponseWriteDataByteAligned_atomic32_T_16 ?
    memoryResponseWriteDataByteAligned_atomic32Src1 : memoryResponseWriteDataByteAligned_atomic32Src2; // @[memAccess.scala 257:12]
  wire [31:0] _memoryResponseWriteDataByteAligned_atomic32_T_9 = memoryResponseWriteDataByteAligned_atomic32Src1 &
    memoryResponseWriteDataByteAligned_atomic32Src2; // @[memAccess.scala 256:22]
  wire [31:0] _memoryResponseWriteDataByteAligned_atomic32_T_8 = memoryResponseWriteDataByteAligned_atomic32Src1 |
    memoryResponseWriteDataByteAligned_atomic32Src2; // @[memAccess.scala 255:22]
  wire [31:0] _memoryResponseWriteDataByteAligned_atomic32_T_7 = memoryResponseWriteDataByteAligned_atomic32Src1 ^
    memoryResponseWriteDataByteAligned_atomic32Src2; // @[memAccess.scala 254:22]
  wire [31:0] _memoryResponseWriteDataByteAligned_atomic32_T_5 = memoryResponseWriteDataByteAligned_atomic32Src1 +
    memoryResponseWriteDataByteAligned_atomic32Src2; // @[memAccess.scala 253:82]
  wire [31:0] _memoryResponseWriteDataByteAligned_atomic32_T_6 = cacheLookUp_query_instruction[27] ?
    memoryResponseWriteDataByteAligned_atomic32Src2 : _memoryResponseWriteDataByteAligned_atomic32_T_5; // @[memAccess.scala 253:12]
  wire [31:0] _GEN_88 = 3'h1 == cacheLookUp_query_instruction[31:29] ? _memoryResponseWriteDataByteAligned_atomic32_T_7
     : _memoryResponseWriteDataByteAligned_atomic32_T_6; // @[memAccess.scala 252:{25,25}]
  wire [31:0] _GEN_89 = 3'h2 == cacheLookUp_query_instruction[31:29] ? _memoryResponseWriteDataByteAligned_atomic32_T_8
     : _GEN_88; // @[memAccess.scala 252:{25,25}]
  wire [31:0] _GEN_90 = 3'h3 == cacheLookUp_query_instruction[31:29] ? _memoryResponseWriteDataByteAligned_atomic32_T_9
     : _GEN_89; // @[memAccess.scala 252:{25,25}]
  wire [31:0] _GEN_91 = 3'h4 == cacheLookUp_query_instruction[31:29] ? _memoryResponseWriteDataByteAligned_atomic32_T_13
     : _GEN_90; // @[memAccess.scala 252:{25,25}]
  wire [31:0] _GEN_92 = 3'h5 == cacheLookUp_query_instruction[31:29] ? _memoryResponseWriteDataByteAligned_atomic32_T_17
     : _GEN_91; // @[memAccess.scala 252:{25,25}]
  wire [31:0] _GEN_93 = 3'h6 == cacheLookUp_query_instruction[31:29] ? _memoryResponseWriteDataByteAligned_atomic32_T_19
     : _GEN_92; // @[memAccess.scala 252:{25,25}]
  wire [31:0] _GEN_94 = 3'h7 == cacheLookUp_query_instruction[31:29] ? _memoryResponseWriteDataByteAligned_atomic32_T_21
     : _GEN_93; // @[memAccess.scala 252:{25,25}]
  wire [31:0] memoryResponseWriteDataByteAligned_atomic32 = cacheLookUp_query_instruction[28] ?
    memoryResponseWriteDataByteAligned_semaphore32 : _GEN_94; // @[memAccess.scala 252:25]
  wire [63:0] _memoryResponseWriteDataByteAligned_postAtomic32_T_3 = {memoryResponseWriteDataByteAligned_atomic32,
    cacheLookUp_cacheDouble[31:0]}; // @[Cat.scala 33:92]
  wire [63:0] _memoryResponseWriteDataByteAligned_postAtomic32_T_1 = {cacheLookUp_cacheDouble[63:32],
    memoryResponseWriteDataByteAligned_atomic32}; // @[Cat.scala 33:92]
  wire [63:0] _GEN_96 = cacheLookUp_query_address[2] ? _memoryResponseWriteDataByteAligned_postAtomic32_T_3 :
    _memoryResponseWriteDataByteAligned_postAtomic32_T_1; // @[memAccess.scala 264:{23,23}]
  wire [63:0] _memoryResponseWriteDataByteAligned_storeData_T_30 = cacheLookUp_write_aligedMask[7] ?
    cacheLookUp_write_dataByteAligned : cacheLookUp_cacheDouble; // @[memAccess.scala 209:51]
  wire [63:0] _memoryResponseWriteDataByteAligned_storeData_T_26 = cacheLookUp_write_aligedMask[6] ?
    cacheLookUp_write_dataByteAligned : cacheLookUp_cacheDouble; // @[memAccess.scala 209:51]
  wire [63:0] _memoryResponseWriteDataByteAligned_storeData_T_22 = cacheLookUp_write_aligedMask[5] ?
    cacheLookUp_write_dataByteAligned : cacheLookUp_cacheDouble; // @[memAccess.scala 209:51]
  wire [63:0] _memoryResponseWriteDataByteAligned_storeData_T_18 = cacheLookUp_write_aligedMask[4] ?
    cacheLookUp_write_dataByteAligned : cacheLookUp_cacheDouble; // @[memAccess.scala 209:51]
  wire [63:0] _memoryResponseWriteDataByteAligned_storeData_T_14 = cacheLookUp_write_aligedMask[3] ?
    cacheLookUp_write_dataByteAligned : cacheLookUp_cacheDouble; // @[memAccess.scala 209:51]
  wire [63:0] _memoryResponseWriteDataByteAligned_storeData_T_10 = cacheLookUp_write_aligedMask[2] ?
    cacheLookUp_write_dataByteAligned : cacheLookUp_cacheDouble; // @[memAccess.scala 209:51]
  wire [63:0] _memoryResponseWriteDataByteAligned_storeData_T_6 = cacheLookUp_write_aligedMask[1] ?
    cacheLookUp_write_dataByteAligned : cacheLookUp_cacheDouble; // @[memAccess.scala 209:51]
  wire [63:0] _memoryResponseWriteDataByteAligned_storeData_T_2 = cacheLookUp_write_aligedMask[0] ?
    cacheLookUp_write_dataByteAligned : cacheLookUp_cacheDouble; // @[memAccess.scala 209:51]
  wire [63:0] memoryResponseWriteDataByteAligned_storeData = {_memoryResponseWriteDataByteAligned_storeData_T_30[63:56],
    _memoryResponseWriteDataByteAligned_storeData_T_26[55:48],_memoryResponseWriteDataByteAligned_storeData_T_22[47:40],
    _memoryResponseWriteDataByteAligned_storeData_T_18[39:32],_memoryResponseWriteDataByteAligned_storeData_T_14[31:24],
    _memoryResponseWriteDataByteAligned_storeData_T_10[23:16],_memoryResponseWriteDataByteAligned_storeData_T_6[15:8],
    _memoryResponseWriteDataByteAligned_storeData_T_2[7:0]}; // @[Cat.scala 33:92]
  wire  _cacheLookUp_cacheDouble_T_10 = cacheLookUp_query_valid & cacheLookUp_query_instruction[5] &
    cacheLookUp_query_address[31:3] == servicing_query_address[31:3]; // @[memAccess.scala 123:75]
  wire  _cacheLookUp_cacheDouble_T_13 = memoryResponse_query_valid & memoryResponse_query_instruction[5]; // @[memAccess.scala 124:35]
  wire  _cacheLookUp_cacheDouble_T_17 = memoryResponse_query_valid & memoryResponse_query_instruction[5] &
    memoryResponse_query_address[31:3] == servicing_query_address[31:3]; // @[memAccess.scala 124:81]
  wire [5:0] _GEN_17 = 3'h1 == cacheLookUp_query_address[2:0] ? 6'h8 : 6'h0; // @[memAccess.scala 132:{55,55}]
  wire [5:0] _GEN_18 = 3'h2 == cacheLookUp_query_address[2:0] ? 6'h10 : _GEN_17; // @[memAccess.scala 132:{55,55}]
  wire [5:0] _GEN_19 = 3'h3 == cacheLookUp_query_address[2:0] ? 6'h18 : _GEN_18; // @[memAccess.scala 132:{55,55}]
  wire [5:0] _GEN_20 = 3'h4 == cacheLookUp_query_address[2:0] ? 6'h20 : _GEN_19; // @[memAccess.scala 132:{55,55}]
  wire [5:0] _GEN_21 = 3'h5 == cacheLookUp_query_address[2:0] ? 6'h28 : _GEN_20; // @[memAccess.scala 132:{55,55}]
  wire [5:0] _GEN_22 = 3'h6 == cacheLookUp_query_address[2:0] ? 6'h30 : _GEN_21; // @[memAccess.scala 132:{55,55}]
  wire [5:0] _GEN_23 = 3'h7 == cacheLookUp_query_address[2:0] ? 6'h38 : _GEN_22; // @[memAccess.scala 132:{55,55}]
  wire  _missHandler_missedRequest_T_1 = ~missHandler_handlerBusy; // @[memAccess.scala 135:12]
  wire  _missHandler_missedRequest_T_4 = |cacheLookUp_hitVector; // @[memAccess.scala 136:92]
  wire  _GEN_24 = cacheLookUp_query_instruction[6:2] == 5'h8 | |cacheLookUp_hitVector ? 1'h0 : cacheLookUp_query_valid; // @[memAccess.scala 136:119 133:25 136:97]
  wire  _GEN_26 = _missHandler_missedRequest_T_4 ? 1'h0 : cacheLookUp_query_valid; // @[memAccess.scala 133:25 141:{41,63}]
  wire  _GEN_27 = cacheLookUp_query_address[31:6] != missHandler_dependencyCheck_requset_address[31:6] ? _GEN_24 :
    _GEN_26; // @[memAccess.scala 137:143]
  wire  _GEN_28 = ~missHandler_handlerBusy ? _GEN_24 : _GEN_27; // @[memAccess.scala 135:38]
  wire  _GEN_29 = ~missHandler_handlerSaturated ? _GEN_28 : cacheLookUp_query_valid; // @[memAccess.scala 133:25 134:41]
  wire  _missHandler_missedRequest_T_18 = missHandler_dependencyCheck_requset_address[31:6] == cacheLookUp_query_address
    [31:6] & _missHandler_missedRequest_T_4; // @[memAccess.scala 146:135]
  wire  _GEN_30 = _missHandler_missedRequest_T_18 ? 1'h0 : _GEN_29; // @[memAccess.scala 148:{31,9}]
  wire  _GEN_31 = missHandler_handlerBusy ? _GEN_30 : _GEN_29; // @[memAccess.scala 144:35]
  wire [3:0] _missHandler_missedRequest_T_19 = branchOps_branchMask & cacheLookUp_query_branchMask; // @[memAccess.scala 150:51]
  wire  _missHandler_missedRequest_T_21 = branchOps_valid & |_missHandler_missedRequest_T_19; // @[memAccess.scala 150:26]
  wire [3:0] _missHandler_missedRequest_request_query_branchMask_T = branchOps_branchMask ^ cacheLookUp_query_branchMask
    ; // @[memAccess.scala 151:81]
  wire [3:0] _GEN_32 = branchOps_passed ? _missHandler_missedRequest_request_query_branchMask_T :
    cacheLookUp_query_branchMask; // @[memAccess.scala 131:19 151:{30,57}]
  wire  _GEN_33 = branchOps_passed & _GEN_31; // @[memAccess.scala 151:30 152:40]
  wire  _missHandler_cachePipelineEmpty_T_1 = scheduler_toCache_queryWithData_query_valid | servicing_query_valid |
    cacheLookUp_query_valid; // @[memAccess.scala 162:14]
  wire  _GEN_37 = 3'h1 == cacheLookUp_query_address[2:0] ? cacheLookUp_cacheDouble[15] : cacheLookUp_cacheDouble[7]; // @[memAccess.scala 186:{24,24}]
  wire  _GEN_38 = 3'h2 == cacheLookUp_query_address[2:0] ? cacheLookUp_cacheDouble[23] : _GEN_37; // @[memAccess.scala 186:{24,24}]
  wire  _GEN_39 = 3'h3 == cacheLookUp_query_address[2:0] ? cacheLookUp_cacheDouble[31] : _GEN_38; // @[memAccess.scala 186:{24,24}]
  wire  _GEN_40 = 3'h4 == cacheLookUp_query_address[2:0] ? cacheLookUp_cacheDouble[39] : _GEN_39; // @[memAccess.scala 186:{24,24}]
  wire  _GEN_41 = 3'h5 == cacheLookUp_query_address[2:0] ? cacheLookUp_cacheDouble[47] : _GEN_40; // @[memAccess.scala 186:{24,24}]
  wire  _GEN_42 = 3'h6 == cacheLookUp_query_address[2:0] ? cacheLookUp_cacheDouble[55] : _GEN_41; // @[memAccess.scala 186:{24,24}]
  wire  _GEN_43 = 3'h7 == cacheLookUp_query_address[2:0] ? cacheLookUp_cacheDouble[63] : _GEN_42; // @[memAccess.scala 186:{24,24}]
  wire  _GEN_45 = 2'h1 == cacheLookUp_query_address[2:1] ? cacheLookUp_cacheDouble[31] : cacheLookUp_cacheDouble[15]; // @[memAccess.scala 186:{24,24}]
  wire  _GEN_46 = 2'h2 == cacheLookUp_query_address[2:1] ? cacheLookUp_cacheDouble[47] : _GEN_45; // @[memAccess.scala 186:{24,24}]
  wire  _GEN_47 = 2'h3 == cacheLookUp_query_address[2:1] ? cacheLookUp_cacheDouble[63] : _GEN_46; // @[memAccess.scala 186:{24,24}]
  wire  _GEN_49 = cacheLookUp_query_address[2] ? cacheLookUp_cacheDouble[63] : cacheLookUp_cacheDouble[31]; // @[memAccess.scala 186:{24,24}]
  wire  _GEN_51 = 2'h1 == cacheLookUp_query_instruction[13:12] ? _GEN_47 : _GEN_43; // @[memAccess.scala 194:{25,25}]
  wire  _GEN_52 = 2'h2 == cacheLookUp_query_instruction[13:12] ? _GEN_49 : _GEN_51; // @[memAccess.scala 194:{25,25}]
  wire  _GEN_53 = 2'h3 == cacheLookUp_query_instruction[13:12] ? cacheLookUp_cacheDouble[63] : _GEN_52; // @[memAccess.scala 194:{25,25}]
  wire  _memoryResponse_readData_T_3 = ~cacheLookUp_query_instruction[14] & _GEN_53; // @[memAccess.scala 194:25]
  wire [55:0] _memoryResponse_readData_T_5 = _memoryResponse_readData_T_3 ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 77:12]
  wire [7:0] _GEN_55 = 3'h1 == cacheLookUp_query_address[2:0] ? cacheLookUp_cacheDouble[15:8] : cacheLookUp_cacheDouble[
    7:0]; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_56 = 3'h2 == cacheLookUp_query_address[2:0] ? cacheLookUp_cacheDouble[23:16] : _GEN_55; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_57 = 3'h3 == cacheLookUp_query_address[2:0] ? cacheLookUp_cacheDouble[31:24] : _GEN_56; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_58 = 3'h4 == cacheLookUp_query_address[2:0] ? cacheLookUp_cacheDouble[39:32] : _GEN_57; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_59 = 3'h5 == cacheLookUp_query_address[2:0] ? cacheLookUp_cacheDouble[47:40] : _GEN_58; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_60 = 3'h6 == cacheLookUp_query_address[2:0] ? cacheLookUp_cacheDouble[55:48] : _GEN_59; // @[Cat.scala 33:{92,92}]
  wire [7:0] _GEN_61 = 3'h7 == cacheLookUp_query_address[2:0] ? cacheLookUp_cacheDouble[63:56] : _GEN_60; // @[Cat.scala 33:{92,92}]
  wire [63:0] _memoryResponse_readData_T_15 = {_memoryResponse_readData_T_5,_GEN_61}; // @[Cat.scala 33:92]
  wire [47:0] _memoryResponse_readData_T_21 = _memoryResponse_readData_T_3 ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 77:12]
  wire [15:0] _GEN_63 = 2'h1 == cacheLookUp_query_address[2:1] ? cacheLookUp_cacheDouble[31:16] :
    cacheLookUp_cacheDouble[15:0]; // @[Cat.scala 33:{92,92}]
  wire [15:0] _GEN_64 = 2'h2 == cacheLookUp_query_address[2:1] ? cacheLookUp_cacheDouble[47:32] : _GEN_63; // @[Cat.scala 33:{92,92}]
  wire [15:0] _GEN_65 = 2'h3 == cacheLookUp_query_address[2:1] ? cacheLookUp_cacheDouble[63:48] : _GEN_64; // @[Cat.scala 33:{92,92}]
  wire [63:0] _memoryResponse_readData_T_27 = {_memoryResponse_readData_T_21,_GEN_65}; // @[Cat.scala 33:92]
  wire [31:0] _memoryResponse_readData_T_33 = _memoryResponse_readData_T_3 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _memoryResponse_readData_T_37 = {_memoryResponse_readData_T_33,
    memoryResponseWriteDataByteAligned_atomic32Src1}; // @[Cat.scala 33:92]
  wire [63:0] _GEN_69 = 2'h1 == cacheLookUp_query_instruction[13:12] ? _memoryResponse_readData_T_27 :
    _memoryResponse_readData_T_15; // @[memAccess.scala 185:{29,29}]
  wire  _memoryResponse_readData_T_44 = reservation64_valid & cacheLookUp_query_instruction[12] &
    _memoryResponseWriteDataByteAligned_semaphore64_T; // @[memAccess.scala 202:73]
  wire  _memoryResponse_readData_T_50 = reservation_valid & ~cacheLookUp_query_instruction[12] &
    _memoryResponseWriteDataByteAligned_semaphore32High_T_1; // @[memAccess.scala 203:72]
  wire  _memoryResponse_readData_T_51 = _memoryResponse_readData_T_44 | _memoryResponse_readData_T_50; // @[memAccess.scala 204:18]
  wire  _memoryResponse_readData_T_53 = ~((reservation_valid | reservation64_valid) & _memoryResponse_readData_T_51); // @[memAccess.scala 201:35]
  wire  _GEN_98 = branchOps_passed & cacheLookUp_query_valid; // @[memAccess.scala 176:26 271:30 272:47]
  wire  _GEN_100 = _missHandler_missedRequest_T_21 ? _GEN_98 : cacheLookUp_query_valid; // @[memAccess.scala 176:26 270:88]
  wire [31:0] _memoryResponse_query_address_T_1 = {missHandler_dependencyCheck_requset_address[31:12],
    missHandler_pushToCache_cacheWriteOut_address,3'h0}; // @[Cat.scala 33:92]
  wire  _GEN_101 = peripheralHandler_readFinished_ready & peripheralHandler_finishedRequest_valid; // @[memAccess.scala 286:52 288:26 168:30]
  wire  _GEN_108 = peripheralHandler_readFinished_ready | memoryResponse_hit; // @[memAccess.scala 286:52 290:24 96:31]
  wire  _GEN_110 = peripheralHandler_readFinished_ready; // @[memAccess.scala 173:40 286:52 293:42]
  wire  _GEN_112 = missHandler_pushToCache_ready ? 1'h0 : _GEN_101; // @[memAccess.scala 274:45 275:32]
  wire  _GEN_114 = missHandler_pushToCache_ready; // @[memAccess.scala 274:45 277:28]
  wire  _GEN_115 = missHandler_pushToCache_ready & missHandler_rlastToCache; // @[memAccess.scala 171:37 274:45 278:39]
  wire  _GEN_128 = missHandler_pushToCache_ready ? 1'h0 : _GEN_110; // @[memAccess.scala 173:40 274:45]
  wire  _GEN_130 = cacheLookUp_query_valid ? _GEN_100 : _GEN_112; // @[memAccess.scala 175:33]
  wire [6:0] _GEN_140 = cacheLookUp_query_valid ? cacheLookUp_query_address[12:6] : {{1'd0},
    memoryResponse_invalidate_cacheIndex}; // @[memAccess.scala 175:33 183:42 96:31]
  wire [2:0] _T_40 = {cacheLookUp_query_instruction[28],cacheLookUp_query_instruction[27],cacheLookUp_query_instruction[
    3]}; // @[Cat.scala 33:92]
  wire  _GEN_153 = cacheLookUp_query_instruction[12] | reservation64_valid; // @[memAccess.scala 300:{54,76} 38:30]
  wire [3:0] _T_50 = {cacheLookUp_query_instruction[28],cacheLookUp_query_instruction[27],cacheLookUp_query_instruction[
    5],cacheLookUp_query_instruction[3]}; // @[Cat.scala 33:92]
  wire  _GEN_157 = cacheLookUp_query_instruction[12] ? 1'h0 : reservation64_valid; // @[memAccess.scala 305:{54,76} 38:30]
  wire  _GEN_158 = cacheLookUp_query_instruction[12] & reservation_valid; // @[memAccess.scala 305:{119,54} 33:28]
  wire  _T_54 = ~missHandler_nonSaturatedReplay; // @[memAccess.scala 311:42]
  wire  _GEN_169 = cacheLookUp_query_address[31:6] == missHandler_dependencyCheck_requset_address[31:6] ? 1'h0 :
    _GEN_130; // @[memAccess.scala 315:136 316:36]
  wire  _GEN_170 = missHandler_handlerBusy & _T_54 ? _GEN_169 : _GEN_130; // @[memAccess.scala 314:76]
  wire  _GEN_171 = missHandler_handlerSaturated & ~missHandler_nonSaturatedReplay ? 1'h0 : _GEN_170; // @[memAccess.scala 311:76 313:34]
  wire  _GEN_172 = missHandler_missedRequest_query_valid ? 1'h0 : _GEN_171; // @[memAccess.scala 319:{49,78}]
  wire  _GEN_173 = cacheLookUp_query_valid ? _GEN_172 : _GEN_130; // @[memAccess.scala 310:33]
  wire  _T_66 = dataQueue_0_valid & dataQueue_1_valid; // @[memAccess.scala 351:45]
  wire  _T_67 = dataQueue_0_valid & dataQueue_1_valid & dataQueue_2_valid; // @[memAccess.scala 351:45]
  wire  dequeueData = scheduler_storeCommit_ready & dataQueue_0_valid & _missHandler_missedRequest_T_1 & ~
    scheduler_cacheStalled & ~scheduler_replaying; // @[memAccess.scala 356:126]
  reg  writeHandler_itWasPeripheral_REG; // @[memAccess.scala 488:58]
  reg  writeHandler_itWasPeripheral_REG_1; // @[memAccess.scala 488:50]
  reg  writeHandler_itWasPeripheral_REG_2; // @[memAccess.scala 488:42]
  wire [3:0] _T_69 = scheduler_toCache_queryWithData_query_branchMask & branchOps_branchMask; // @[memAccess.scala 507:58]
  wire  _T_70 = |_T_69; // @[memAccess.scala 507:82]
  wire [3:0] _servicing_query_branchMask_T = scheduler_toCache_queryWithData_query_branchMask ^ branchOps_branchMask; // @[memAccess.scala 507:107]
  wire [3:0] _T_71 = servicing_query_branchMask & branchOps_branchMask; // @[memAccess.scala 507:58]
  wire  _T_72 = |_T_71; // @[memAccess.scala 507:82]
  wire [3:0] _cacheLookUp_query_branchMask_T = servicing_query_branchMask ^ branchOps_branchMask; // @[memAccess.scala 507:107]
  wire [3:0] _T_80 = cacheLookUp_query_branchMask & branchOps_branchMask; // @[memAccess.scala 518:62]
  reg  waitForFenceData; // @[memAccess.scala 523:33]
  wire  _T_89 = ~(_missHandler_cachePipelineEmpty_T_1 | memoryResponse_query_valid) & (scheduler_clean &
    missHandler_clean & writeHandler_clean); // @[memAccess.scala 528:154]
  queryScheduler scheduler ( // @[memAccess.scala 13:25]
    .clock(scheduler_clock),
    .reset(scheduler_reset),
    .toCache_queryWithData_query_valid(scheduler_toCache_queryWithData_query_valid),
    .toCache_queryWithData_query_address(scheduler_toCache_queryWithData_query_address),
    .toCache_queryWithData_query_instruction(scheduler_toCache_queryWithData_query_instruction),
    .toCache_queryWithData_query_branchMask(scheduler_toCache_queryWithData_query_branchMask),
    .toCache_queryWithData_query_robAddr(scheduler_toCache_queryWithData_query_robAddr),
    .toCache_queryWithData_query_prfDest(scheduler_toCache_queryWithData_query_prfDest),
    .toCache_queryWithData_data(scheduler_toCache_queryWithData_data),
    .toCache_replaying(scheduler_toCache_replaying),
    .storeCommit_ready(scheduler_storeCommit_ready),
    .storeCommit_fired(scheduler_storeCommit_fired),
    .replaying(scheduler_replaying),
    .cacheStalled(scheduler_cacheStalled),
    .replayQueue_query_valid(scheduler_replayQueue_query_valid),
    .replayQueue_query_address(scheduler_replayQueue_query_address),
    .replayQueue_query_instruction(scheduler_replayQueue_query_instruction),
    .replayQueue_query_branchMask(scheduler_replayQueue_query_branchMask),
    .replayQueue_query_robAddr(scheduler_replayQueue_query_robAddr),
    .replayQueue_query_prfDest(scheduler_replayQueue_query_prfDest),
    .replayQueue_data(scheduler_replayQueue_data),
    .branchOps_valid(scheduler_branchOps_valid),
    .branchOps_branchMask(scheduler_branchOps_branchMask),
    .branchOps_passed(scheduler_branchOps_passed),
    .peripheral_ready(scheduler_peripheral_ready),
    .peripheral_bits_valid(scheduler_peripheral_bits_valid),
    .peripheral_bits_address(scheduler_peripheral_bits_address),
    .peripheral_bits_instruction(scheduler_peripheral_bits_instruction),
    .peripheral_bits_branchMask(scheduler_peripheral_bits_branchMask),
    .peripheral_bits_robAddr(scheduler_peripheral_bits_robAddr),
    .peripheral_bits_prfDest(scheduler_peripheral_bits_prfDest),
    .newInstruction_valid(scheduler_newInstruction_valid),
    .newInstruction_address(scheduler_newInstruction_address),
    .newInstruction_instruction(scheduler_newInstruction_instruction),
    .newInstruction_branchMask(scheduler_newInstruction_branchMask),
    .newInstruction_robAddr(scheduler_newInstruction_robAddr),
    .newInstruction_prfDest(scheduler_newInstruction_prfDest),
    .canAllocate(scheduler_canAllocate),
    .clean(scheduler_clean)
  );
  peripheralHandler peripheralHandler ( // @[memAccess.scala 19:33]
    .clock(peripheralHandler_clock),
    .reset(peripheralHandler_reset),
    .request_valid(peripheralHandler_request_valid),
    .request_address(peripheralHandler_request_address),
    .request_instruction(peripheralHandler_request_instruction),
    .request_branchMask(peripheralHandler_request_branchMask),
    .request_robAddr(peripheralHandler_request_robAddr),
    .request_prfDest(peripheralHandler_request_prfDest),
    .finishedRequest_valid(peripheralHandler_finishedRequest_valid),
    .finishedRequest_address(peripheralHandler_finishedRequest_address),
    .finishedRequest_instruction(peripheralHandler_finishedRequest_instruction),
    .finishedRequest_robAddr(peripheralHandler_finishedRequest_robAddr),
    .finishedRequest_prfDest(peripheralHandler_finishedRequest_prfDest),
    .ready(peripheralHandler_ready),
    .branchOps_valid(peripheralHandler_branchOps_valid),
    .branchOps_branchMask(peripheralHandler_branchOps_branchMask),
    .branchOps_passed(peripheralHandler_branchOps_passed),
    .axi_AWADDR(peripheralHandler_axi_AWADDR),
    .axi_AWLEN(peripheralHandler_axi_AWLEN),
    .axi_AWSIZE(peripheralHandler_axi_AWSIZE),
    .axi_AWVALID(peripheralHandler_axi_AWVALID),
    .axi_AWREADY(peripheralHandler_axi_AWREADY),
    .axi_WDATA(peripheralHandler_axi_WDATA),
    .axi_WSTRB(peripheralHandler_axi_WSTRB),
    .axi_WLAST(peripheralHandler_axi_WLAST),
    .axi_WVALID(peripheralHandler_axi_WVALID),
    .axi_WREADY(peripheralHandler_axi_WREADY),
    .axi_BVALID(peripheralHandler_axi_BVALID),
    .axi_BREADY(peripheralHandler_axi_BREADY),
    .axi_ARADDR(peripheralHandler_axi_ARADDR),
    .axi_ARLEN(peripheralHandler_axi_ARLEN),
    .axi_ARSIZE(peripheralHandler_axi_ARSIZE),
    .axi_ARVALID(peripheralHandler_axi_ARVALID),
    .axi_ARREADY(peripheralHandler_axi_ARREADY),
    .axi_RDATA(peripheralHandler_axi_RDATA),
    .axi_RLAST(peripheralHandler_axi_RLAST),
    .axi_RVALID(peripheralHandler_axi_RVALID),
    .axi_RREADY(peripheralHandler_axi_RREADY),
    .readFinished_ready(peripheralHandler_readFinished_ready),
    .readFinished_fired(peripheralHandler_readFinished_fired),
    .readDataOut(peripheralHandler_readDataOut),
    .writeIn_valid(peripheralHandler_writeIn_valid),
    .writeIn_data(peripheralHandler_writeIn_data)
  );
  zeroWriteLatencyCache cache ( // @[memAccess.scala 46:21]
    .clock(cache_clock),
    .reset(cache_reset),
    .readAddress(cache_readAddress),
    .readOut_0_data(cache_readOut_0_data),
    .readOut_0_tag(cache_readOut_0_tag),
    .readOut_0_valid(cache_readOut_0_valid),
    .readOut_1_data(cache_readOut_1_data),
    .readOut_1_tag(cache_readOut_1_tag),
    .readOut_1_valid(cache_readOut_1_valid),
    .writePorts_0_enable(cache_writePorts_0_enable),
    .writePorts_0_cacheAddress(cache_writePorts_0_cacheAddress),
    .writePorts_0_data(cache_writePorts_0_data),
    .writePorts_1_enable(cache_writePorts_1_enable),
    .writePorts_1_cacheAddress(cache_writePorts_1_cacheAddress),
    .writePorts_1_data(cache_writePorts_1_data),
    .invalidateSet_valid(cache_invalidateSet_valid),
    .invalidateSet_cacheIndex(cache_invalidateSet_cacheIndex),
    .invalidateSet_invalidateVector_0(cache_invalidateSet_invalidateVector_0),
    .invalidateSet_invalidateVector_1(cache_invalidateSet_invalidateVector_1),
    .cacheFillDone_valid(cache_cacheFillDone_valid),
    .cacheFillDone_cacheIndex(cache_cacheFillDone_cacheIndex),
    .cacheFillDone_validateVector_0(cache_cacheFillDone_validateVector_0),
    .cacheFillDone_validateVector_1(cache_cacheFillDone_validateVector_1),
    .cacheFillDone_tag(cache_cacheFillDone_tag)
  );
  missHandler missHandler ( // @[memAccess.scala 128:27]
    .clock(missHandler_clock),
    .reset(missHandler_reset),
    .replayOut_query_valid(missHandler_replayOut_query_valid),
    .replayOut_query_address(missHandler_replayOut_query_address),
    .replayOut_query_instruction(missHandler_replayOut_query_instruction),
    .replayOut_query_branchMask(missHandler_replayOut_query_branchMask),
    .replayOut_query_robAddr(missHandler_replayOut_query_robAddr),
    .replayOut_query_prfDest(missHandler_replayOut_query_prfDest),
    .replayOut_data(missHandler_replayOut_data),
    .replayingQuries(missHandler_replayingQuries),
    .branchOps_valid(missHandler_branchOps_valid),
    .branchOps_branchMask(missHandler_branchOps_branchMask),
    .branchOps_passed(missHandler_branchOps_passed),
    .cachePipelineEmpty(missHandler_cachePipelineEmpty),
    .missedRequest_query_valid(missHandler_missedRequest_query_valid),
    .missedRequest_query_address(missHandler_missedRequest_query_address),
    .missedRequest_query_instruction(missHandler_missedRequest_query_instruction),
    .missedRequest_query_branchMask(missHandler_missedRequest_query_branchMask),
    .missedRequest_query_robAddr(missHandler_missedRequest_query_robAddr),
    .missedRequest_query_prfDest(missHandler_missedRequest_query_prfDest),
    .missedRequest_data(missHandler_missedRequest_data),
    .pushToCache_ready(missHandler_pushToCache_ready),
    .pushToCache_fired(missHandler_pushToCache_fired),
    .pushToCache_cacheWriteOut_data(missHandler_pushToCache_cacheWriteOut_data),
    .pushToCache_cacheWriteOut_address(missHandler_pushToCache_cacheWriteOut_address),
    .pushToCache_cacheWriteOut_setSelVector(missHandler_pushToCache_cacheWriteOut_setSelVector),
    .axi_ARADDR(missHandler_axi_ARADDR),
    .axi_ARVALID(missHandler_axi_ARVALID),
    .axi_ARREADY(missHandler_axi_ARREADY),
    .axi_RDATA(missHandler_axi_RDATA),
    .axi_RLAST(missHandler_axi_RLAST),
    .axi_RVALID(missHandler_axi_RVALID),
    .axi_RREADY(missHandler_axi_RREADY),
    .dependencyCheck_requset_valid(missHandler_dependencyCheck_requset_valid),
    .dependencyCheck_requset_address(missHandler_dependencyCheck_requset_address),
    .dependencyCheck_free(missHandler_dependencyCheck_free),
    .rlastToCache(missHandler_rlastToCache),
    .setInvalidateVector(missHandler_setInvalidateVector),
    .setFillStatus(missHandler_setFillStatus),
    .handlerBusy(missHandler_handlerBusy),
    .handlerSaturated(missHandler_handlerSaturated),
    .clean(missHandler_clean),
    .nonSaturatedReplay(missHandler_nonSaturatedReplay)
  );
  writeHandler writeHandler ( // @[memAccess.scala 378:28]
    .clock(writeHandler_clock),
    .reset(writeHandler_reset),
    .itWasPeripheral(writeHandler_itWasPeripheral),
    .writeCommit_ready(writeHandler_writeCommit_ready),
    .writeCommit_fired(writeHandler_writeCommit_fired),
    .axi_AWADDR(writeHandler_axi_AWADDR),
    .axi_AWLEN(writeHandler_axi_AWLEN),
    .axi_AWSIZE(writeHandler_axi_AWSIZE),
    .axi_AWVALID(writeHandler_axi_AWVALID),
    .axi_AWREADY(writeHandler_axi_AWREADY),
    .axi_WDATA(writeHandler_axi_WDATA),
    .axi_WSTRB(writeHandler_axi_WSTRB),
    .axi_WLAST(writeHandler_axi_WLAST),
    .axi_WVALID(writeHandler_axi_WVALID),
    .axi_WREADY(writeHandler_axi_WREADY),
    .axi_BVALID(writeHandler_axi_BVALID),
    .axi_BREADY(writeHandler_axi_BREADY),
    .request_valid(writeHandler_request_valid),
    .request_address(writeHandler_request_address),
    .request_instruction(writeHandler_request_instruction),
    .request_alignedData(writeHandler_request_alignedData),
    .request_mask(writeHandler_request_mask),
    .dependencyCheck_requset_valid(writeHandler_dependencyCheck_requset_valid),
    .dependencyCheck_requset_address(writeHandler_dependencyCheck_requset_address),
    .dependencyCheck_free(writeHandler_dependencyCheck_free),
    .clean(writeHandler_clean)
  );
  assign peripheral_AWADDR = peripheralHandler_axi_AWADDR; // @[memAccess.scala 22:14]
  assign peripheral_AWLEN = peripheralHandler_axi_AWLEN; // @[memAccess.scala 22:14]
  assign peripheral_AWSIZE = peripheralHandler_axi_AWSIZE; // @[memAccess.scala 22:14]
  assign peripheral_AWVALID = peripheralHandler_axi_AWVALID; // @[memAccess.scala 22:14]
  assign peripheral_WDATA = peripheralHandler_axi_WDATA; // @[memAccess.scala 22:14]
  assign peripheral_WSTRB = peripheralHandler_axi_WSTRB; // @[memAccess.scala 22:14]
  assign peripheral_WLAST = peripheralHandler_axi_WLAST; // @[memAccess.scala 22:14]
  assign peripheral_WVALID = peripheralHandler_axi_WVALID; // @[memAccess.scala 22:14]
  assign peripheral_BREADY = peripheralHandler_axi_BREADY; // @[memAccess.scala 22:14]
  assign peripheral_ARADDR = peripheralHandler_axi_ARADDR; // @[memAccess.scala 22:14]
  assign peripheral_ARLEN = peripheralHandler_axi_ARLEN; // @[memAccess.scala 22:14]
  assign peripheral_ARSIZE = peripheralHandler_axi_ARSIZE; // @[memAccess.scala 22:14]
  assign peripheral_ARVALID = peripheralHandler_axi_ARVALID; // @[memAccess.scala 22:14]
  assign peripheral_RREADY = peripheralHandler_axi_RREADY; // @[memAccess.scala 22:14]
  assign responseOut_valid = memoryResponse_query_valid & memoryResponse_hit & memoryResponse_query_instruction[6:5] != 2'h1
    ; // @[memAccess.scala 344:73]
  assign responseOut_prfDest = memoryResponse_query_prfDest; // @[memAccess.scala 345:23]
  assign responseOut_robAddr = memoryResponse_query_robAddr; // @[memAccess.scala 346:23]
  assign responseOut_result = memoryResponse_readData; // @[memAccess.scala 347:22]
  assign responseOut_instruction = memoryResponse_query_instruction; // @[memAccess.scala 348:27]
  assign dPort_AWADDR = writeHandler_axi_AWADDR; // @[memAccess.scala 473:51]
  assign dPort_AWLEN = writeHandler_axi_AWLEN; // @[memAccess.scala 473:51]
  assign dPort_AWSIZE = writeHandler_axi_AWSIZE; // @[memAccess.scala 473:51]
  assign dPort_AWVALID = writeHandler_axi_AWVALID; // @[memAccess.scala 473:51]
  assign dPort_WDATA = writeHandler_axi_WDATA; // @[memAccess.scala 473:51]
  assign dPort_WSTRB = writeHandler_axi_WSTRB; // @[memAccess.scala 473:51]
  assign dPort_WLAST = writeHandler_axi_WLAST; // @[memAccess.scala 473:51]
  assign dPort_WVALID = writeHandler_axi_WVALID; // @[memAccess.scala 473:51]
  assign dPort_BREADY = writeHandler_axi_BREADY; // @[memAccess.scala 473:51]
  assign dPort_ARADDR = missHandler_axi_ARADDR; // @[memAccess.scala 473:51]
  assign dPort_ARVALID = missHandler_axi_ARVALID; // @[memAccess.scala 473:51]
  assign dPort_RREADY = missHandler_axi_RREADY; // @[memAccess.scala 473:51]
  assign writeCommit_ready = writeHandler_writeCommit_ready & ~(scheduler_cacheStalled | scheduler_replaying); // @[memAccess.scala 492:55]
  assign canAllocate = scheduler_canAllocate; // @[memAccess.scala 496:15]
  assign fenceInstructions_ready = ~waitForFenceData ? 1'h0 : _T_89; // @[memAccess.scala 525:27 527:27]
  assign scheduler_clock = clock;
  assign scheduler_reset = reset;
  assign scheduler_storeCommit_fired = scheduler_storeCommit_ready & dataQueue_0_valid & _missHandler_missedRequest_T_1
     & ~scheduler_cacheStalled & ~scheduler_replaying; // @[memAccess.scala 356:126]
  assign scheduler_replaying = missHandler_replayingQuries; // @[memAccess.scala 371:23]
  assign scheduler_cacheStalled = missHandler_handlerSaturated; // @[memAccess.scala 367:26]
  assign scheduler_replayQueue_query_valid = missHandler_replayOut_query_valid; // @[memAccess.scala 373:25]
  assign scheduler_replayQueue_query_address = missHandler_replayOut_query_address; // @[memAccess.scala 373:25]
  assign scheduler_replayQueue_query_instruction = missHandler_replayOut_query_instruction; // @[memAccess.scala 373:25]
  assign scheduler_replayQueue_query_branchMask = missHandler_replayOut_query_branchMask; // @[memAccess.scala 373:25]
  assign scheduler_replayQueue_query_robAddr = missHandler_replayOut_query_robAddr; // @[memAccess.scala 373:25]
  assign scheduler_replayQueue_query_prfDest = missHandler_replayOut_query_prfDest; // @[memAccess.scala 373:25]
  assign scheduler_replayQueue_data = missHandler_replayOut_data; // @[memAccess.scala 373:25]
  assign scheduler_branchOps_valid = branchOps_valid; // @[memAccess.scala 44:23]
  assign scheduler_branchOps_branchMask = branchOps_branchMask; // @[memAccess.scala 44:23]
  assign scheduler_branchOps_passed = branchOps_passed; // @[memAccess.scala 44:23]
  assign scheduler_peripheral_ready = peripheralHandler_ready; // @[memAccess.scala 24:30]
  assign scheduler_newInstruction_valid = request_valid; // @[memAccess.scala 376:28]
  assign scheduler_newInstruction_address = request_address; // @[memAccess.scala 376:28]
  assign scheduler_newInstruction_instruction = request_instruction; // @[memAccess.scala 376:28]
  assign scheduler_newInstruction_branchMask = request_branchMask; // @[memAccess.scala 376:28]
  assign scheduler_newInstruction_robAddr = request_robAddr; // @[memAccess.scala 376:28]
  assign scheduler_newInstruction_prfDest = request_prfDest; // @[memAccess.scala 376:28]
  assign peripheralHandler_clock = clock;
  assign peripheralHandler_reset = reset;
  assign peripheralHandler_request_valid = scheduler_peripheral_bits_valid; // @[memAccess.scala 25:29]
  assign peripheralHandler_request_address = scheduler_peripheral_bits_address; // @[memAccess.scala 25:29]
  assign peripheralHandler_request_instruction = scheduler_peripheral_bits_instruction; // @[memAccess.scala 25:29]
  assign peripheralHandler_request_branchMask = scheduler_peripheral_bits_branchMask; // @[memAccess.scala 25:29]
  assign peripheralHandler_request_robAddr = scheduler_peripheral_bits_robAddr; // @[memAccess.scala 25:29]
  assign peripheralHandler_request_prfDest = scheduler_peripheral_bits_prfDest; // @[memAccess.scala 25:29]
  assign peripheralHandler_branchOps_valid = branchOps_valid; // @[memAccess.scala 493:31]
  assign peripheralHandler_branchOps_branchMask = branchOps_branchMask; // @[memAccess.scala 493:31]
  assign peripheralHandler_branchOps_passed = branchOps_passed; // @[memAccess.scala 493:31]
  assign peripheralHandler_axi_AWREADY = peripheral_AWREADY; // @[memAccess.scala 22:14]
  assign peripheralHandler_axi_WREADY = peripheral_WREADY; // @[memAccess.scala 22:14]
  assign peripheralHandler_axi_BVALID = peripheral_BVALID; // @[memAccess.scala 22:14]
  assign peripheralHandler_axi_ARREADY = peripheral_ARREADY; // @[memAccess.scala 22:14]
  assign peripheralHandler_axi_RDATA = peripheral_RDATA; // @[memAccess.scala 22:14]
  assign peripheralHandler_axi_RLAST = peripheral_RLAST; // @[memAccess.scala 22:14]
  assign peripheralHandler_axi_RVALID = peripheral_RVALID; // @[memAccess.scala 22:14]
  assign peripheralHandler_readFinished_fired = cacheLookUp_query_valid ? 1'h0 : _GEN_128; // @[memAccess.scala 175:33 173:40]
  assign peripheralHandler_writeIn_valid = ~_T_2 & (scheduler_toCache_queryWithData_query_valid &
    scheduler_toCache_queryWithData_query_instruction[5]); // @[memAccess.scala 72:35 73:68 75:37]
  assign peripheralHandler_writeIn_data = dataToCache; // @[memAccess.scala 77:34]
  assign cache_clock = clock;
  assign cache_reset = reset;
  assign cache_readAddress = scheduler_toCache_queryWithData_query_address; // @[memAccess.scala 48:21]
  assign cache_writePorts_0_enable = memoryResponse_hitVector[0] & (_cacheLookUp_cacheDouble_T_13 |
    memoryResponse_filling); // @[memAccess.scala 327:32]
  assign cache_writePorts_0_cacheAddress = memoryResponse_query_address; // @[memAccess.scala 328:28]
  assign cache_writePorts_0_data = memoryResponse_write_dataByteAligned; // @[memAccess.scala 329:20]
  assign cache_writePorts_1_enable = memoryResponse_hitVector[1] & (_cacheLookUp_cacheDouble_T_13 |
    memoryResponse_filling); // @[memAccess.scala 327:32]
  assign cache_writePorts_1_cacheAddress = memoryResponse_query_address; // @[memAccess.scala 328:28]
  assign cache_writePorts_1_data = memoryResponse_write_dataByteAligned; // @[memAccess.scala 329:20]
  assign cache_invalidateSet_valid = memoryResponse_invalidate_valid; // @[memAccess.scala 334:23]
  assign cache_invalidateSet_cacheIndex = memoryResponse_invalidate_cacheIndex; // @[memAccess.scala 334:23]
  assign cache_invalidateSet_invalidateVector_0 = memoryResponse_invalidate_invalidateVector_0; // @[memAccess.scala 334:23]
  assign cache_invalidateSet_invalidateVector_1 = memoryResponse_invalidate_invalidateVector_1; // @[memAccess.scala 334:23]
  assign cache_cacheFillDone_valid = memoryResponse_cacheSetFill_valid; // @[memAccess.scala 332:23]
  assign cache_cacheFillDone_cacheIndex = memoryResponse_cacheSetFill_cacheIndex; // @[memAccess.scala 332:23]
  assign cache_cacheFillDone_validateVector_0 = memoryResponse_cacheSetFill_validateVector_0; // @[memAccess.scala 332:23]
  assign cache_cacheFillDone_validateVector_1 = memoryResponse_cacheSetFill_validateVector_1; // @[memAccess.scala 332:23]
  assign cache_cacheFillDone_tag = memoryResponse_cacheSetFill_tag; // @[memAccess.scala 332:23]
  assign missHandler_clock = clock;
  assign missHandler_reset = reset;
  assign missHandler_branchOps_valid = branchOps_valid; // @[memAccess.scala 166:25]
  assign missHandler_branchOps_branchMask = branchOps_branchMask; // @[memAccess.scala 166:25]
  assign missHandler_branchOps_passed = branchOps_passed; // @[memAccess.scala 166:25]
  assign missHandler_cachePipelineEmpty = ~_missHandler_cachePipelineEmpty_T_1; // @[memAccess.scala 158:37]
  assign missHandler_missedRequest_query_valid = branchOps_valid & |_missHandler_missedRequest_T_19 ? _GEN_33 : _GEN_31; // @[memAccess.scala 150:88]
  assign missHandler_missedRequest_query_address = cacheLookUp_query_address; // @[memAccess.scala 130:23 131:19]
  assign missHandler_missedRequest_query_instruction = cacheLookUp_query_instruction; // @[memAccess.scala 130:23 131:19]
  assign missHandler_missedRequest_query_branchMask = branchOps_valid & |_missHandler_missedRequest_T_19 ? _GEN_32 :
    cacheLookUp_query_branchMask; // @[memAccess.scala 131:19 150:88]
  assign missHandler_missedRequest_query_robAddr = cacheLookUp_query_robAddr; // @[memAccess.scala 130:23 131:19]
  assign missHandler_missedRequest_query_prfDest = cacheLookUp_query_prfDest; // @[memAccess.scala 130:23 131:19]
  assign missHandler_missedRequest_data = cacheLookUp_write_dataByteAligned >> _GEN_23; // @[memAccess.scala 132:55]
  assign missHandler_pushToCache_fired = missHandler_pushToCache_ready & ~cacheLookUp_query_valid; // @[memAccess.scala 321:66]
  assign missHandler_axi_ARREADY = dPort_ARREADY; // @[memAccess.scala 473:51]
  assign missHandler_axi_RDATA = dPort_RDATA; // @[memAccess.scala 473:51]
  assign missHandler_axi_RLAST = dPort_RLAST; // @[memAccess.scala 473:51]
  assign missHandler_axi_RVALID = dPort_RVALID; // @[memAccess.scala 473:51]
  assign missHandler_dependencyCheck_free = writeHandler_dependencyCheck_free; // @[memAccess.scala 389:32]
  assign missHandler_setFillStatus = cacheLookUp_setFillVector; // @[memAccess.scala 164:29]
  assign writeHandler_clock = clock;
  assign writeHandler_reset = reset;
  assign writeHandler_itWasPeripheral = writeHandler_itWasPeripheral_REG_2; // @[memAccess.scala 488:32]
  assign writeHandler_writeCommit_fired = writeCommit_fired; // @[memAccess.scala 491:15]
  assign writeHandler_axi_AWREADY = dPort_AWREADY; // @[memAccess.scala 473:51]
  assign writeHandler_axi_WREADY = dPort_WREADY; // @[memAccess.scala 473:51]
  assign writeHandler_axi_BVALID = dPort_BVALID; // @[memAccess.scala 473:51]
  assign writeHandler_request_valid = memoryResponse_query_valid & memoryResponse_query_instruction[5]; // @[memAccess.scala 387:60]
  assign writeHandler_request_address = memoryResponse_query_address; // @[memAccess.scala 380:32]
  assign writeHandler_request_instruction = memoryResponse_query_instruction; // @[memAccess.scala 382:36]
  assign writeHandler_request_alignedData = memoryResponse_write_dataByteAligned; // @[memAccess.scala 385:36]
  assign writeHandler_request_mask = memoryResponse_write_aligedMask; // @[memAccess.scala 386:29]
  assign writeHandler_dependencyCheck_requset_valid = missHandler_dependencyCheck_requset_valid; // @[memAccess.scala 389:32]
  assign writeHandler_dependencyCheck_requset_address = missHandler_dependencyCheck_requset_address; // @[memAccess.scala 389:32]
  always @(posedge clock) begin
    if (reset) begin // @[memAccess.scala 33:28]
      reservation_valid <= 1'h0; // @[memAccess.scala 33:28]
    end else if (cacheLookUp_query_valid & _missHandler_missedRequest_T_4) begin // @[memAccess.scala 298:62]
      if (_T_40 == 3'h5) begin // @[memAccess.scala 299:86]
        if (!(cacheLookUp_query_instruction[12])) begin // @[memAccess.scala 300:54]
          reservation_valid <= 1'h1; // @[memAccess.scala 300:118]
        end
      end else if (_T_50 == 4'hf) begin // @[memAccess.scala 304:97]
        reservation_valid <= _GEN_158;
      end
    end
    if (cacheLookUp_query_valid & _missHandler_missedRequest_T_4) begin // @[memAccess.scala 298:62]
      if (_T_40 == 3'h5) begin // @[memAccess.scala 299:86]
        if (!(cacheLookUp_query_instruction[12])) begin // @[memAccess.scala 301:54]
          reservation_address <= cacheLookUp_query_address; // @[memAccess.scala 303:41]
        end
      end
    end
    if (reset) begin // @[memAccess.scala 38:30]
      reservation64_valid <= 1'h0; // @[memAccess.scala 38:30]
    end else if (cacheLookUp_query_valid & _missHandler_missedRequest_T_4) begin // @[memAccess.scala 298:62]
      if (_T_40 == 3'h5) begin // @[memAccess.scala 299:86]
        reservation64_valid <= _GEN_153;
      end else if (_T_50 == 4'hf) begin // @[memAccess.scala 304:97]
        reservation64_valid <= _GEN_157;
      end
    end
    if (cacheLookUp_query_valid & _missHandler_missedRequest_T_4) begin // @[memAccess.scala 298:62]
      if (_T_40 == 3'h5) begin // @[memAccess.scala 299:86]
        if (cacheLookUp_query_instruction[12]) begin // @[memAccess.scala 301:54]
          reservation64_address <= cacheLookUp_query_address; // @[memAccess.scala 302:31]
        end
      end
    end
    if (reset) begin // @[memAccess.scala 52:26]
      dataQueue_0_valid <= 1'h0; // @[memAccess.scala 52:26]
    end else if (dequeueData) begin // @[memAccess.scala 361:21]
      if (dataQueue_0_valid & ~dataQueue_1_valid) begin // @[memAccess.scala 354:18]
        dataQueue_0_valid <= writeDataIn_valid;
      end else begin
        dataQueue_0_valid <= dataQueue_1_valid;
      end
    end else if (~dataQueue_0_valid) begin // @[memAccess.scala 354:18]
      dataQueue_0_valid <= writeDataIn_valid;
    end
    if (dequeueData) begin // @[memAccess.scala 361:21]
      if (dataQueue_0_valid & ~dataQueue_1_valid) begin // @[memAccess.scala 354:18]
        dataQueue_0_data <= writeDataIn_data;
      end else begin
        dataQueue_0_data <= dataQueue_1_data;
      end
    end else if (~dataQueue_0_valid) begin // @[memAccess.scala 354:18]
      dataQueue_0_data <= writeDataIn_data;
    end
    if (reset) begin // @[memAccess.scala 52:26]
      dataQueue_1_valid <= 1'h0; // @[memAccess.scala 52:26]
    end else if (dequeueData) begin // @[memAccess.scala 361:21]
      if (_T_66 & ~dataQueue_2_valid) begin // @[memAccess.scala 354:18]
        dataQueue_1_valid <= writeDataIn_valid;
      end else begin
        dataQueue_1_valid <= dataQueue_2_valid;
      end
    end else if (dataQueue_0_valid & ~dataQueue_1_valid) begin // @[memAccess.scala 354:18]
      dataQueue_1_valid <= writeDataIn_valid;
    end
    if (dequeueData) begin // @[memAccess.scala 361:21]
      if (_T_66 & ~dataQueue_2_valid) begin // @[memAccess.scala 354:18]
        dataQueue_1_data <= writeDataIn_data;
      end else begin
        dataQueue_1_data <= dataQueue_2_data;
      end
    end else if (dataQueue_0_valid & ~dataQueue_1_valid) begin // @[memAccess.scala 354:18]
      dataQueue_1_data <= writeDataIn_data;
    end
    if (reset) begin // @[memAccess.scala 52:26]
      dataQueue_2_valid <= 1'h0; // @[memAccess.scala 52:26]
    end else if (dequeueData) begin // @[memAccess.scala 361:21]
      if (_T_67 & ~dataQueue_3_valid) begin // @[memAccess.scala 354:18]
        dataQueue_2_valid <= writeDataIn_valid;
      end else begin
        dataQueue_2_valid <= dataQueue_3_valid;
      end
    end else if (_T_66 & ~dataQueue_2_valid) begin // @[memAccess.scala 354:18]
      dataQueue_2_valid <= writeDataIn_valid;
    end
    if (dequeueData) begin // @[memAccess.scala 361:21]
      if (_T_67 & ~dataQueue_3_valid) begin // @[memAccess.scala 354:18]
        dataQueue_2_data <= writeDataIn_data;
      end else begin
        dataQueue_2_data <= dataQueue_3_data;
      end
    end else if (_T_66 & ~dataQueue_2_valid) begin // @[memAccess.scala 354:18]
      dataQueue_2_data <= writeDataIn_data;
    end
    if (reset) begin // @[memAccess.scala 52:26]
      dataQueue_3_valid <= 1'h0; // @[memAccess.scala 52:26]
    end else if (dequeueData) begin // @[memAccess.scala 361:21]
      dataQueue_3_valid <= 1'h0; // @[memAccess.scala 363:41]
    end else if (_T_67 & ~dataQueue_3_valid) begin // @[memAccess.scala 354:18]
      dataQueue_3_valid <= writeDataIn_valid;
    end
    if (_T_67 & ~dataQueue_3_valid) begin // @[memAccess.scala 354:18]
      dataQueue_3_data <= writeDataIn_data;
    end
    if (dequeueData) begin // @[memAccess.scala 361:21]
      dataToCache <= dataQueue_0_data; // @[memAccess.scala 364:17]
    end
    if (reset) begin // @[memAccess.scala 61:26]
      servicing_query_valid <= 1'h0; // @[memAccess.scala 61:26]
    end else if (branchOps_valid) begin // @[memAccess.scala 498:25]
      if (~branchOps_passed) begin // @[memAccess.scala 509:29]
        if (_T_70) begin // @[memAccess.scala 518:91]
          servicing_query_valid <= 1'h0; // @[memAccess.scala 518:102]
        end else begin
          servicing_query_valid <= _GEN_2;
        end
      end else begin
        servicing_query_valid <= _GEN_2;
      end
    end else begin
      servicing_query_valid <= _GEN_2;
    end
    servicing_query_address <= scheduler_toCache_queryWithData_query_address; // @[memAccess.scala 63:19]
    servicing_query_instruction <= scheduler_toCache_queryWithData_query_instruction; // @[memAccess.scala 63:19]
    if (branchOps_valid) begin // @[memAccess.scala 498:25]
      if (|_T_69) begin // @[memAccess.scala 507:87]
        servicing_query_branchMask <= _servicing_query_branchMask_T; // @[memAccess.scala 507:96]
      end else begin
        servicing_query_branchMask <= scheduler_toCache_queryWithData_query_branchMask; // @[memAccess.scala 63:19]
      end
    end else begin
      servicing_query_branchMask <= scheduler_toCache_queryWithData_query_branchMask; // @[memAccess.scala 63:19]
    end
    servicing_query_robAddr <= scheduler_toCache_queryWithData_query_robAddr; // @[memAccess.scala 63:19]
    servicing_query_prfDest <= scheduler_toCache_queryWithData_query_prfDest; // @[memAccess.scala 63:19]
    if (scheduler_toCache_replaying) begin // @[memAccess.scala 64:37]
      servicing_data <= scheduler_toCache_queryWithData_data; // @[memAccess.scala 64:54]
    end else if (|scheduler_toCache_queryWithData_query_instruction[24:20]) begin // @[memAccess.scala 67:73]
      servicing_data <= dataToCache; // @[memAccess.scala 68:22]
    end else begin
      servicing_data <= 64'h0; // @[memAccess.scala 66:20]
    end
    if (reset) begin // @[memAccess.scala 79:28]
      cacheLookUp_query_valid <= 1'h0; // @[memAccess.scala 79:28]
    end else if (branchOps_valid) begin // @[memAccess.scala 498:25]
      if (~branchOps_passed) begin // @[memAccess.scala 509:29]
        if (_T_72) begin // @[memAccess.scala 518:91]
          cacheLookUp_query_valid <= 1'h0; // @[memAccess.scala 518:102]
        end else begin
          cacheLookUp_query_valid <= servicing_query_valid; // @[memAccess.scala 89:21]
        end
      end else begin
        cacheLookUp_query_valid <= servicing_query_valid; // @[memAccess.scala 89:21]
      end
    end else begin
      cacheLookUp_query_valid <= servicing_query_valid; // @[memAccess.scala 89:21]
    end
    cacheLookUp_query_address <= servicing_query_address; // @[memAccess.scala 89:21]
    cacheLookUp_query_instruction <= servicing_query_instruction; // @[memAccess.scala 89:21]
    if (branchOps_valid) begin // @[memAccess.scala 498:25]
      if (|_T_71) begin // @[memAccess.scala 507:87]
        cacheLookUp_query_branchMask <= _cacheLookUp_query_branchMask_T; // @[memAccess.scala 507:96]
      end else begin
        cacheLookUp_query_branchMask <= servicing_query_branchMask; // @[memAccess.scala 89:21]
      end
    end else begin
      cacheLookUp_query_branchMask <= servicing_query_branchMask; // @[memAccess.scala 89:21]
    end
    cacheLookUp_query_robAddr <= servicing_query_robAddr; // @[memAccess.scala 89:21]
    cacheLookUp_query_prfDest <= servicing_query_prfDest; // @[memAccess.scala 89:21]
    cacheLookUp_write_dataByteAligned <= _cacheLookUp_write_dataByteAligned_T_1[63:0]; // @[memAccess.scala 92:37]
    cacheLookUp_write_aligedMask <= _cacheLookUp_write_aligedMask_T_2[7:0]; // @[memAccess.scala 93:32]
    cacheLookUp_hitVector <= {_cacheLookUp_hitVector_T_5,_cacheLookUp_hitVector_T_2}; // @[Cat.scala 33:92]
    cacheLookUp_setFillVector <= {cache_readOut_1_valid,cache_readOut_0_valid}; // @[Cat.scala 33:92]
    if (_cacheLookUp_cacheDouble_T_10) begin // @[Mux.scala 101:16]
      if (cacheLookUp_query_valid) begin // @[memAccess.scala 175:33]
        if (cacheLookUp_query_instruction[3]) begin // @[memAccess.scala 266:10]
          if (cacheLookUp_query_instruction[12]) begin // @[memAccess.scala 264:23]
            cacheLookUp_cacheDouble <= memoryResponseWriteDataByteAligned_atomic64;
          end else begin
            cacheLookUp_cacheDouble <= _GEN_96;
          end
        end else begin
          cacheLookUp_cacheDouble <= memoryResponseWriteDataByteAligned_storeData;
        end
      end else begin
        cacheLookUp_cacheDouble <= 64'h0;
      end
    end else if (_cacheLookUp_cacheDouble_T_17) begin // @[Mux.scala 101:16]
      cacheLookUp_cacheDouble <= memoryResponse_write_dataByteAligned;
    end else if (_cacheLookUp_hitVector_T_5) begin // @[Mux.scala 101:16]
      cacheLookUp_cacheDouble <= cache_readOut_1_data;
    end else begin
      cacheLookUp_cacheDouble <= cache_readOut_0_data;
    end
    if (reset) begin // @[memAccess.scala 96:31]
      memoryResponse_query_valid <= 1'h0; // @[memAccess.scala 96:31]
    end else if (branchOps_valid) begin // @[memAccess.scala 498:25]
      if (~branchOps_passed) begin // @[memAccess.scala 509:29]
        if (|_T_80) begin // @[memAccess.scala 518:91]
          memoryResponse_query_valid <= 1'h0; // @[memAccess.scala 518:102]
        end else begin
          memoryResponse_query_valid <= _GEN_173;
        end
      end else begin
        memoryResponse_query_valid <= _GEN_173;
      end
    end else begin
      memoryResponse_query_valid <= _GEN_173;
    end
    if (cacheLookUp_query_valid) begin // @[memAccess.scala 175:33]
      memoryResponse_query_address <= cacheLookUp_query_address; // @[memAccess.scala 176:26]
    end else if (missHandler_pushToCache_ready) begin // @[memAccess.scala 274:45]
      memoryResponse_query_address <= _memoryResponse_query_address_T_1; // @[memAccess.scala 276:34]
    end else if (peripheralHandler_readFinished_ready) begin // @[memAccess.scala 286:52]
      memoryResponse_query_address <= peripheralHandler_finishedRequest_address; // @[memAccess.scala 288:26]
    end
    if (cacheLookUp_query_valid) begin // @[memAccess.scala 175:33]
      memoryResponse_query_instruction <= cacheLookUp_query_instruction; // @[memAccess.scala 176:26]
    end else if (!(missHandler_pushToCache_ready)) begin // @[memAccess.scala 274:45]
      if (peripheralHandler_readFinished_ready) begin // @[memAccess.scala 286:52]
        memoryResponse_query_instruction <= peripheralHandler_finishedRequest_instruction; // @[memAccess.scala 288:26]
      end
    end
    if (cacheLookUp_query_valid) begin // @[memAccess.scala 175:33]
      memoryResponse_query_robAddr <= cacheLookUp_query_robAddr; // @[memAccess.scala 176:26]
    end else if (!(missHandler_pushToCache_ready)) begin // @[memAccess.scala 274:45]
      if (peripheralHandler_readFinished_ready) begin // @[memAccess.scala 286:52]
        memoryResponse_query_robAddr <= peripheralHandler_finishedRequest_robAddr; // @[memAccess.scala 288:26]
      end
    end
    if (cacheLookUp_query_valid) begin // @[memAccess.scala 175:33]
      memoryResponse_query_prfDest <= cacheLookUp_query_prfDest; // @[memAccess.scala 176:26]
    end else if (!(missHandler_pushToCache_ready)) begin // @[memAccess.scala 274:45]
      if (peripheralHandler_readFinished_ready) begin // @[memAccess.scala 286:52]
        memoryResponse_query_prfDest <= peripheralHandler_finishedRequest_prfDest; // @[memAccess.scala 288:26]
      end
    end
    if (cacheLookUp_query_valid) begin // @[memAccess.scala 175:33]
      if (cacheLookUp_query_valid) begin // @[memAccess.scala 175:33]
        if (cacheLookUp_query_instruction[3]) begin // @[memAccess.scala 266:10]
          if (cacheLookUp_query_instruction[12]) begin // @[memAccess.scala 264:23]
            memoryResponse_write_dataByteAligned <= memoryResponseWriteDataByteAligned_atomic64;
          end else begin
            memoryResponse_write_dataByteAligned <= _GEN_96;
          end
        end else begin
          memoryResponse_write_dataByteAligned <= memoryResponseWriteDataByteAligned_storeData;
        end
      end else begin
        memoryResponse_write_dataByteAligned <= 64'h0;
      end
    end else if (missHandler_pushToCache_ready) begin // @[memAccess.scala 274:45]
      memoryResponse_write_dataByteAligned <= missHandler_pushToCache_cacheWriteOut_data; // @[memAccess.scala 284:42]
    end
    if (cacheLookUp_query_valid) begin // @[memAccess.scala 175:33]
      memoryResponse_write_aligedMask <= cacheLookUp_write_aligedMask; // @[memAccess.scala 269:37]
    end
    if (cacheLookUp_query_valid) begin // @[memAccess.scala 175:33]
      memoryResponse_hit <= _missHandler_missedRequest_T_4; // @[memAccess.scala 179:24]
    end else if (missHandler_pushToCache_ready) begin // @[memAccess.scala 274:45]
      memoryResponse_hit <= 1'h0; // @[memAccess.scala 281:24]
    end else begin
      memoryResponse_hit <= _GEN_108;
    end
    if (cacheLookUp_query_valid) begin // @[memAccess.scala 175:33]
      memoryResponse_hitVector <= cacheLookUp_hitVector; // @[memAccess.scala 206:30]
    end else if (missHandler_pushToCache_ready) begin // @[memAccess.scala 274:45]
      memoryResponse_hitVector <= missHandler_pushToCache_cacheWriteOut_setSelVector; // @[memAccess.scala 282:30]
    end else if (peripheralHandler_readFinished_ready) begin // @[memAccess.scala 286:52]
      memoryResponse_hitVector <= 2'h1; // @[memAccess.scala 291:30]
    end
    if (cacheLookUp_query_valid) begin // @[memAccess.scala 175:33]
      if (cacheLookUp_query_instruction[3]) begin // @[memAccess.scala 200:51]
        memoryResponse_readData <= {{63'd0}, _memoryResponse_readData_T_53}; // @[memAccess.scala 201:31]
      end else if (2'h3 == cacheLookUp_query_instruction[13:12]) begin // @[memAccess.scala 185:29]
        memoryResponse_readData <= cacheLookUp_cacheDouble; // @[memAccess.scala 185:29]
      end else if (2'h2 == cacheLookUp_query_instruction[13:12]) begin // @[memAccess.scala 185:29]
        memoryResponse_readData <= _memoryResponse_readData_T_37; // @[memAccess.scala 185:29]
      end else begin
        memoryResponse_readData <= _GEN_69;
      end
    end else if (!(missHandler_pushToCache_ready)) begin // @[memAccess.scala 274:45]
      if (peripheralHandler_readFinished_ready) begin // @[memAccess.scala 286:52]
        memoryResponse_readData <= peripheralHandler_readDataOut; // @[memAccess.scala 294:29]
      end
    end
    memoryResponse_invalidate_valid <= cacheLookUp_query_valid & (&cacheLookUp_setFillVector &
      _missHandler_missedRequest_T_1 & cacheLookUp_query_valid & ~_missHandler_missedRequest_T_4); // @[memAccess.scala 175:33 182:37]
    memoryResponse_invalidate_cacheIndex <= _GEN_140[5:0];
    if (cacheLookUp_query_valid) begin // @[memAccess.scala 175:33]
      memoryResponse_invalidate_invalidateVector_0 <= missHandler_setInvalidateVector[0]; // @[memAccess.scala 184:48]
    end
    if (cacheLookUp_query_valid) begin // @[memAccess.scala 175:33]
      memoryResponse_invalidate_invalidateVector_1 <= missHandler_setInvalidateVector[1]; // @[memAccess.scala 184:48]
    end
    if (cacheLookUp_query_valid) begin // @[memAccess.scala 175:33]
      memoryResponse_cacheSetFill_valid <= 1'h0; // @[memAccess.scala 177:39]
    end else begin
      memoryResponse_cacheSetFill_valid <= _GEN_115;
    end
    if (!(cacheLookUp_query_valid)) begin // @[memAccess.scala 175:33]
      if (missHandler_pushToCache_ready) begin // @[memAccess.scala 274:45]
        memoryResponse_cacheSetFill_cacheIndex <= missHandler_pushToCache_cacheWriteOut_address[8:3]; // @[memAccess.scala 279:44]
      end
    end
    if (!(cacheLookUp_query_valid)) begin // @[memAccess.scala 175:33]
      if (missHandler_pushToCache_ready) begin // @[memAccess.scala 274:45]
        memoryResponse_cacheSetFill_validateVector_0 <= missHandler_pushToCache_cacheWriteOut_setSelVector[0]; // @[memAccess.scala 280:48]
      end
    end
    if (!(cacheLookUp_query_valid)) begin // @[memAccess.scala 175:33]
      if (missHandler_pushToCache_ready) begin // @[memAccess.scala 274:45]
        memoryResponse_cacheSetFill_validateVector_1 <= missHandler_pushToCache_cacheWriteOut_setSelVector[1]; // @[memAccess.scala 280:48]
      end
    end
    if (!(cacheLookUp_query_valid)) begin // @[memAccess.scala 175:33]
      if (missHandler_pushToCache_ready) begin // @[memAccess.scala 274:45]
        memoryResponse_cacheSetFill_tag <= missHandler_dependencyCheck_requset_address[31:12]; // @[memAccess.scala 285:37]
      end
    end
    if (reset) begin // @[memAccess.scala 96:31]
      memoryResponse_filling <= 1'h0; // @[memAccess.scala 96:31]
    end else if (cacheLookUp_query_valid) begin // @[memAccess.scala 175:33]
      memoryResponse_filling <= 1'h0; // @[memAccess.scala 180:28]
    end else begin
      memoryResponse_filling <= _GEN_114;
    end
    if (reset) begin // @[memAccess.scala 488:58]
      writeHandler_itWasPeripheral_REG <= 1'h0; // @[memAccess.scala 488:58]
    end else begin
      writeHandler_itWasPeripheral_REG <= peripheralHandler_writeIn_valid; // @[memAccess.scala 488:58]
    end
    if (reset) begin // @[memAccess.scala 488:50]
      writeHandler_itWasPeripheral_REG_1 <= 1'h0; // @[memAccess.scala 488:50]
    end else begin
      writeHandler_itWasPeripheral_REG_1 <= writeHandler_itWasPeripheral_REG; // @[memAccess.scala 488:50]
    end
    if (reset) begin // @[memAccess.scala 488:42]
      writeHandler_itWasPeripheral_REG_2 <= 1'h0; // @[memAccess.scala 488:42]
    end else begin
      writeHandler_itWasPeripheral_REG_2 <= writeHandler_itWasPeripheral_REG_1; // @[memAccess.scala 488:42]
    end
    if (reset) begin // @[memAccess.scala 523:33]
      waitForFenceData <= 1'h0; // @[memAccess.scala 523:33]
    end else if (~waitForFenceData) begin // @[memAccess.scala 527:27]
      waitForFenceData <= initiateFence; // @[memAccess.scala 527:46]
    end else if (~(_missHandler_cachePipelineEmpty_T_1 | memoryResponse_query_valid) & (scheduler_clean &
      missHandler_clean & writeHandler_clean)) begin // @[memAccess.scala 528:233]
      if (fenceInstructions_fired) begin // @[memAccess.scala 530:35]
        waitForFenceData <= 1'h0; // @[memAccess.scala 530:54]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reservation_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reservation_address = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reservation64_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  reservation64_address = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  dataQueue_0_valid = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  dataQueue_0_data = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  dataQueue_1_valid = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  dataQueue_1_data = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  dataQueue_2_valid = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  dataQueue_2_data = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  dataQueue_3_valid = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  dataQueue_3_data = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  dataToCache = _RAND_12[63:0];
  _RAND_13 = {1{`RANDOM}};
  servicing_query_valid = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  servicing_query_address = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  servicing_query_instruction = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  servicing_query_branchMask = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  servicing_query_robAddr = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  servicing_query_prfDest = _RAND_18[5:0];
  _RAND_19 = {2{`RANDOM}};
  servicing_data = _RAND_19[63:0];
  _RAND_20 = {1{`RANDOM}};
  cacheLookUp_query_valid = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  cacheLookUp_query_address = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  cacheLookUp_query_instruction = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  cacheLookUp_query_branchMask = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  cacheLookUp_query_robAddr = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  cacheLookUp_query_prfDest = _RAND_25[5:0];
  _RAND_26 = {2{`RANDOM}};
  cacheLookUp_write_dataByteAligned = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  cacheLookUp_write_aligedMask = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  cacheLookUp_hitVector = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  cacheLookUp_setFillVector = _RAND_29[1:0];
  _RAND_30 = {2{`RANDOM}};
  cacheLookUp_cacheDouble = _RAND_30[63:0];
  _RAND_31 = {1{`RANDOM}};
  memoryResponse_query_valid = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  memoryResponse_query_address = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  memoryResponse_query_instruction = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  memoryResponse_query_robAddr = _RAND_34[3:0];
  _RAND_35 = {1{`RANDOM}};
  memoryResponse_query_prfDest = _RAND_35[5:0];
  _RAND_36 = {2{`RANDOM}};
  memoryResponse_write_dataByteAligned = _RAND_36[63:0];
  _RAND_37 = {1{`RANDOM}};
  memoryResponse_write_aligedMask = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  memoryResponse_hit = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  memoryResponse_hitVector = _RAND_39[1:0];
  _RAND_40 = {2{`RANDOM}};
  memoryResponse_readData = _RAND_40[63:0];
  _RAND_41 = {1{`RANDOM}};
  memoryResponse_invalidate_valid = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  memoryResponse_invalidate_cacheIndex = _RAND_42[5:0];
  _RAND_43 = {1{`RANDOM}};
  memoryResponse_invalidate_invalidateVector_0 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  memoryResponse_invalidate_invalidateVector_1 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  memoryResponse_cacheSetFill_valid = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  memoryResponse_cacheSetFill_cacheIndex = _RAND_46[5:0];
  _RAND_47 = {1{`RANDOM}};
  memoryResponse_cacheSetFill_validateVector_0 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  memoryResponse_cacheSetFill_validateVector_1 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  memoryResponse_cacheSetFill_tag = _RAND_49[19:0];
  _RAND_50 = {1{`RANDOM}};
  memoryResponse_filling = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  writeHandler_itWasPeripheral_REG = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  writeHandler_itWasPeripheral_REG_1 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  writeHandler_itWasPeripheral_REG_2 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  waitForFenceData = _RAND_54[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReadWriteSmem(
  input         clock,
  input         io_wenable,
  input         io_renable,
  input  [5:0]  io_raddr,
  input  [5:0]  io_waddr,
  input  [63:0] io_dataIn,
  output [63:0] io_dataOut
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mem [0:63]; // @[SRAM_block.scala 15:24]
  wire  mem_io_dataOut_MPORT_en; // @[SRAM_block.scala 15:24]
  wire [5:0] mem_io_dataOut_MPORT_addr; // @[SRAM_block.scala 15:24]
  wire [63:0] mem_io_dataOut_MPORT_data; // @[SRAM_block.scala 15:24]
  wire [63:0] mem_MPORT_data; // @[SRAM_block.scala 15:24]
  wire [5:0] mem_MPORT_addr; // @[SRAM_block.scala 15:24]
  wire  mem_MPORT_mask; // @[SRAM_block.scala 15:24]
  wire  mem_MPORT_en; // @[SRAM_block.scala 15:24]
  reg  mem_io_dataOut_MPORT_en_pipe_0;
  reg [5:0] mem_io_dataOut_MPORT_addr_pipe_0;
  assign mem_io_dataOut_MPORT_en = mem_io_dataOut_MPORT_en_pipe_0;
  assign mem_io_dataOut_MPORT_addr = mem_io_dataOut_MPORT_addr_pipe_0;
  assign mem_io_dataOut_MPORT_data = mem[mem_io_dataOut_MPORT_addr]; // @[SRAM_block.scala 15:24]
  assign mem_MPORT_data = io_dataIn;
  assign mem_MPORT_addr = io_waddr;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_wenable;
  assign io_dataOut = mem_io_dataOut_MPORT_data; // @[SRAM_block.scala 21:14]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SRAM_block.scala 15:24]
    end
    mem_io_dataOut_MPORT_en_pipe_0 <= io_renable;
    if (io_renable) begin
      mem_io_dataOut_MPORT_addr_pipe_0 <= io_raddr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    mem[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_dataOut_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_dataOut_MPORT_addr_pipe_0 = _RAND_2[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LVT_set(
  input         clock,
  input         io_wenable,
  input         io_r1enable,
  input         io_r2enable,
  input         io_r3enable,
  input  [5:0]  io_r1addr,
  input  [5:0]  io_r2addr,
  input  [5:0]  io_r3addr,
  input  [5:0]  io_waddr,
  input  [63:0] io_wdata,
  output [63:0] io_r1data,
  output [63:0] io_r2data,
  output [63:0] io_r3data
);
  wire  b1_clock; // @[LVT_set.scala 20:18]
  wire  b1_io_wenable; // @[LVT_set.scala 20:18]
  wire  b1_io_renable; // @[LVT_set.scala 20:18]
  wire [5:0] b1_io_raddr; // @[LVT_set.scala 20:18]
  wire [5:0] b1_io_waddr; // @[LVT_set.scala 20:18]
  wire [63:0] b1_io_dataIn; // @[LVT_set.scala 20:18]
  wire [63:0] b1_io_dataOut; // @[LVT_set.scala 20:18]
  wire  b2_clock; // @[LVT_set.scala 21:18]
  wire  b2_io_wenable; // @[LVT_set.scala 21:18]
  wire  b2_io_renable; // @[LVT_set.scala 21:18]
  wire [5:0] b2_io_raddr; // @[LVT_set.scala 21:18]
  wire [5:0] b2_io_waddr; // @[LVT_set.scala 21:18]
  wire [63:0] b2_io_dataIn; // @[LVT_set.scala 21:18]
  wire [63:0] b2_io_dataOut; // @[LVT_set.scala 21:18]
  wire  b3_clock; // @[LVT_set.scala 22:18]
  wire  b3_io_wenable; // @[LVT_set.scala 22:18]
  wire  b3_io_renable; // @[LVT_set.scala 22:18]
  wire [5:0] b3_io_raddr; // @[LVT_set.scala 22:18]
  wire [5:0] b3_io_waddr; // @[LVT_set.scala 22:18]
  wire [63:0] b3_io_dataIn; // @[LVT_set.scala 22:18]
  wire [63:0] b3_io_dataOut; // @[LVT_set.scala 22:18]
  ReadWriteSmem b1 ( // @[LVT_set.scala 20:18]
    .clock(b1_clock),
    .io_wenable(b1_io_wenable),
    .io_renable(b1_io_renable),
    .io_raddr(b1_io_raddr),
    .io_waddr(b1_io_waddr),
    .io_dataIn(b1_io_dataIn),
    .io_dataOut(b1_io_dataOut)
  );
  ReadWriteSmem b2 ( // @[LVT_set.scala 21:18]
    .clock(b2_clock),
    .io_wenable(b2_io_wenable),
    .io_renable(b2_io_renable),
    .io_raddr(b2_io_raddr),
    .io_waddr(b2_io_waddr),
    .io_dataIn(b2_io_dataIn),
    .io_dataOut(b2_io_dataOut)
  );
  ReadWriteSmem b3 ( // @[LVT_set.scala 22:18]
    .clock(b3_clock),
    .io_wenable(b3_io_wenable),
    .io_renable(b3_io_renable),
    .io_raddr(b3_io_raddr),
    .io_waddr(b3_io_waddr),
    .io_dataIn(b3_io_dataIn),
    .io_dataOut(b3_io_dataOut)
  );
  assign io_r1data = b1_io_dataOut; // @[LVT_set.scala 35:13]
  assign io_r2data = b2_io_dataOut; // @[LVT_set.scala 36:13]
  assign io_r3data = b3_io_dataOut; // @[LVT_set.scala 37:13]
  assign b1_clock = clock;
  assign b1_io_wenable = io_wenable; // @[LVT_set.scala 24:17]
  assign b1_io_renable = io_r1enable; // @[LVT_set.scala 31:17]
  assign b1_io_raddr = io_r1addr; // @[LVT_set.scala 39:15]
  assign b1_io_waddr = io_waddr; // @[LVT_set.scala 43:15]
  assign b1_io_dataIn = io_wdata; // @[LVT_set.scala 27:16]
  assign b2_clock = clock;
  assign b2_io_wenable = io_wenable; // @[LVT_set.scala 25:17]
  assign b2_io_renable = io_r2enable; // @[LVT_set.scala 32:17]
  assign b2_io_raddr = io_r2addr; // @[LVT_set.scala 40:15]
  assign b2_io_waddr = io_waddr; // @[LVT_set.scala 44:15]
  assign b2_io_dataIn = io_wdata; // @[LVT_set.scala 28:16]
  assign b3_clock = clock;
  assign b3_io_wenable = io_wenable; // @[LVT_set.scala 26:17]
  assign b3_io_renable = io_r3enable; // @[LVT_set.scala 33:17]
  assign b3_io_raddr = io_r3addr; // @[LVT_set.scala 41:15]
  assign b3_io_waddr = io_waddr; // @[LVT_set.scala 45:15]
  assign b3_io_dataIn = io_wdata; // @[LVT_set.scala 29:16]
endmodule
module LVT_Mem(
  input         clock,
  input         reset,
  input  [5:0]  io_R1_addr,
  output [63:0] io_R1_data,
  input         io_R1_en,
  input  [5:0]  io_R2_addr,
  output [63:0] io_R2_data,
  input         io_R2_en,
  input  [5:0]  io_R3_addr,
  output [63:0] io_R3_data,
  input         io_R3_en,
  input  [5:0]  io_W1_addr,
  input  [63:0] io_W1_data,
  input         io_W1_en,
  input  [5:0]  io_W2_addr,
  input  [63:0] io_W2_data,
  input         io_W2_en,
  input  [5:0]  io_W3_addr,
  input  [63:0] io_W3_data,
  input         io_W3_en,
  input  [5:0]  io_W4_addr,
  input  [63:0] io_W4_data,
  input         io_W4_en
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] LVT [0:63]; // @[LVT_Mem.scala 32:16]
  wire  LVT_r1_sel_reg_MPORT_en; // @[LVT_Mem.scala 32:16]
  wire [5:0] LVT_r1_sel_reg_MPORT_addr; // @[LVT_Mem.scala 32:16]
  wire [1:0] LVT_r1_sel_reg_MPORT_data; // @[LVT_Mem.scala 32:16]
  wire  LVT_r2_sel_reg_MPORT_en; // @[LVT_Mem.scala 32:16]
  wire [5:0] LVT_r2_sel_reg_MPORT_addr; // @[LVT_Mem.scala 32:16]
  wire [1:0] LVT_r2_sel_reg_MPORT_data; // @[LVT_Mem.scala 32:16]
  wire  LVT_r3_sel_reg_MPORT_en; // @[LVT_Mem.scala 32:16]
  wire [5:0] LVT_r3_sel_reg_MPORT_addr; // @[LVT_Mem.scala 32:16]
  wire [1:0] LVT_r3_sel_reg_MPORT_data; // @[LVT_Mem.scala 32:16]
  wire [1:0] LVT_MPORT_data; // @[LVT_Mem.scala 32:16]
  wire [5:0] LVT_MPORT_addr; // @[LVT_Mem.scala 32:16]
  wire  LVT_MPORT_mask; // @[LVT_Mem.scala 32:16]
  wire  LVT_MPORT_en; // @[LVT_Mem.scala 32:16]
  wire [1:0] LVT_MPORT_1_data; // @[LVT_Mem.scala 32:16]
  wire [5:0] LVT_MPORT_1_addr; // @[LVT_Mem.scala 32:16]
  wire  LVT_MPORT_1_mask; // @[LVT_Mem.scala 32:16]
  wire  LVT_MPORT_1_en; // @[LVT_Mem.scala 32:16]
  wire [1:0] LVT_MPORT_2_data; // @[LVT_Mem.scala 32:16]
  wire [5:0] LVT_MPORT_2_addr; // @[LVT_Mem.scala 32:16]
  wire  LVT_MPORT_2_mask; // @[LVT_Mem.scala 32:16]
  wire  LVT_MPORT_2_en; // @[LVT_Mem.scala 32:16]
  wire [1:0] LVT_MPORT_3_data; // @[LVT_Mem.scala 32:16]
  wire [5:0] LVT_MPORT_3_addr; // @[LVT_Mem.scala 32:16]
  wire  LVT_MPORT_3_mask; // @[LVT_Mem.scala 32:16]
  wire  LVT_MPORT_3_en; // @[LVT_Mem.scala 32:16]
  wire  s1_clock; // @[LVT_Mem.scala 35:18]
  wire  s1_io_wenable; // @[LVT_Mem.scala 35:18]
  wire  s1_io_r1enable; // @[LVT_Mem.scala 35:18]
  wire  s1_io_r2enable; // @[LVT_Mem.scala 35:18]
  wire  s1_io_r3enable; // @[LVT_Mem.scala 35:18]
  wire [5:0] s1_io_r1addr; // @[LVT_Mem.scala 35:18]
  wire [5:0] s1_io_r2addr; // @[LVT_Mem.scala 35:18]
  wire [5:0] s1_io_r3addr; // @[LVT_Mem.scala 35:18]
  wire [5:0] s1_io_waddr; // @[LVT_Mem.scala 35:18]
  wire [63:0] s1_io_wdata; // @[LVT_Mem.scala 35:18]
  wire [63:0] s1_io_r1data; // @[LVT_Mem.scala 35:18]
  wire [63:0] s1_io_r2data; // @[LVT_Mem.scala 35:18]
  wire [63:0] s1_io_r3data; // @[LVT_Mem.scala 35:18]
  wire  s2_clock; // @[LVT_Mem.scala 36:18]
  wire  s2_io_wenable; // @[LVT_Mem.scala 36:18]
  wire  s2_io_r1enable; // @[LVT_Mem.scala 36:18]
  wire  s2_io_r2enable; // @[LVT_Mem.scala 36:18]
  wire  s2_io_r3enable; // @[LVT_Mem.scala 36:18]
  wire [5:0] s2_io_r1addr; // @[LVT_Mem.scala 36:18]
  wire [5:0] s2_io_r2addr; // @[LVT_Mem.scala 36:18]
  wire [5:0] s2_io_r3addr; // @[LVT_Mem.scala 36:18]
  wire [5:0] s2_io_waddr; // @[LVT_Mem.scala 36:18]
  wire [63:0] s2_io_wdata; // @[LVT_Mem.scala 36:18]
  wire [63:0] s2_io_r1data; // @[LVT_Mem.scala 36:18]
  wire [63:0] s2_io_r2data; // @[LVT_Mem.scala 36:18]
  wire [63:0] s2_io_r3data; // @[LVT_Mem.scala 36:18]
  wire  s3_clock; // @[LVT_Mem.scala 37:18]
  wire  s3_io_wenable; // @[LVT_Mem.scala 37:18]
  wire  s3_io_r1enable; // @[LVT_Mem.scala 37:18]
  wire  s3_io_r2enable; // @[LVT_Mem.scala 37:18]
  wire  s3_io_r3enable; // @[LVT_Mem.scala 37:18]
  wire [5:0] s3_io_r1addr; // @[LVT_Mem.scala 37:18]
  wire [5:0] s3_io_r2addr; // @[LVT_Mem.scala 37:18]
  wire [5:0] s3_io_r3addr; // @[LVT_Mem.scala 37:18]
  wire [5:0] s3_io_waddr; // @[LVT_Mem.scala 37:18]
  wire [63:0] s3_io_wdata; // @[LVT_Mem.scala 37:18]
  wire [63:0] s3_io_r1data; // @[LVT_Mem.scala 37:18]
  wire [63:0] s3_io_r2data; // @[LVT_Mem.scala 37:18]
  wire [63:0] s3_io_r3data; // @[LVT_Mem.scala 37:18]
  wire  s4_clock; // @[LVT_Mem.scala 38:18]
  wire  s4_io_wenable; // @[LVT_Mem.scala 38:18]
  wire  s4_io_r1enable; // @[LVT_Mem.scala 38:18]
  wire  s4_io_r2enable; // @[LVT_Mem.scala 38:18]
  wire  s4_io_r3enable; // @[LVT_Mem.scala 38:18]
  wire [5:0] s4_io_r1addr; // @[LVT_Mem.scala 38:18]
  wire [5:0] s4_io_r2addr; // @[LVT_Mem.scala 38:18]
  wire [5:0] s4_io_r3addr; // @[LVT_Mem.scala 38:18]
  wire [5:0] s4_io_waddr; // @[LVT_Mem.scala 38:18]
  wire [63:0] s4_io_wdata; // @[LVT_Mem.scala 38:18]
  wire [63:0] s4_io_r1data; // @[LVT_Mem.scala 38:18]
  wire [63:0] s4_io_r2data; // @[LVT_Mem.scala 38:18]
  wire [63:0] s4_io_r3data; // @[LVT_Mem.scala 38:18]
  reg [1:0] r1_sel_reg; // @[LVT_Mem.scala 69:27]
  reg [1:0] r2_sel_reg; // @[LVT_Mem.scala 70:27]
  reg [1:0] r3_sel_reg; // @[LVT_Mem.scala 71:27]
  wire  _io_R1_data_T = r1_sel_reg == 2'h0; // @[LVT_Mem.scala 110:45]
  wire  _io_R1_data_T_1 = r1_sel_reg == 2'h1; // @[LVT_Mem.scala 110:79]
  wire  _io_R1_data_T_2 = r1_sel_reg == 2'h2; // @[LVT_Mem.scala 110:113]
  wire  _io_R1_data_T_3 = r1_sel_reg == 2'h3; // @[LVT_Mem.scala 110:147]
  wire [63:0] _io_R1_data_T_4 = _io_R1_data_T_3 ? s4_io_r1data : 64'h0; // @[Mux.scala 101:16]
  wire [63:0] _io_R1_data_T_5 = _io_R1_data_T_2 ? s3_io_r1data : _io_R1_data_T_4; // @[Mux.scala 101:16]
  wire [63:0] _io_R1_data_T_6 = _io_R1_data_T_1 ? s2_io_r1data : _io_R1_data_T_5; // @[Mux.scala 101:16]
  wire  _io_R2_data_T = r2_sel_reg == 2'h0; // @[LVT_Mem.scala 111:45]
  wire  _io_R2_data_T_1 = r2_sel_reg == 2'h1; // @[LVT_Mem.scala 111:79]
  wire  _io_R2_data_T_2 = r2_sel_reg == 2'h2; // @[LVT_Mem.scala 111:113]
  wire  _io_R2_data_T_3 = r2_sel_reg == 2'h3; // @[LVT_Mem.scala 111:147]
  wire [63:0] _io_R2_data_T_4 = _io_R2_data_T_3 ? s4_io_r2data : 64'h0; // @[Mux.scala 101:16]
  wire [63:0] _io_R2_data_T_5 = _io_R2_data_T_2 ? s3_io_r2data : _io_R2_data_T_4; // @[Mux.scala 101:16]
  wire [63:0] _io_R2_data_T_6 = _io_R2_data_T_1 ? s2_io_r2data : _io_R2_data_T_5; // @[Mux.scala 101:16]
  wire  _io_R3_data_T = r3_sel_reg == 2'h0; // @[LVT_Mem.scala 112:45]
  wire  _io_R3_data_T_1 = r3_sel_reg == 2'h1; // @[LVT_Mem.scala 112:79]
  wire  _io_R3_data_T_2 = r3_sel_reg == 2'h2; // @[LVT_Mem.scala 112:113]
  wire  _io_R3_data_T_3 = r3_sel_reg == 2'h3; // @[LVT_Mem.scala 112:147]
  wire [63:0] _io_R3_data_T_4 = _io_R3_data_T_3 ? s4_io_r3data : 64'h0; // @[Mux.scala 101:16]
  wire [63:0] _io_R3_data_T_5 = _io_R3_data_T_2 ? s3_io_r3data : _io_R3_data_T_4; // @[Mux.scala 101:16]
  wire [63:0] _io_R3_data_T_6 = _io_R3_data_T_1 ? s2_io_r3data : _io_R3_data_T_5; // @[Mux.scala 101:16]
  LVT_set s1 ( // @[LVT_Mem.scala 35:18]
    .clock(s1_clock),
    .io_wenable(s1_io_wenable),
    .io_r1enable(s1_io_r1enable),
    .io_r2enable(s1_io_r2enable),
    .io_r3enable(s1_io_r3enable),
    .io_r1addr(s1_io_r1addr),
    .io_r2addr(s1_io_r2addr),
    .io_r3addr(s1_io_r3addr),
    .io_waddr(s1_io_waddr),
    .io_wdata(s1_io_wdata),
    .io_r1data(s1_io_r1data),
    .io_r2data(s1_io_r2data),
    .io_r3data(s1_io_r3data)
  );
  LVT_set s2 ( // @[LVT_Mem.scala 36:18]
    .clock(s2_clock),
    .io_wenable(s2_io_wenable),
    .io_r1enable(s2_io_r1enable),
    .io_r2enable(s2_io_r2enable),
    .io_r3enable(s2_io_r3enable),
    .io_r1addr(s2_io_r1addr),
    .io_r2addr(s2_io_r2addr),
    .io_r3addr(s2_io_r3addr),
    .io_waddr(s2_io_waddr),
    .io_wdata(s2_io_wdata),
    .io_r1data(s2_io_r1data),
    .io_r2data(s2_io_r2data),
    .io_r3data(s2_io_r3data)
  );
  LVT_set s3 ( // @[LVT_Mem.scala 37:18]
    .clock(s3_clock),
    .io_wenable(s3_io_wenable),
    .io_r1enable(s3_io_r1enable),
    .io_r2enable(s3_io_r2enable),
    .io_r3enable(s3_io_r3enable),
    .io_r1addr(s3_io_r1addr),
    .io_r2addr(s3_io_r2addr),
    .io_r3addr(s3_io_r3addr),
    .io_waddr(s3_io_waddr),
    .io_wdata(s3_io_wdata),
    .io_r1data(s3_io_r1data),
    .io_r2data(s3_io_r2data),
    .io_r3data(s3_io_r3data)
  );
  LVT_set s4 ( // @[LVT_Mem.scala 38:18]
    .clock(s4_clock),
    .io_wenable(s4_io_wenable),
    .io_r1enable(s4_io_r1enable),
    .io_r2enable(s4_io_r2enable),
    .io_r3enable(s4_io_r3enable),
    .io_r1addr(s4_io_r1addr),
    .io_r2addr(s4_io_r2addr),
    .io_r3addr(s4_io_r3addr),
    .io_waddr(s4_io_waddr),
    .io_wdata(s4_io_wdata),
    .io_r1data(s4_io_r1data),
    .io_r2data(s4_io_r2data),
    .io_r3data(s4_io_r3data)
  );
  assign LVT_r1_sel_reg_MPORT_en = 1'h1;
  assign LVT_r1_sel_reg_MPORT_addr = io_R1_addr;
  assign LVT_r1_sel_reg_MPORT_data = LVT[LVT_r1_sel_reg_MPORT_addr]; // @[LVT_Mem.scala 32:16]
  assign LVT_r2_sel_reg_MPORT_en = 1'h1;
  assign LVT_r2_sel_reg_MPORT_addr = io_R2_addr;
  assign LVT_r2_sel_reg_MPORT_data = LVT[LVT_r2_sel_reg_MPORT_addr]; // @[LVT_Mem.scala 32:16]
  assign LVT_r3_sel_reg_MPORT_en = 1'h1;
  assign LVT_r3_sel_reg_MPORT_addr = io_R3_addr;
  assign LVT_r3_sel_reg_MPORT_data = LVT[LVT_r3_sel_reg_MPORT_addr]; // @[LVT_Mem.scala 32:16]
  assign LVT_MPORT_data = 2'h0;
  assign LVT_MPORT_addr = io_W1_addr;
  assign LVT_MPORT_mask = 1'h1;
  assign LVT_MPORT_en = io_W1_en;
  assign LVT_MPORT_1_data = 2'h1;
  assign LVT_MPORT_1_addr = io_W2_addr;
  assign LVT_MPORT_1_mask = 1'h1;
  assign LVT_MPORT_1_en = io_W2_en;
  assign LVT_MPORT_2_data = 2'h2;
  assign LVT_MPORT_2_addr = io_W3_addr;
  assign LVT_MPORT_2_mask = 1'h1;
  assign LVT_MPORT_2_en = io_W3_en;
  assign LVT_MPORT_3_data = 2'h3;
  assign LVT_MPORT_3_addr = io_W4_addr;
  assign LVT_MPORT_3_mask = 1'h1;
  assign LVT_MPORT_3_en = io_W4_en;
  assign io_R1_data = _io_R1_data_T ? s1_io_r1data : _io_R1_data_T_6; // @[Mux.scala 101:16]
  assign io_R2_data = _io_R2_data_T ? s1_io_r2data : _io_R2_data_T_6; // @[Mux.scala 101:16]
  assign io_R3_data = _io_R3_data_T ? s1_io_r3data : _io_R3_data_T_6; // @[Mux.scala 101:16]
  assign s1_clock = clock;
  assign s1_io_wenable = io_W1_en; // @[LVT_Mem.scala 55:17]
  assign s1_io_r1enable = io_R1_en; // @[LVT_Mem.scala 93:18]
  assign s1_io_r2enable = io_R2_en; // @[LVT_Mem.scala 98:18]
  assign s1_io_r3enable = io_R3_en; // @[LVT_Mem.scala 103:18]
  assign s1_io_r1addr = io_R1_addr; // @[LVT_Mem.scala 78:16]
  assign s1_io_r2addr = io_R2_addr; // @[LVT_Mem.scala 83:16]
  assign s1_io_r3addr = io_R3_addr; // @[LVT_Mem.scala 88:16]
  assign s1_io_waddr = io_W1_addr; // @[LVT_Mem.scala 63:15]
  assign s1_io_wdata = io_W1_data; // @[LVT_Mem.scala 59:15]
  assign s2_clock = clock;
  assign s2_io_wenable = io_W2_en; // @[LVT_Mem.scala 56:17]
  assign s2_io_r1enable = io_R1_en; // @[LVT_Mem.scala 94:18]
  assign s2_io_r2enable = io_R2_en; // @[LVT_Mem.scala 99:18]
  assign s2_io_r3enable = io_R3_en; // @[LVT_Mem.scala 104:18]
  assign s2_io_r1addr = io_R1_addr; // @[LVT_Mem.scala 79:16]
  assign s2_io_r2addr = io_R2_addr; // @[LVT_Mem.scala 84:16]
  assign s2_io_r3addr = io_R3_addr; // @[LVT_Mem.scala 89:16]
  assign s2_io_waddr = io_W2_addr; // @[LVT_Mem.scala 64:15]
  assign s2_io_wdata = io_W2_data; // @[LVT_Mem.scala 60:15]
  assign s3_clock = clock;
  assign s3_io_wenable = io_W3_en; // @[LVT_Mem.scala 57:17]
  assign s3_io_r1enable = io_R1_en; // @[LVT_Mem.scala 95:18]
  assign s3_io_r2enable = io_R2_en; // @[LVT_Mem.scala 100:18]
  assign s3_io_r3enable = io_R3_en; // @[LVT_Mem.scala 105:18]
  assign s3_io_r1addr = io_R1_addr; // @[LVT_Mem.scala 80:16]
  assign s3_io_r2addr = io_R2_addr; // @[LVT_Mem.scala 85:16]
  assign s3_io_r3addr = io_R3_addr; // @[LVT_Mem.scala 90:16]
  assign s3_io_waddr = io_W3_addr; // @[LVT_Mem.scala 65:15]
  assign s3_io_wdata = io_W3_data; // @[LVT_Mem.scala 61:15]
  assign s4_clock = clock;
  assign s4_io_wenable = io_W4_en; // @[LVT_Mem.scala 58:17]
  assign s4_io_r1enable = io_R1_en; // @[LVT_Mem.scala 96:18]
  assign s4_io_r2enable = io_R2_en; // @[LVT_Mem.scala 101:18]
  assign s4_io_r3enable = io_R3_en; // @[LVT_Mem.scala 106:18]
  assign s4_io_r1addr = io_R1_addr; // @[LVT_Mem.scala 81:16]
  assign s4_io_r2addr = io_R2_addr; // @[LVT_Mem.scala 86:16]
  assign s4_io_r3addr = io_R3_addr; // @[LVT_Mem.scala 91:16]
  assign s4_io_waddr = io_W4_addr; // @[LVT_Mem.scala 66:15]
  assign s4_io_wdata = io_W4_data; // @[LVT_Mem.scala 62:15]
  always @(posedge clock) begin
    if (LVT_MPORT_en & LVT_MPORT_mask) begin
      LVT[LVT_MPORT_addr] <= LVT_MPORT_data; // @[LVT_Mem.scala 32:16]
    end
    if (LVT_MPORT_1_en & LVT_MPORT_1_mask) begin
      LVT[LVT_MPORT_1_addr] <= LVT_MPORT_1_data; // @[LVT_Mem.scala 32:16]
    end
    if (LVT_MPORT_2_en & LVT_MPORT_2_mask) begin
      LVT[LVT_MPORT_2_addr] <= LVT_MPORT_2_data; // @[LVT_Mem.scala 32:16]
    end
    if (LVT_MPORT_3_en & LVT_MPORT_3_mask) begin
      LVT[LVT_MPORT_3_addr] <= LVT_MPORT_3_data; // @[LVT_Mem.scala 32:16]
    end
    if (reset) begin // @[LVT_Mem.scala 69:27]
      r1_sel_reg <= 2'h0; // @[LVT_Mem.scala 69:27]
    end else begin
      r1_sel_reg <= LVT_r1_sel_reg_MPORT_data; // @[LVT_Mem.scala 73:14]
    end
    if (reset) begin // @[LVT_Mem.scala 70:27]
      r2_sel_reg <= 2'h0; // @[LVT_Mem.scala 70:27]
    end else begin
      r2_sel_reg <= LVT_r2_sel_reg_MPORT_data; // @[LVT_Mem.scala 74:14]
    end
    if (reset) begin // @[LVT_Mem.scala 71:27]
      r3_sel_reg <= 2'h0; // @[LVT_Mem.scala 71:27]
    end else begin
      r3_sel_reg <= LVT_r3_sel_reg_MPORT_data; // @[LVT_Mem.scala 75:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    LVT[initvar] = _RAND_0[1:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  r1_sel_reg = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  r2_sel_reg = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  r3_sel_reg = _RAND_3[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PRF(
  input         clock,
  input         reset,
  input  [5:0]  w1_addr,
  input  [63:0] w1_data,
  input         w1_en,
  input  [5:0]  w2_addr,
  input  [63:0] w2_data,
  input         w2_en,
  input  [5:0]  w3_addr,
  input  [63:0] w3_data,
  input         w3_en,
  input  [5:0]  w4_addr,
  input  [63:0] w4_data,
  input         w4_en,
  input         execRead_valid,
  input  [31:0] execRead_instruction,
  input  [3:0]  execRead_branchmask,
  input  [5:0]  execRead_rs1Addr,
  input  [5:0]  execRead_rs2Addr,
  input  [5:0]  execRead_robAddr,
  input  [5:0]  execRead_prfDest,
  output        toExec_valid,
  output [31:0] toExec_instruction,
  output [3:0]  toExec_branchmask,
  output [5:0]  toExec_rs1Addr,
  output [63:0] toExec_rs1Data,
  output [5:0]  toExec_rs2Addr,
  output [63:0] toExec_rs2Data,
  output [5:0]  toExec_robAddr,
  output [5:0]  toExec_prfDest,
  input         fromStore_valid,
  input  [5:0]  fromStore_rs2Addr,
  output        toStore_valid,
  output [63:0] toStore_rs2Data,
  input         branchCheck_pass,
  input  [3:0]  branchCheck_branchmask,
  input         branchCheck_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  prf_clock; // @[PRF.scala 72:19]
  wire  prf_reset; // @[PRF.scala 72:19]
  wire [5:0] prf_io_R1_addr; // @[PRF.scala 72:19]
  wire [63:0] prf_io_R1_data; // @[PRF.scala 72:19]
  wire  prf_io_R1_en; // @[PRF.scala 72:19]
  wire [5:0] prf_io_R2_addr; // @[PRF.scala 72:19]
  wire [63:0] prf_io_R2_data; // @[PRF.scala 72:19]
  wire  prf_io_R2_en; // @[PRF.scala 72:19]
  wire [5:0] prf_io_R3_addr; // @[PRF.scala 72:19]
  wire [63:0] prf_io_R3_data; // @[PRF.scala 72:19]
  wire  prf_io_R3_en; // @[PRF.scala 72:19]
  wire [5:0] prf_io_W1_addr; // @[PRF.scala 72:19]
  wire [63:0] prf_io_W1_data; // @[PRF.scala 72:19]
  wire  prf_io_W1_en; // @[PRF.scala 72:19]
  wire [5:0] prf_io_W2_addr; // @[PRF.scala 72:19]
  wire [63:0] prf_io_W2_data; // @[PRF.scala 72:19]
  wire  prf_io_W2_en; // @[PRF.scala 72:19]
  wire [5:0] prf_io_W3_addr; // @[PRF.scala 72:19]
  wire [63:0] prf_io_W3_data; // @[PRF.scala 72:19]
  wire  prf_io_W3_en; // @[PRF.scala 72:19]
  wire [5:0] prf_io_W4_addr; // @[PRF.scala 72:19]
  wire [63:0] prf_io_W4_data; // @[PRF.scala 72:19]
  wire  prf_io_W4_en; // @[PRF.scala 72:19]
  reg [5:0] toExec_robAddr_REG; // @[PRF.scala 81:28]
  reg [5:0] toExec_rs1Addr_REG; // @[PRF.scala 82:28]
  reg [5:0] toExec_rs2Addr_REG; // @[PRF.scala 83:28]
  reg [31:0] toExec_instruction_REG; // @[PRF.scala 84:32]
  reg [5:0] toExec_prfDest_REG; // @[PRF.scala 86:28]
  reg  toExec_valid_; // @[PRF.scala 103:29]
  reg [3:0] toExec_mask; // @[PRF.scala 106:28]
  wire [3:0] _T = branchCheck_branchmask & execRead_branchmask; // @[PRF.scala 114:36]
  wire [3:0] _toExec_mask_T = branchCheck_branchmask ^ execRead_branchmask; // @[PRF.scala 115:47]
  reg  toStore_valid_REG_1; // @[PRF.scala 139:27]
  LVT_Mem prf ( // @[PRF.scala 72:19]
    .clock(prf_clock),
    .reset(prf_reset),
    .io_R1_addr(prf_io_R1_addr),
    .io_R1_data(prf_io_R1_data),
    .io_R1_en(prf_io_R1_en),
    .io_R2_addr(prf_io_R2_addr),
    .io_R2_data(prf_io_R2_data),
    .io_R2_en(prf_io_R2_en),
    .io_R3_addr(prf_io_R3_addr),
    .io_R3_data(prf_io_R3_data),
    .io_R3_en(prf_io_R3_en),
    .io_W1_addr(prf_io_W1_addr),
    .io_W1_data(prf_io_W1_data),
    .io_W1_en(prf_io_W1_en),
    .io_W2_addr(prf_io_W2_addr),
    .io_W2_data(prf_io_W2_data),
    .io_W2_en(prf_io_W2_en),
    .io_W3_addr(prf_io_W3_addr),
    .io_W3_data(prf_io_W3_data),
    .io_W3_en(prf_io_W3_en),
    .io_W4_addr(prf_io_W4_addr),
    .io_W4_data(prf_io_W4_data),
    .io_W4_en(prf_io_W4_en)
  );
  assign toExec_valid = toExec_valid_; // @[PRF.scala 135:16]
  assign toExec_instruction = toExec_instruction_REG; // @[PRF.scala 84:22]
  assign toExec_branchmask = toExec_mask; // @[PRF.scala 136:21]
  assign toExec_rs1Addr = toExec_rs1Addr_REG; // @[PRF.scala 82:18]
  assign toExec_rs1Data = prf_io_R1_data; // @[PRF.scala 92:18]
  assign toExec_rs2Addr = toExec_rs2Addr_REG; // @[PRF.scala 83:18]
  assign toExec_rs2Data = prf_io_R2_data; // @[PRF.scala 96:18]
  assign toExec_robAddr = toExec_robAddr_REG; // @[PRF.scala 81:18]
  assign toExec_prfDest = toExec_prfDest_REG; // @[PRF.scala 86:18]
  assign toStore_valid = toStore_valid_REG_1; // @[PRF.scala 139:17]
  assign toStore_rs2Data = prf_io_R3_data; // @[PRF.scala 100:19]
  assign prf_clock = clock;
  assign prf_reset = reset;
  assign prf_io_R1_addr = execRead_rs1Addr; // @[PRF.scala 91:18]
  assign prf_io_R1_en = execRead_valid; // @[PRF.scala 90:16]
  assign prf_io_R2_addr = execRead_rs2Addr; // @[PRF.scala 95:18]
  assign prf_io_R2_en = execRead_valid; // @[PRF.scala 94:16]
  assign prf_io_R3_addr = fromStore_rs2Addr; // @[PRF.scala 99:18]
  assign prf_io_R3_en = fromStore_valid; // @[PRF.scala 98:16]
  assign prf_io_W1_addr = w1_addr; // @[PRF.scala 75:13]
  assign prf_io_W1_data = w1_data; // @[PRF.scala 75:13]
  assign prf_io_W1_en = w1_en; // @[PRF.scala 75:13]
  assign prf_io_W2_addr = w2_addr; // @[PRF.scala 76:13]
  assign prf_io_W2_data = w2_data; // @[PRF.scala 76:13]
  assign prf_io_W2_en = w2_en; // @[PRF.scala 76:13]
  assign prf_io_W3_addr = w3_addr; // @[PRF.scala 77:13]
  assign prf_io_W3_data = w3_data; // @[PRF.scala 77:13]
  assign prf_io_W3_en = w3_en; // @[PRF.scala 77:13]
  assign prf_io_W4_addr = w4_addr; // @[PRF.scala 78:13]
  assign prf_io_W4_data = w4_data; // @[PRF.scala 78:13]
  assign prf_io_W4_en = w4_en; // @[PRF.scala 78:13]
  always @(posedge clock) begin
    toExec_robAddr_REG <= execRead_robAddr; // @[PRF.scala 81:28]
    toExec_rs1Addr_REG <= execRead_rs1Addr; // @[PRF.scala 82:28]
    toExec_rs2Addr_REG <= execRead_rs2Addr; // @[PRF.scala 83:28]
    toExec_instruction_REG <= execRead_instruction; // @[PRF.scala 84:32]
    toExec_prfDest_REG <= execRead_prfDest; // @[PRF.scala 86:28]
    if (reset) begin // @[PRF.scala 103:29]
      toExec_valid_ <= 1'h0; // @[PRF.scala 103:29]
    end else if (branchCheck_valid) begin // @[PRF.scala 109:27]
      if (branchCheck_pass) begin // @[PRF.scala 111:28]
        toExec_valid_ <= execRead_valid; // @[PRF.scala 112:20]
      end else begin
        toExec_valid_ <= _T == 4'h0 & execRead_valid; // @[PRF.scala 121:20]
      end
    end else begin
      toExec_valid_ <= execRead_valid; // @[PRF.scala 128:18]
    end
    if (reset) begin // @[PRF.scala 106:28]
      toExec_mask <= 4'h0; // @[PRF.scala 106:28]
    end else if (branchCheck_valid) begin // @[PRF.scala 109:27]
      if (branchCheck_pass) begin // @[PRF.scala 111:28]
        if (|_T) begin // @[PRF.scala 114:64]
          toExec_mask <= _toExec_mask_T; // @[PRF.scala 115:21]
        end else begin
          toExec_mask <= execRead_branchmask; // @[PRF.scala 113:19]
        end
      end else begin
        toExec_mask <= execRead_branchmask; // @[PRF.scala 122:19]
      end
    end else begin
      toExec_mask <= execRead_branchmask; // @[PRF.scala 129:17]
    end
    if (reset) begin // @[PRF.scala 139:27]
      toStore_valid_REG_1 <= 1'h0; // @[PRF.scala 139:27]
    end else begin
      toStore_valid_REG_1 <= fromStore_valid; // @[PRF.scala 139:27]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  toExec_robAddr_REG = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  toExec_rs1Addr_REG = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  toExec_rs2Addr_REG = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  toExec_instruction_REG = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  toExec_prfDest_REG = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  toExec_valid_ = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  toExec_mask = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  toStore_valid_REG_1 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module core(
  input         clock,
  input         reset,
  output        iPort_AWID,
  output [31:0] iPort_AWADDR,
  output [7:0]  iPort_AWLEN,
  output [2:0]  iPort_AWSIZE,
  output [1:0]  iPort_AWBURST,
  output        iPort_AWLOCK,
  output [3:0]  iPort_AWCACHE,
  output [2:0]  iPort_AWPROT,
  output [3:0]  iPort_AWQOS,
  output        iPort_AWVALID,
  input         iPort_AWREADY,
  output [31:0] iPort_WDATA,
  output [3:0]  iPort_WSTRB,
  output        iPort_WLAST,
  output        iPort_WVALID,
  input         iPort_WREADY,
  input         iPort_BID,
  input  [1:0]  iPort_BRESP,
  input         iPort_BVALID,
  output        iPort_BREADY,
  output        iPort_ARID,
  output [31:0] iPort_ARADDR,
  output [7:0]  iPort_ARLEN,
  output [2:0]  iPort_ARSIZE,
  output [1:0]  iPort_ARBURST,
  output        iPort_ARLOCK,
  output [3:0]  iPort_ARCACHE,
  output [2:0]  iPort_ARPROT,
  output [3:0]  iPort_ARQOS,
  output        iPort_ARVALID,
  input         iPort_ARREADY,
  input         iPort_RID,
  input  [31:0] iPort_RDATA,
  input  [1:0]  iPort_RRESP,
  input         iPort_RLAST,
  input         iPort_RVALID,
  output        iPort_RREADY,
  output        dPort_AWID,
  output [31:0] dPort_AWADDR,
  output [7:0]  dPort_AWLEN,
  output [2:0]  dPort_AWSIZE,
  output [1:0]  dPort_AWBURST,
  output        dPort_AWLOCK,
  output [3:0]  dPort_AWCACHE,
  output [2:0]  dPort_AWPROT,
  output [3:0]  dPort_AWQOS,
  output        dPort_AWVALID,
  input         dPort_AWREADY,
  output [31:0] dPort_WDATA,
  output [3:0]  dPort_WSTRB,
  output        dPort_WLAST,
  output        dPort_WVALID,
  input         dPort_WREADY,
  input         dPort_BID,
  input  [1:0]  dPort_BRESP,
  input         dPort_BVALID,
  output        dPort_BREADY,
  output        dPort_ARID,
  output [31:0] dPort_ARADDR,
  output [7:0]  dPort_ARLEN,
  output [2:0]  dPort_ARSIZE,
  output [1:0]  dPort_ARBURST,
  output        dPort_ARLOCK,
  output [3:0]  dPort_ARCACHE,
  output [2:0]  dPort_ARPROT,
  output [3:0]  dPort_ARQOS,
  output        dPort_ARVALID,
  input         dPort_ARREADY,
  input         dPort_RID,
  input  [31:0] dPort_RDATA,
  input  [1:0]  dPort_RRESP,
  input         dPort_RLAST,
  input         dPort_RVALID,
  output        dPort_RREADY,
  output        peripheral_AWID,
  output [31:0] peripheral_AWADDR,
  output [7:0]  peripheral_AWLEN,
  output [2:0]  peripheral_AWSIZE,
  output [1:0]  peripheral_AWBURST,
  output        peripheral_AWLOCK,
  output [3:0]  peripheral_AWCACHE,
  output [2:0]  peripheral_AWPROT,
  output [3:0]  peripheral_AWQOS,
  output        peripheral_AWVALID,
  input         peripheral_AWREADY,
  output [31:0] peripheral_WDATA,
  output [3:0]  peripheral_WSTRB,
  output        peripheral_WLAST,
  output        peripheral_WVALID,
  input         peripheral_WREADY,
  input         peripheral_BID,
  input  [1:0]  peripheral_BRESP,
  input         peripheral_BVALID,
  output        peripheral_BREADY,
  output        peripheral_ARID,
  output [31:0] peripheral_ARADDR,
  output [7:0]  peripheral_ARLEN,
  output [2:0]  peripheral_ARSIZE,
  output [1:0]  peripheral_ARBURST,
  output        peripheral_ARLOCK,
  output [3:0]  peripheral_ARCACHE,
  output [2:0]  peripheral_ARPROT,
  output [3:0]  peripheral_ARQOS,
  output        peripheral_ARVALID,
  input         peripheral_ARREADY,
  input         peripheral_RID,
  input  [31:0] peripheral_RDATA,
  input  [1:0]  peripheral_RRESP,
  input         peripheral_RLAST,
  input         peripheral_RVALID,
  output        peripheral_RREADY,
  output        core_sample0,
  output        core_sample1,
  input         MTIP
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [95:0] _RAND_47;
  reg [95:0] _RAND_48;
  reg [95:0] _RAND_49;
  reg [95:0] _RAND_50;
  reg [95:0] _RAND_51;
  reg [95:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [95:0] _RAND_62;
  reg [95:0] _RAND_63;
  reg [95:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
`endif // RANDOMIZE_REG_INIT
  wire  icache_clock; // @[core.scala 19:22]
  wire  icache_reset; // @[core.scala 19:22]
  wire  icache_fromFetch_req_ready; // @[core.scala 19:22]
  wire  icache_fromFetch_req_valid; // @[core.scala 19:22]
  wire [63:0] icache_fromFetch_req_bits; // @[core.scala 19:22]
  wire  icache_fromFetch_resp_ready; // @[core.scala 19:22]
  wire  icache_fromFetch_resp_valid; // @[core.scala 19:22]
  wire [31:0] icache_fromFetch_resp_bits; // @[core.scala 19:22]
  wire  icache_updateAllCachelines_ready; // @[core.scala 19:22]
  wire  icache_updateAllCachelines_fired; // @[core.scala 19:22]
  wire  icache_cachelinesUpdatesResp_ready; // @[core.scala 19:22]
  wire  icache_cachelinesUpdatesResp_fired; // @[core.scala 19:22]
  wire [31:0] icache_lowLevelMem_ARADDR; // @[core.scala 19:22]
  wire  icache_lowLevelMem_ARVALID; // @[core.scala 19:22]
  wire  icache_lowLevelMem_ARREADY; // @[core.scala 19:22]
  wire [31:0] icache_lowLevelMem_RDATA; // @[core.scala 19:22]
  wire  icache_lowLevelMem_RLAST; // @[core.scala 19:22]
  wire  icache_lowLevelMem_RVALID; // @[core.scala 19:22]
  wire  icache_lowLevelMem_RREADY; // @[core.scala 19:22]
  wire  fetch_clock; // @[core.scala 28:21]
  wire  fetch_reset; // @[core.scala 28:21]
  wire  fetch_cache_req_ready; // @[core.scala 28:21]
  wire  fetch_cache_req_valid; // @[core.scala 28:21]
  wire [63:0] fetch_cache_req_bits; // @[core.scala 28:21]
  wire  fetch_cache_resp_ready; // @[core.scala 28:21]
  wire  fetch_cache_resp_valid; // @[core.scala 28:21]
  wire [31:0] fetch_cache_resp_bits; // @[core.scala 28:21]
  wire  fetch_toDecode_ready; // @[core.scala 28:21]
  wire  fetch_toDecode_fired; // @[core.scala 28:21]
  wire [63:0] fetch_toDecode_pc; // @[core.scala 28:21]
  wire [31:0] fetch_toDecode_instruction; // @[core.scala 28:21]
  wire  fetch_toDecode_expected_valid; // @[core.scala 28:21]
  wire [63:0] fetch_toDecode_expected_pc; // @[core.scala 28:21]
  wire  fetch_branchRes_fired; // @[core.scala 28:21]
  wire  fetch_branchRes_branchTaken; // @[core.scala 28:21]
  wire [63:0] fetch_branchRes_pc; // @[core.scala 28:21]
  wire [63:0] fetch_branchRes_pcAfterBrnach; // @[core.scala 28:21]
  wire  fetch_carryOutFence_ready; // @[core.scala 28:21]
  wire  fetch_carryOutFence_fired; // @[core.scala 28:21]
  wire  fetch_updateAllCachelines_ready; // @[core.scala 28:21]
  wire  fetch_updateAllCachelines_fired; // @[core.scala 28:21]
  wire  fetch_cachelinesUpdatesResp_ready; // @[core.scala 28:21]
  wire  fetch_cachelinesUpdatesResp_fired; // @[core.scala 28:21]
  wire  decode_clock; // @[core.scala 38:22]
  wire  decode_reset; // @[core.scala 38:22]
  wire  decode_fromFetch_ready; // @[core.scala 38:22]
  wire  decode_fromFetch_fired; // @[core.scala 38:22]
  wire [63:0] decode_fromFetch_pc; // @[core.scala 38:22]
  wire [31:0] decode_fromFetch_instruction; // @[core.scala 38:22]
  wire  decode_fromFetch_expected_valid; // @[core.scala 38:22]
  wire [63:0] decode_fromFetch_expected_pc; // @[core.scala 38:22]
  wire  decode_toExec_ready; // @[core.scala 38:22]
  wire  decode_toExec_fired; // @[core.scala 38:22]
  wire [31:0] decode_toExec_instruction; // @[core.scala 38:22]
  wire [63:0] decode_toExec_pc; // @[core.scala 38:22]
  wire [5:0] decode_toExec_PRFDest; // @[core.scala 38:22]
  wire [5:0] decode_toExec_rs1Addr; // @[core.scala 38:22]
  wire  decode_toExec_rs1Ready; // @[core.scala 38:22]
  wire [5:0] decode_toExec_rs2Addr; // @[core.scala 38:22]
  wire  decode_toExec_rs2Ready; // @[core.scala 38:22]
  wire [3:0] decode_toExec_branchMask; // @[core.scala 38:22]
  wire  decode_writeBackResult_fired; // @[core.scala 38:22]
  wire [31:0] decode_writeBackResult_instruction; // @[core.scala 38:22]
  wire [4:0] decode_writeBackResult_rdAddr; // @[core.scala 38:22]
  wire [5:0] decode_writeBackResult_PRFDest; // @[core.scala 38:22]
  wire [63:0] decode_writeBackResult_data; // @[core.scala 38:22]
  wire [5:0] decode_writeAddrPRF_exec1Addr; // @[core.scala 38:22]
  wire [5:0] decode_writeAddrPRF_exec2Addr; // @[core.scala 38:22]
  wire [5:0] decode_writeAddrPRF_exec3Addr; // @[core.scala 38:22]
  wire  decode_writeAddrPRF_exec1Valid; // @[core.scala 38:22]
  wire  decode_writeAddrPRF_exec2Valid; // @[core.scala 38:22]
  wire  decode_writeAddrPRF_exec3Valid; // @[core.scala 38:22]
  wire  decode_jumpAddrWrite_ready; // @[core.scala 38:22]
  wire  decode_jumpAddrWrite_fired; // @[core.scala 38:22]
  wire [5:0] decode_jumpAddrWrite_PRFDest; // @[core.scala 38:22]
  wire [63:0] decode_jumpAddrWrite_linkAddr; // @[core.scala 38:22]
  wire  decode_branchPCs_branchPCReady; // @[core.scala 38:22]
  wire [63:0] decode_branchPCs_branchPC; // @[core.scala 38:22]
  wire  decode_branchPCs_predictedPCReady; // @[core.scala 38:22]
  wire [63:0] decode_branchPCs_predictedPC; // @[core.scala 38:22]
  wire [3:0] decode_branchPCs_branchMask; // @[core.scala 38:22]
  wire  decode_branchEvalIn_fired; // @[core.scala 38:22]
  wire  decode_branchEvalIn_passFail; // @[core.scala 38:22]
  wire [3:0] decode_branchEvalIn_branchMask; // @[core.scala 38:22]
  wire [63:0] decode_branchEvalIn_targetPC; // @[core.scala 38:22]
  wire [63:0] decode_interruptedPC; // @[core.scala 38:22]
  wire  decode_canTakeInterrupt; // @[core.scala 38:22]
  wire  dataQueue_clock; // @[core.scala 52:25]
  wire  dataQueue_reset; // @[core.scala 52:25]
  wire  dataQueue_fromROB_readyNow; // @[core.scala 52:25]
  wire  dataQueue_fromBranch_passOrFail; // @[core.scala 52:25]
  wire [3:0] dataQueue_fromBranch_robAddr; // @[core.scala 52:25]
  wire  dataQueue_fromBranch_valid; // @[core.scala 52:25]
  wire  dataQueue_fromDecode_ready; // @[core.scala 52:25]
  wire  dataQueue_fromDecode_valid; // @[core.scala 52:25]
  wire [5:0] dataQueue_fromDecode_rs2Addr; // @[core.scala 52:25]
  wire [3:0] dataQueue_fromDecode_branchMask; // @[core.scala 52:25]
  wire  dataQueue_toPRF_valid; // @[core.scala 52:25]
  wire [5:0] dataQueue_toPRF_rs2Addr; // @[core.scala 52:25]
  wire  dataQueue_robMapUpdate_valid; // @[core.scala 52:25]
  wire [3:0] dataQueue_robMapUpdate_robAddr; // @[core.scala 52:25]
  wire  rob_clock; // @[core.scala 53:19]
  wire  rob_reset; // @[core.scala 53:19]
  wire  rob_allocate_ready; // @[core.scala 53:19]
  wire  rob_allocate_fired; // @[core.scala 53:19]
  wire [63:0] rob_allocate_pc; // @[core.scala 53:19]
  wire [31:0] rob_allocate_instruction; // @[core.scala 53:19]
  wire [5:0] rob_allocate_prfDest; // @[core.scala 53:19]
  wire [3:0] rob_allocate_robAddr; // @[core.scala 53:19]
  wire  rob_allocate_isReady; // @[core.scala 53:19]
  wire  rob_commit_ready; // @[core.scala 53:19]
  wire  rob_commit_fired; // @[core.scala 53:19]
  wire [5:0] rob_commit_prfDest; // @[core.scala 53:19]
  wire [31:0] rob_commit_instruction; // @[core.scala 53:19]
  wire  rob_commit_exceptionOccurred; // @[core.scala 53:19]
  wire [63:0] rob_commit_mtval; // @[core.scala 53:19]
  wire  rob_commit_isStore; // @[core.scala 53:19]
  wire  rob_commit_is_fence; // @[core.scala 53:19]
  wire [3:0] rob_commit_robAddr; // @[core.scala 53:19]
  wire  rob_branch_valid; // @[core.scala 53:19]
  wire  rob_branch_pass; // @[core.scala 53:19]
  wire [3:0] rob_branch_robAddr; // @[core.scala 53:19]
  wire [3:0] rob_execPorts_0_robAddr; // @[core.scala 53:19]
  wire [63:0] rob_execPorts_0_mtval; // @[core.scala 53:19]
  wire  rob_execPorts_0_valid; // @[core.scala 53:19]
  wire [3:0] rob_execPorts_1_robAddr; // @[core.scala 53:19]
  wire  rob_execPorts_1_valid; // @[core.scala 53:19]
  wire [3:0] rob_execPorts_2_robAddr; // @[core.scala 53:19]
  wire  rob_execPorts_2_valid; // @[core.scala 53:19]
  wire [3:0] rob_execPorts_3_robAddr; // @[core.scala 53:19]
  wire  rob_execPorts_3_valid; // @[core.scala 53:19]
  wire  scheduler_clock; // @[core.scala 54:25]
  wire  scheduler_reset; // @[core.scala 54:25]
  wire  scheduler_allocate_ready; // @[core.scala 54:25]
  wire  scheduler_allocate_fired; // @[core.scala 54:25]
  wire [31:0] scheduler_allocate_instruction; // @[core.scala 54:25]
  wire [3:0] scheduler_allocate_branchMask; // @[core.scala 54:25]
  wire  scheduler_allocate_rs1_ready; // @[core.scala 54:25]
  wire [5:0] scheduler_allocate_rs1_prfAddr; // @[core.scala 54:25]
  wire  scheduler_allocate_rs2_ready; // @[core.scala 54:25]
  wire [5:0] scheduler_allocate_rs2_prfAddr; // @[core.scala 54:25]
  wire [5:0] scheduler_allocate_prfDest; // @[core.scala 54:25]
  wire [3:0] scheduler_allocate_robAddr; // @[core.scala 54:25]
  wire  scheduler_release_ready; // @[core.scala 54:25]
  wire  scheduler_release_fired; // @[core.scala 54:25]
  wire [31:0] scheduler_release_instruction; // @[core.scala 54:25]
  wire [3:0] scheduler_release_branchMask; // @[core.scala 54:25]
  wire [5:0] scheduler_release_rs1prfAddr; // @[core.scala 54:25]
  wire [5:0] scheduler_release_rs2prfAddr; // @[core.scala 54:25]
  wire [5:0] scheduler_release_prfDest; // @[core.scala 54:25]
  wire [3:0] scheduler_release_robAddr; // @[core.scala 54:25]
  wire  scheduler_wakeUpExt_0_valid; // @[core.scala 54:25]
  wire [5:0] scheduler_wakeUpExt_0_prfAddr; // @[core.scala 54:25]
  wire  scheduler_wakeUpExt_1_valid; // @[core.scala 54:25]
  wire [5:0] scheduler_wakeUpExt_1_prfAddr; // @[core.scala 54:25]
  wire  scheduler_branchOps_valid; // @[core.scala 54:25]
  wire [3:0] scheduler_branchOps_branchMask; // @[core.scala 54:25]
  wire  scheduler_branchOps_passed; // @[core.scala 54:25]
  wire  scheduler_memoryReady; // @[core.scala 54:25]
  wire  scheduler_multuplyAndDivideReady; // @[core.scala 54:25]
  wire  scheduler_instrRetired_valid; // @[core.scala 54:25]
  wire [5:0] scheduler_instrRetired_prfAddr; // @[core.scala 54:25]
  wire  memAccess_clock; // @[core.scala 55:25]
  wire  memAccess_reset; // @[core.scala 55:25]
  wire [31:0] memAccess_peripheral_AWADDR; // @[core.scala 55:25]
  wire [7:0] memAccess_peripheral_AWLEN; // @[core.scala 55:25]
  wire [2:0] memAccess_peripheral_AWSIZE; // @[core.scala 55:25]
  wire  memAccess_peripheral_AWVALID; // @[core.scala 55:25]
  wire  memAccess_peripheral_AWREADY; // @[core.scala 55:25]
  wire [31:0] memAccess_peripheral_WDATA; // @[core.scala 55:25]
  wire [3:0] memAccess_peripheral_WSTRB; // @[core.scala 55:25]
  wire  memAccess_peripheral_WLAST; // @[core.scala 55:25]
  wire  memAccess_peripheral_WVALID; // @[core.scala 55:25]
  wire  memAccess_peripheral_WREADY; // @[core.scala 55:25]
  wire  memAccess_peripheral_BVALID; // @[core.scala 55:25]
  wire  memAccess_peripheral_BREADY; // @[core.scala 55:25]
  wire [31:0] memAccess_peripheral_ARADDR; // @[core.scala 55:25]
  wire [7:0] memAccess_peripheral_ARLEN; // @[core.scala 55:25]
  wire [2:0] memAccess_peripheral_ARSIZE; // @[core.scala 55:25]
  wire  memAccess_peripheral_ARVALID; // @[core.scala 55:25]
  wire  memAccess_peripheral_ARREADY; // @[core.scala 55:25]
  wire [31:0] memAccess_peripheral_RDATA; // @[core.scala 55:25]
  wire  memAccess_peripheral_RLAST; // @[core.scala 55:25]
  wire  memAccess_peripheral_RVALID; // @[core.scala 55:25]
  wire  memAccess_peripheral_RREADY; // @[core.scala 55:25]
  wire  memAccess_branchOps_valid; // @[core.scala 55:25]
  wire [3:0] memAccess_branchOps_branchMask; // @[core.scala 55:25]
  wire  memAccess_branchOps_passed; // @[core.scala 55:25]
  wire  memAccess_writeDataIn_valid; // @[core.scala 55:25]
  wire [63:0] memAccess_writeDataIn_data; // @[core.scala 55:25]
  wire  memAccess_responseOut_valid; // @[core.scala 55:25]
  wire [5:0] memAccess_responseOut_prfDest; // @[core.scala 55:25]
  wire [3:0] memAccess_responseOut_robAddr; // @[core.scala 55:25]
  wire [63:0] memAccess_responseOut_result; // @[core.scala 55:25]
  wire [31:0] memAccess_responseOut_instruction; // @[core.scala 55:25]
  wire  memAccess_request_valid; // @[core.scala 55:25]
  wire [31:0] memAccess_request_address; // @[core.scala 55:25]
  wire [31:0] memAccess_request_instruction; // @[core.scala 55:25]
  wire [3:0] memAccess_request_branchMask; // @[core.scala 55:25]
  wire [3:0] memAccess_request_robAddr; // @[core.scala 55:25]
  wire [5:0] memAccess_request_prfDest; // @[core.scala 55:25]
  wire [31:0] memAccess_dPort_AWADDR; // @[core.scala 55:25]
  wire [7:0] memAccess_dPort_AWLEN; // @[core.scala 55:25]
  wire [2:0] memAccess_dPort_AWSIZE; // @[core.scala 55:25]
  wire  memAccess_dPort_AWVALID; // @[core.scala 55:25]
  wire  memAccess_dPort_AWREADY; // @[core.scala 55:25]
  wire [31:0] memAccess_dPort_WDATA; // @[core.scala 55:25]
  wire [3:0] memAccess_dPort_WSTRB; // @[core.scala 55:25]
  wire  memAccess_dPort_WLAST; // @[core.scala 55:25]
  wire  memAccess_dPort_WVALID; // @[core.scala 55:25]
  wire  memAccess_dPort_WREADY; // @[core.scala 55:25]
  wire  memAccess_dPort_BVALID; // @[core.scala 55:25]
  wire  memAccess_dPort_BREADY; // @[core.scala 55:25]
  wire [31:0] memAccess_dPort_ARADDR; // @[core.scala 55:25]
  wire  memAccess_dPort_ARVALID; // @[core.scala 55:25]
  wire  memAccess_dPort_ARREADY; // @[core.scala 55:25]
  wire [31:0] memAccess_dPort_RDATA; // @[core.scala 55:25]
  wire  memAccess_dPort_RLAST; // @[core.scala 55:25]
  wire  memAccess_dPort_RVALID; // @[core.scala 55:25]
  wire  memAccess_dPort_RREADY; // @[core.scala 55:25]
  wire  memAccess_writeCommit_ready; // @[core.scala 55:25]
  wire  memAccess_writeCommit_fired; // @[core.scala 55:25]
  wire  memAccess_canAllocate; // @[core.scala 55:25]
  wire  memAccess_initiateFence; // @[core.scala 55:25]
  wire  memAccess_fenceInstructions_ready; // @[core.scala 55:25]
  wire  memAccess_fenceInstructions_fired; // @[core.scala 55:25]
  wire  prf_clock; // @[core.scala 119:19]
  wire  prf_reset; // @[core.scala 119:19]
  wire [5:0] prf_w1_addr; // @[core.scala 119:19]
  wire [63:0] prf_w1_data; // @[core.scala 119:19]
  wire  prf_w1_en; // @[core.scala 119:19]
  wire [5:0] prf_w2_addr; // @[core.scala 119:19]
  wire [63:0] prf_w2_data; // @[core.scala 119:19]
  wire  prf_w2_en; // @[core.scala 119:19]
  wire [5:0] prf_w3_addr; // @[core.scala 119:19]
  wire [63:0] prf_w3_data; // @[core.scala 119:19]
  wire  prf_w3_en; // @[core.scala 119:19]
  wire [5:0] prf_w4_addr; // @[core.scala 119:19]
  wire [63:0] prf_w4_data; // @[core.scala 119:19]
  wire  prf_w4_en; // @[core.scala 119:19]
  wire  prf_execRead_valid; // @[core.scala 119:19]
  wire [31:0] prf_execRead_instruction; // @[core.scala 119:19]
  wire [3:0] prf_execRead_branchmask; // @[core.scala 119:19]
  wire [5:0] prf_execRead_rs1Addr; // @[core.scala 119:19]
  wire [5:0] prf_execRead_rs2Addr; // @[core.scala 119:19]
  wire [5:0] prf_execRead_robAddr; // @[core.scala 119:19]
  wire [5:0] prf_execRead_prfDest; // @[core.scala 119:19]
  wire  prf_toExec_valid; // @[core.scala 119:19]
  wire [31:0] prf_toExec_instruction; // @[core.scala 119:19]
  wire [3:0] prf_toExec_branchmask; // @[core.scala 119:19]
  wire [5:0] prf_toExec_rs1Addr; // @[core.scala 119:19]
  wire [63:0] prf_toExec_rs1Data; // @[core.scala 119:19]
  wire [5:0] prf_toExec_rs2Addr; // @[core.scala 119:19]
  wire [63:0] prf_toExec_rs2Data; // @[core.scala 119:19]
  wire [5:0] prf_toExec_robAddr; // @[core.scala 119:19]
  wire [5:0] prf_toExec_prfDest; // @[core.scala 119:19]
  wire  prf_fromStore_valid; // @[core.scala 119:19]
  wire [5:0] prf_fromStore_rs2Addr; // @[core.scala 119:19]
  wire  prf_toStore_valid; // @[core.scala 119:19]
  wire [63:0] prf_toStore_rs2Data; // @[core.scala 119:19]
  wire  prf_branchCheck_pass; // @[core.scala 119:19]
  wire [3:0] prf_branchCheck_branchmask; // @[core.scala 119:19]
  wire  prf_branchCheck_valid; // @[core.scala 119:19]
  wire  _fetch_toDecode_fired_T_3 = ~decode_fromFetch_expected_valid | decode_fromFetch_expected_pc == fetch_toDecode_pc
    ; // @[core.scala 45:40]
  wire  instructionDecodedReady = 5'h3 == decode_toExec_instruction[6:2] | 5'h5 == decode_toExec_instruction[6:2] | 5'hd
     == decode_toExec_instruction[6:2]; // @[core.scala 77:125]
  wire [6:0] _scheduler_allocate_rs2_ready_T_1 = decode_toExec_instruction[6:0] & 7'h77; // @[core.scala 90:72]
  wire  _GEN_0 = instructionDecodedReady ? 1'h0 : decode_toExec_ready & rob_allocate_ready & scheduler_allocate_ready &
    (decode_toExec_instruction[6:4] != 3'h2 | dataQueue_fromDecode_ready); // @[core.scala 99:{33,60} 79:7]
  reg [3:0] branchEvals_branchMask; // @[core.scala 509:28]
  wire [3:0] _scheduler_allocate_branchMask_T = decode_toExec_branchMask ^ branchEvals_branchMask; // @[core.scala 101:62]
  reg  branchEvals_passed; // @[core.scala 509:28]
  wire  _T = ~branchEvals_passed; // @[core.scala 103:9]
  wire  _GEN_1 = ~branchEvals_passed ? 1'h0 : _GEN_0; // @[core.scala 103:28 104:30]
  wire  _GEN_2 = ~branchEvals_passed ? 1'h0 : decode_toExec_ready & rob_allocate_ready & scheduler_allocate_ready & (
    decode_toExec_instruction[6:4] != 3'h2 | dataQueue_fromDecode_ready); // @[core.scala 103:28 105:24 79:7]
  wire  _GEN_3 = ~branchEvals_passed ? 1'h0 : scheduler_allocate_fired & decode_toExec_instruction[6:4] == 3'h2; // @[core.scala 103:28 106:32 98:30]
  reg  branchEvals_valid; // @[core.scala 509:28]
  wire [5:0] wakeUps_0_prfAddr = scheduler_instrRetired_prfAddr; // @[core.scala 71:21 757:20]
  wire  _GEN_9 = decode_toExec_rs1Addr == wakeUps_0_prfAddr | decode_toExec_rs1Ready; // @[core.scala 112:{55,86} 88:32]
  wire  _GEN_10 = decode_toExec_rs2Addr == wakeUps_0_prfAddr | (7'h13 == _scheduler_allocate_rs2_ready_T_1 |
    decode_toExec_rs2Ready); // @[core.scala 113:{55,86} 90:32]
  wire  wakeUps_0_valid = scheduler_instrRetired_valid; // @[core.scala 71:21 758:18]
  wire  _GEN_11 = wakeUps_0_valid ? _GEN_9 : decode_toExec_rs1Ready; // @[core.scala 111:24 88:32]
  wire  _GEN_12 = wakeUps_0_valid ? _GEN_10 : 7'h13 == _scheduler_allocate_rs2_ready_T_1 | decode_toExec_rs2Ready; // @[core.scala 111:24 90:32]
  wire [5:0] wakeUps_1_prfAddr = memAccess_responseOut_prfDest; // @[core.scala 71:21 757:20]
  wire  _GEN_13 = decode_toExec_rs1Addr == wakeUps_1_prfAddr | _GEN_11; // @[core.scala 112:{55,86}]
  wire  _GEN_14 = decode_toExec_rs2Addr == wakeUps_1_prfAddr | _GEN_12; // @[core.scala 113:{55,86}]
  wire  _T_181 = |memAccess_responseOut_instruction[11:7]; // @[core.scala 752:77]
  wire  wakeUps_1_valid = memAccess_responseOut_valid & |memAccess_responseOut_instruction[11:7]; // @[core.scala 752:33]
  wire  _GEN_15 = wakeUps_1_valid ? _GEN_13 : _GEN_11; // @[core.scala 111:24]
  wire  _GEN_16 = wakeUps_1_valid ? _GEN_14 : _GEN_12; // @[core.scala 111:24]
  reg [5:0] extnMResponse_prfDest; // @[core.scala 211:30]
  wire  _GEN_17 = decode_toExec_rs1Addr == extnMResponse_prfDest | _GEN_15; // @[core.scala 112:{55,86}]
  wire  _GEN_18 = decode_toExec_rs2Addr == extnMResponse_prfDest | _GEN_16; // @[core.scala 113:{55,86}]
  reg  extnMResponse_valid; // @[core.scala 211:30]
  reg [31:0] extnResponseInstruction; // @[core.scala 350:36]
  wire  _T_184 = |extnResponseInstruction[11:7]; // @[core.scala 753:59]
  wire  wakeUps_2_valid = extnMResponse_valid & |extnResponseInstruction[11:7]; // @[core.scala 753:25]
  reg  mExtensionReady; // @[core.scala 117:32]
  wire [3:0] _scheduler_release_fired_T_2 = {scheduler_release_instruction[25],scheduler_release_instruction[6:4]}; // @[Cat.scala 33:92]
  wire  _scheduler_release_fired_T_5 = ~(_scheduler_release_fired_T_2 == 4'hb) | mExtensionReady; // @[core.scala 123:99]
  wire  _GEN_21 = scheduler_release_instruction[1:0] == 2'h0 ? 1'h0 : scheduler_release_fired; // @[core.scala 130:22 132:{57,78}]
  reg  addressGenerationInput_valid; // @[core.scala 140:39]
  reg [63:0] addressGenerationInput_rs1; // @[core.scala 140:39]
  reg [31:0] addressGenerationInput_instruction; // @[core.scala 140:39]
  reg [5:0] addressGenerationInput_prfDest; // @[core.scala 140:39]
  reg [3:0] addressGenerationInput_robAddr; // @[core.scala 140:39]
  reg [3:0] addressGenerationInput_branchMask; // @[core.scala 140:39]
  wire [3:0] _T_9 = prf_toExec_branchmask & branchEvals_branchMask; // @[core.scala 157:33]
  wire  _T_10 = |_T_9; // @[core.scala 157:57]
  wire [3:0] _addressGenerationInput_branchMask_T = prf_toExec_branchmask ^ branchEvals_branchMask; // @[core.scala 158:66]
  wire [3:0] _GEN_22 = |_T_9 ? _addressGenerationInput_branchMask_T : prf_toExec_branchmask; // @[core.scala 154:37 157:62 158:41]
  wire  _T_14 = _T & _T_10; // @[core.scala 160:28]
  wire [3:0] _GEN_24 = branchEvals_valid ? _GEN_22 : prf_toExec_branchmask; // @[core.scala 156:25 154:37]
  reg  memoryRequest_valid; // @[core.scala 163:30]
  reg [31:0] memoryRequest_address; // @[core.scala 163:30]
  reg [31:0] memoryRequest_instruction; // @[core.scala 163:30]
  reg [3:0] memoryRequest_branchMask; // @[core.scala 163:30]
  reg [3:0] memoryRequest_robAddr; // @[core.scala 163:30]
  reg [5:0] memoryRequest_prfDest; // @[core.scala 163:30]
  wire [51:0] _memoryRequest_address_T_2 = addressGenerationInput_instruction[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _memoryRequest_address_T_4 = {_memoryRequest_address_T_2,addressGenerationInput_instruction[31:20]}; // @[Cat.scala 33:92]
  wire [63:0] _memoryRequest_address_T_10 = {_memoryRequest_address_T_2,addressGenerationInput_instruction[31:25],
    addressGenerationInput_instruction[11:7]}; // @[Cat.scala 33:92]
  wire [1:0] _memoryRequest_address_T_13 = {addressGenerationInput_instruction[3],addressGenerationInput_instruction[5]}
    ; // @[Cat.scala 33:92]
  wire [63:0] _GEN_27 = 2'h1 == _memoryRequest_address_T_13 ? _memoryRequest_address_T_10 : _memoryRequest_address_T_4; // @[core.scala 164:{55,55}]
  wire [63:0] _GEN_28 = 2'h2 == _memoryRequest_address_T_13 ? 64'h0 : _GEN_27; // @[core.scala 164:{55,55}]
  wire [63:0] _GEN_29 = 2'h3 == _memoryRequest_address_T_13 ? 64'h0 : _GEN_28; // @[core.scala 164:{55,55}]
  wire [63:0] _memoryRequest_address_T_15 = addressGenerationInput_rs1 + _GEN_29; // @[core.scala 164:55]
  wire [3:0] _T_15 = addressGenerationInput_branchMask & branchEvals_branchMask; // @[core.scala 176:45]
  wire  _T_16 = |_T_15; // @[core.scala 176:69]
  wire [3:0] _memoryRequest_branchMask_T = addressGenerationInput_branchMask ^ branchEvals_branchMask; // @[core.scala 177:69]
  reg  singleCycleArithmeticRequest_valid; // @[core.scala 185:45]
  reg [63:0] singleCycleArithmeticRequest_rs1; // @[core.scala 185:45]
  reg [63:0] singleCycleArithmeticRequest_rs2; // @[core.scala 185:45]
  reg [31:0] singleCycleArithmeticRequest_instruction; // @[core.scala 185:45]
  reg [5:0] singleCycleArithmeticRequest_prfDest; // @[core.scala 185:45]
  reg [3:0] singleCycleArithmeticRequest_robAddr; // @[core.scala 185:45]
  reg [3:0] singleCycleArithmeticRequest_branchMask; // @[core.scala 185:45]
  reg  singleCycleArithmeticResponse_valid; // @[core.scala 195:46]
  reg [63:0] singleCycleArithmeticResponse_result; // @[core.scala 195:46]
  reg [5:0] singleCycleArithmeticResponse_prfDest; // @[core.scala 195:46]
  reg [3:0] singleCycleArithmeticResponse_robAddr; // @[core.scala 195:46]
  reg  extnMRequest_valid; // @[core.scala 202:29]
  reg [63:0] extnMRequest_rs1; // @[core.scala 202:29]
  reg [63:0] extnMRequest_rs2; // @[core.scala 202:29]
  reg [31:0] extnMRequest_instruction; // @[core.scala 202:29]
  reg [5:0] extnMRequest_prfDest; // @[core.scala 202:29]
  reg [3:0] extnMRequest_robAddr; // @[core.scala 202:29]
  reg [3:0] extnMRequest_branchMask; // @[core.scala 202:29]
  reg  extnMServicing_valid; // @[core.scala 204:31]
  reg [31:0] extnMServicing_instruction; // @[core.scala 204:31]
  reg [5:0] extnMServicing_prfDest; // @[core.scala 204:31]
  reg [3:0] extnMServicing_robAddr; // @[core.scala 204:31]
  reg [3:0] extnMServicing_branchMask; // @[core.scala 204:31]
  reg  extnMPartialServicing_valid; // @[core.scala 205:38]
  reg [31:0] extnMPartialServicing_instruction; // @[core.scala 205:38]
  reg [5:0] extnMPartialServicing_prfDest; // @[core.scala 205:38]
  reg [3:0] extnMPartialServicing_robAddr; // @[core.scala 205:38]
  reg [3:0] extnMPartialServicing_branchMask; // @[core.scala 205:38]
  reg [95:0] muls_0; // @[core.scala 206:17]
  reg [95:0] muls_1; // @[core.scala 206:17]
  reg [95:0] muls_2; // @[core.scala 206:17]
  reg [95:0] muls_3; // @[core.scala 206:17]
  reg [95:0] muls_4; // @[core.scala 206:17]
  reg [95:0] muls_5; // @[core.scala 206:17]
  reg [63:0] extnMResponse_result; // @[core.scala 211:30]
  reg [3:0] extnMResponse_robAddr; // @[core.scala 211:30]
  reg  division_request_valid; // @[core.scala 213:25]
  reg [63:0] division_request_rs1; // @[core.scala 213:25]
  reg [63:0] division_request_rs2; // @[core.scala 213:25]
  reg [31:0] division_request_instruction; // @[core.scala 213:25]
  reg [5:0] division_request_prfDest; // @[core.scala 213:25]
  reg [3:0] division_request_robAddr; // @[core.scala 213:25]
  reg [3:0] division_request_branchMask; // @[core.scala 213:25]
  reg [64:0] division_quotient; // @[core.scala 213:25]
  reg [64:0] division_remainder; // @[core.scala 213:25]
  reg [64:0] division_divisor; // @[core.scala 213:25]
  reg [6:0] division_counter; // @[core.scala 213:25]
  reg  fwdBuffers_0_valid; // @[core.scala 222:27]
  reg [5:0] fwdBuffers_0_prfDest; // @[core.scala 222:27]
  reg [63:0] fwdBuffers_0_result; // @[core.scala 222:27]
  reg  fwdBuffers_1_valid; // @[core.scala 222:27]
  reg [5:0] fwdBuffers_1_prfDest; // @[core.scala 222:27]
  reg [63:0] fwdBuffers_1_result; // @[core.scala 222:27]
  wire  _fwdFrom_0_valid_T_1 = |singleCycleArithmeticRequest_instruction[11:7]; // @[core.scala 231:109]
  wire  fwdFrom_0_valid = singleCycleArithmeticRequest_valid & |singleCycleArithmeticRequest_instruction[11:7]; // @[core.scala 231:58]
  wire  _addressGenerationInput_rs1_T_1 = |prf_toExec_instruction[19:15]; // @[core.scala 235:68]
  wire  _addressGenerationInput_rs1_T_3 = fwdFrom_0_valid & singleCycleArithmeticRequest_prfDest == prf_toExec_rs1Addr; // @[core.scala 236:34]
  wire  _addressGenerationInput_rs1_T_5 = fwdBuffers_0_valid & fwdBuffers_0_prfDest == prf_toExec_rs1Addr; // @[core.scala 236:34]
  wire  _addressGenerationInput_rs1_T_7 = fwdBuffers_1_valid & fwdBuffers_1_prfDest == prf_toExec_rs1Addr; // @[core.scala 236:34]
  wire [1:0] _arithmeticResult_arithmetic32_T_56 = {singleCycleArithmeticRequest_instruction[14],
    singleCycleArithmeticRequest_instruction[12]}; // @[Cat.scala 33:92]
  wire [31:0] _arithmeticResult_arithmetic32_T_36 = singleCycleArithmeticRequest_rs1[31:0]; // @[core.scala 251:69]
  wire [31:0] _arithmeticResult_arithmetic32_T_39 = $signed(_arithmeticResult_arithmetic32_T_36) >>>
    singleCycleArithmeticRequest_rs2[4:0]; // @[core.scala 251:90]
  wire [31:0] _arithmeticResult_arithmetic32_T_42 = _arithmeticResult_arithmetic32_T_39[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _arithmeticResult_arithmetic32_T_44 = {_arithmeticResult_arithmetic32_T_42,
    _arithmeticResult_arithmetic32_T_39}; // @[Cat.scala 33:92]
  wire [31:0] _arithmeticResult_arithmetic32_T_47 = singleCycleArithmeticRequest_rs1[31:0] >>
    singleCycleArithmeticRequest_rs2[4:0]; // @[core.scala 251:122]
  wire [31:0] _arithmeticResult_arithmetic32_T_50 = _arithmeticResult_arithmetic32_T_47[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _arithmeticResult_arithmetic32_T_52 = {_arithmeticResult_arithmetic32_T_50,
    _arithmeticResult_arithmetic32_T_47}; // @[Cat.scala 33:92]
  wire [63:0] _arithmeticResult_arithmetic32_T_53 = singleCycleArithmeticRequest_instruction[30] ?
    _arithmeticResult_arithmetic32_T_44 : _arithmeticResult_arithmetic32_T_52; // @[core.scala 251:20]
  wire [94:0] _GEN_250 = {{31'd0}, singleCycleArithmeticRequest_rs1}; // @[core.scala 250:34]
  wire [94:0] _arithmeticResult_arithmetic32_T_27 = _GEN_250 << singleCycleArithmeticRequest_rs2[4:0]; // @[core.scala 250:34]
  wire [31:0] _arithmeticResult_arithmetic32_T_30 = _arithmeticResult_arithmetic32_T_27[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _arithmeticResult_arithmetic32_T_32 = {_arithmeticResult_arithmetic32_T_30,
    _arithmeticResult_arithmetic32_T_27[31:0]}; // @[Cat.scala 33:92]
  wire [1:0] _arithmeticResult_arithmetic32_T_2 = {singleCycleArithmeticRequest_instruction[30],
    singleCycleArithmeticRequest_instruction[5]}; // @[Cat.scala 33:92]
  wire  _arithmeticResult_arithmetic32_T_3 = _arithmeticResult_arithmetic32_T_2 == 2'h3; // @[core.scala 248:58]
  wire [63:0] _arithmeticResult_arithmetic32_T_5 = singleCycleArithmeticRequest_rs1 - singleCycleArithmeticRequest_rs2; // @[core.scala 248:87]
  wire [31:0] _arithmeticResult_arithmetic32_T_8 = _arithmeticResult_arithmetic32_T_5[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _arithmeticResult_arithmetic32_T_10 = {_arithmeticResult_arithmetic32_T_8,
    _arithmeticResult_arithmetic32_T_5[31:0]}; // @[Cat.scala 33:92]
  wire [63:0] _arithmeticResult_arithmetic32_T_12 = singleCycleArithmeticRequest_rs1 + singleCycleArithmeticRequest_rs2; // @[core.scala 248:111]
  wire [31:0] _arithmeticResult_arithmetic32_T_15 = _arithmeticResult_arithmetic32_T_12[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _arithmeticResult_arithmetic32_T_17 = {_arithmeticResult_arithmetic32_T_15,
    _arithmeticResult_arithmetic32_T_12[31:0]}; // @[Cat.scala 33:92]
  wire [63:0] _arithmeticResult_arithmetic32_T_18 = _arithmeticResult_arithmetic32_T_2 == 2'h3 ?
    _arithmeticResult_arithmetic32_T_10 : _arithmeticResult_arithmetic32_T_17; // @[core.scala 248:20]
  wire [63:0] _GEN_36 = 2'h1 == _arithmeticResult_arithmetic32_T_56 ? _arithmeticResult_arithmetic32_T_32 :
    _arithmeticResult_arithmetic32_T_18; // @[core.scala 267:{8,8}]
  wire [63:0] _GEN_37 = 2'h2 == _arithmeticResult_arithmetic32_T_56 ? _arithmeticResult_arithmetic32_T_32 : _GEN_36; // @[core.scala 267:{8,8}]
  wire [63:0] _GEN_38 = 2'h3 == _arithmeticResult_arithmetic32_T_56 ? _arithmeticResult_arithmetic32_T_53 : _GEN_37; // @[core.scala 267:{8,8}]
  wire [63:0] _arithmeticResult_arithmetic64_T_26 = singleCycleArithmeticRequest_rs1 & singleCycleArithmeticRequest_rs2; // @[core.scala 265:22]
  wire [126:0] _arithmeticResult_arithmetic64_WIRE_7 = {{63'd0}, _arithmeticResult_arithmetic64_T_26}; // @[core.scala 257:{43,43}]
  wire [63:0] _arithmeticResult_arithmetic64_T_25 = singleCycleArithmeticRequest_rs1 | singleCycleArithmeticRequest_rs2; // @[core.scala 264:22]
  wire [126:0] _arithmeticResult_arithmetic64_WIRE_6 = {{63'd0}, _arithmeticResult_arithmetic64_T_25}; // @[core.scala 257:{43,43}]
  wire [63:0] _arithmeticResult_arithmetic64_T_21 = $signed(singleCycleArithmeticRequest_rs1) >>>
    singleCycleArithmeticRequest_rs2[5:0]; // @[core.scala 263:71]
  wire [63:0] _arithmeticResult_arithmetic64_T_23 = singleCycleArithmeticRequest_rs1 >> singleCycleArithmeticRequest_rs2
    [5:0]; // @[core.scala 263:84]
  wire [63:0] _arithmeticResult_arithmetic64_T_24 = singleCycleArithmeticRequest_instruction[30] ?
    _arithmeticResult_arithmetic64_T_21 : _arithmeticResult_arithmetic64_T_23; // @[core.scala 263:20]
  wire [126:0] _arithmeticResult_arithmetic64_WIRE_5 = {{63'd0}, _arithmeticResult_arithmetic64_T_24}; // @[core.scala 257:{43,43}]
  wire [63:0] _arithmeticResult_arithmetic64_T_15 = singleCycleArithmeticRequest_rs1 ^ singleCycleArithmeticRequest_rs2; // @[core.scala 262:22]
  wire [126:0] _arithmeticResult_arithmetic64_WIRE_4 = {{63'd0}, _arithmeticResult_arithmetic64_T_15}; // @[core.scala 257:{43,43}]
  wire  _arithmeticResult_arithmetic64_T_14 = singleCycleArithmeticRequest_rs1 < singleCycleArithmeticRequest_rs2; // @[core.scala 261:22]
  wire [126:0] _arithmeticResult_arithmetic64_WIRE_3 = {{126'd0}, _arithmeticResult_arithmetic64_T_14}; // @[core.scala 257:{43,43}]
  wire  _arithmeticResult_arithmetic64_T_13 = $signed(singleCycleArithmeticRequest_rs1) < $signed(
    singleCycleArithmeticRequest_rs2); // @[core.scala 260:29]
  wire [126:0] _arithmeticResult_arithmetic64_WIRE_2 = {{126'd0}, _arithmeticResult_arithmetic64_T_13}; // @[core.scala 257:{43,43}]
  wire [126:0] _GEN_252 = {{63'd0}, singleCycleArithmeticRequest_rs1}; // @[core.scala 259:22]
  wire [126:0] _arithmeticResult_arithmetic64_T_10 = _GEN_252 << singleCycleArithmeticRequest_rs2[5:0]; // @[core.scala 259:22]
  wire [63:0] _arithmeticResult_arithmetic64_T_8 = _arithmeticResult_arithmetic32_T_3 ?
    _arithmeticResult_arithmetic32_T_5 : _arithmeticResult_arithmetic32_T_12; // @[core.scala 258:20]
  wire [126:0] _arithmeticResult_arithmetic64_WIRE_0 = {{63'd0}, _arithmeticResult_arithmetic64_T_8}; // @[core.scala 257:{43,43}]
  wire [126:0] _GEN_40 = 3'h1 == singleCycleArithmeticRequest_instruction[14:12] ? _arithmeticResult_arithmetic64_T_10
     : _arithmeticResult_arithmetic64_WIRE_0; // @[core.scala 267:{8,8}]
  wire [126:0] _GEN_41 = 3'h2 == singleCycleArithmeticRequest_instruction[14:12] ? _arithmeticResult_arithmetic64_WIRE_2
     : _GEN_40; // @[core.scala 267:{8,8}]
  wire [126:0] _GEN_42 = 3'h3 == singleCycleArithmeticRequest_instruction[14:12] ? _arithmeticResult_arithmetic64_WIRE_3
     : _GEN_41; // @[core.scala 267:{8,8}]
  wire [126:0] _GEN_43 = 3'h4 == singleCycleArithmeticRequest_instruction[14:12] ? _arithmeticResult_arithmetic64_WIRE_4
     : _GEN_42; // @[core.scala 267:{8,8}]
  wire [126:0] _GEN_44 = 3'h5 == singleCycleArithmeticRequest_instruction[14:12] ? _arithmeticResult_arithmetic64_WIRE_5
     : _GEN_43; // @[core.scala 267:{8,8}]
  wire [126:0] _GEN_45 = 3'h6 == singleCycleArithmeticRequest_instruction[14:12] ? _arithmeticResult_arithmetic64_WIRE_6
     : _GEN_44; // @[core.scala 267:{8,8}]
  wire [126:0] _GEN_46 = 3'h7 == singleCycleArithmeticRequest_instruction[14:12] ? _arithmeticResult_arithmetic64_WIRE_7
     : _GEN_45; // @[core.scala 267:{8,8}]
  wire [126:0] arithmeticResult = singleCycleArithmeticRequest_instruction[3] ? {{63'd0}, _GEN_38} : _GEN_46; // @[core.scala 267:8]
  wire [63:0] fwdFrom_0_result = arithmeticResult[63:0]; // @[core.scala 228:33 269:21]
  wire [51:0] _arithmeticImm_T_2 = prf_toExec_instruction[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 77:12]
  wire [63:0] arithmeticImm = {_arithmeticImm_T_2,prf_toExec_instruction[31:20]}; // @[Cat.scala 33:92]
  wire [2:0] _singleCycleArithmeticRequest_valid_T_1 = prf_toExec_instruction[4:2] & 3'h5; // @[core.scala 274:91]
  wire  _singleCycleArithmeticRequest_rs2_T_5 = fwdFrom_0_valid & singleCycleArithmeticRequest_prfDest ==
    prf_toExec_rs2Addr; // @[core.scala 283:34]
  wire  _singleCycleArithmeticRequest_rs2_T_7 = fwdBuffers_0_valid & fwdBuffers_0_prfDest == prf_toExec_rs2Addr; // @[core.scala 283:34]
  wire  _singleCycleArithmeticRequest_rs2_T_9 = fwdBuffers_1_valid & fwdBuffers_1_prfDest == prf_toExec_rs2Addr; // @[core.scala 283:34]
  wire [63:0] _singleCycleArithmeticRequest_rs2_T_10 = _singleCycleArithmeticRequest_rs2_T_9 ? fwdBuffers_1_result :
    prf_toExec_rs2Data; // @[Mux.scala 101:16]
  wire [3:0] _T_30 = branchEvals_branchMask & singleCycleArithmeticRequest_branchMask; // @[core.scala 302:53]
  wire [4:0] _extnMRequest_valid_T_1 = prf_toExec_instruction[6:2] & 5'h1d; // @[core.scala 308:75]
  wire  _GEN_54 = _T_14 ? 1'h0 : prf_toExec_valid & 5'hc == _extnMRequest_valid_T_1 & prf_toExec_instruction[25]; // @[core.scala 308:22 315:83 316:26]
  wire  _GEN_56 = branchEvals_valid ? _GEN_54 : prf_toExec_valid & 5'hc == _extnMRequest_valid_T_1 &
    prf_toExec_instruction[25]; // @[core.scala 308:22 311:25]
  wire [32:0] _partialMuls32x32_T_7 = {extnMRequest_rs1[63],extnMRequest_rs1[63:32]}; // @[core.scala 331:57]
  wire [32:0] _partialMuls32x32_T_10 = {1'h0,extnMRequest_rs2[31:0]}; // @[core.scala 331:105]
  wire [32:0] _partialMuls32x32_T_15 = {1'h0,extnMRequest_rs1[31:0]}; // @[core.scala 333:44]
  wire [32:0] _partialMuls32x32_T_19 = {extnMRequest_rs2[63],extnMRequest_rs2[63:32]}; // @[core.scala 333:105]
  wire [32:0] _partialMuls32x32_T_28 = {1'h0,extnMRequest_rs2[63:32]}; // @[core.scala 335:106]
  wire [31:0] _partialMuls32x32_T_30 = extnMRequest_rs1[63:32]; // @[core.scala 336:30]
  wire [31:0] _partialMuls32x32_T_32 = extnMRequest_rs2[63:32]; // @[core.scala 336:64]
  wire [31:0] _partialMuls32x32_T_34 = extnMRequest_rs1[31:0]; // @[core.scala 337:29]
  wire [31:0] _partialMuls32x32_T_36 = extnMRequest_rs2[31:0]; // @[core.scala 337:62]
  reg [63:0] narrowMuls_0; // @[core.scala 339:23]
  reg [63:0] narrowMuls_1; // @[core.scala 339:23]
  reg [63:0] narrowMuls_2; // @[core.scala 339:23]
  reg [63:0] narrowMuls_3; // @[core.scala 339:23]
  reg [63:0] narrowMuls_4; // @[core.scala 339:23]
  reg [63:0] narrowMuls_5; // @[core.scala 339:23]
  reg [63:0] narrowMuls_6; // @[core.scala 339:23]
  reg [63:0] narrowMuls_7; // @[core.scala 339:23]
  reg [63:0] narrowMuls_8; // @[core.scala 339:23]
  wire [65:0] _T_39 = $signed(_partialMuls32x32_T_7) * $signed(_partialMuls32x32_T_10); // @[core.scala 340:41]
  wire [65:0] _T_40 = $signed(_partialMuls32x32_T_15) * $signed(_partialMuls32x32_T_19); // @[core.scala 340:41]
  wire [65:0] _T_41 = $signed(_partialMuls32x32_T_7) * $signed(_partialMuls32x32_T_28); // @[core.scala 340:41]
  wire [95:0] _muls_0_T = {narrowMuls_1,32'h0}; // @[Cat.scala 33:92]
  wire [95:0] _GEN_94 = {{32'd0}, narrowMuls_0}; // @[core.scala 343:29]
  wire [95:0] _muls_1_T = {narrowMuls_5,32'h0}; // @[Cat.scala 33:92]
  wire [95:0] _GEN_108 = {{32'd0}, narrowMuls_3}; // @[core.scala 344:28]
  wire [95:0] _muls_2_T = {narrowMuls_6,32'h0}; // @[Cat.scala 33:92]
  wire [31:0] _muls_3_T_2 = narrowMuls_4[63] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [95:0] _muls_3_T_3 = {_muls_3_T_2,narrowMuls_4}; // @[Cat.scala 33:92]
  wire [95:0] _muls_3_T_4 = {narrowMuls_7,32'h0}; // @[Cat.scala 33:92]
  wire [95:0] _muls_4_T = {narrowMuls_2,32'h0}; // @[Cat.scala 33:92]
  wire [31:0] _extnMResponse_result_T_4 = muls_5[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _extnMResponse_result_T_6 = {_extnMResponse_result_T_4,muls_5[31:0]}; // @[Cat.scala 33:92]
  wire [31:0] _extnMResponse_result_T_9 = muls_4[95] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [127:0] _extnMResponse_result_T_10 = {_extnMResponse_result_T_9,muls_4}; // @[Cat.scala 33:92]
  wire [127:0] _extnMResponse_result_T_11 = {muls_3,32'h0}; // @[Cat.scala 33:92]
  wire [127:0] _extnMResponse_result_T_13 = _extnMResponse_result_T_10 + _extnMResponse_result_T_11; // @[core.scala 355:42]
  wire [127:0] _extnMResponse_result_T_27 = {muls_2,32'h0}; // @[Cat.scala 33:92]
  wire [127:0] _extnMResponse_result_T_29 = _extnMResponse_result_T_10 + _extnMResponse_result_T_27; // @[core.scala 357:42]
  wire [127:0] _extnMResponse_result_T_31 = {muls_1,32'h0}; // @[Cat.scala 33:92]
  wire [127:0] _GEN_144 = {{32'd0}, muls_0}; // @[core.scala 358:14]
  wire [127:0] _extnMResponse_result_T_33 = _GEN_144 + _extnMResponse_result_T_31; // @[core.scala 358:14]
  wire [63:0] _GEN_58 = 2'h1 == extnMServicing_instruction[13:12] ? _extnMResponse_result_T_13[127:64] :
    _extnMResponse_result_T_13[63:0]; // @[core.scala 353:{30,30}]
  wire [63:0] _GEN_59 = 2'h2 == extnMServicing_instruction[13:12] ? _extnMResponse_result_T_29[127:64] : _GEN_58; // @[core.scala 353:{30,30}]
  wire [63:0] _GEN_60 = 2'h3 == extnMServicing_instruction[13:12] ? _extnMResponse_result_T_33[127:64] : _GEN_59; // @[core.scala 353:{30,30}]
  wire [63:0] _extnMResponse_result_T_36 = extnMServicing_instruction[3] ? _extnMResponse_result_T_6 : _GEN_60; // @[core.scala 353:30]
  wire [63:0] _GEN_61 = extnMServicing_valid & (~(|extnMServicing_instruction[24:20]) | ~(|extnMServicing_instruction[19
    :15])) ? 64'h0 : _extnMResponse_result_T_36; // @[core.scala 360:118 353:24 361:26]
  wire [3:0] _T_55 = extnMRequest_branchMask ^ branchEvals_branchMask; // @[core.scala 368:103]
  wire [3:0] _T_56 = extnMRequest_branchMask & branchEvals_branchMask; // @[core.scala 368:130]
  wire  _T_57 = |_T_56; // @[core.scala 368:154]
  wire [3:0] _T_58 = extnMPartialServicing_branchMask ^ branchEvals_branchMask; // @[core.scala 368:103]
  wire [3:0] _T_59 = extnMPartialServicing_branchMask & branchEvals_branchMask; // @[core.scala 368:130]
  wire  _T_60 = |_T_59; // @[core.scala 368:154]
  wire [3:0] _T_64 = extnMServicing_branchMask & branchEvals_branchMask; // @[core.scala 374:93]
  wire  _T_67 = |_T_64; // @[core.scala 374:123]
  wire  _GEN_67 = _T_67 & extnMServicing_valid ? 1'h0 : extnMServicing_valid; // @[core.scala 376:{101,107} 364:23]
  reg [3:0] divBranchMask; // @[core.scala 380:26]
  wire [4:0] _T_74 = {scheduler_release_instruction[25],scheduler_release_instruction[14],scheduler_release_instruction[
    6:4]}; // @[Cat.scala 33:92]
  wire  _T_75 = _T_74 == 5'h1b; // @[core.scala 382:115]
  wire  _T_76 = scheduler_release_fired & _T_75; // @[core.scala 381:32]
  wire [3:0] _mExtensionReady_T = branchEvals_branchMask & scheduler_release_branchMask; // @[core.scala 384:77]
  wire  _mExtensionReady_T_2 = branchEvals_valid & |_mExtensionReady_T; // @[core.scala 384:52]
  wire [3:0] _divBranchMask_T_3 = scheduler_release_branchMask ^ branchEvals_branchMask; // @[core.scala 386:133]
  wire [3:0] _divBranchMask_T_4 = _mExtensionReady_T_2 ? _divBranchMask_T_3 : scheduler_release_branchMask; // @[core.scala 386:25]
  wire  _GEN_77 = _T_76 ? branchEvals_valid & |_mExtensionReady_T & _T : mExtensionReady; // @[core.scala 382:132 384:21 117:32]
  wire [3:0] _GEN_78 = _T_76 ? _divBranchMask_T_4 : divBranchMask; // @[core.scala 382:132 386:19 380:26]
  wire [3:0] _T_78 = branchEvals_branchMask & divBranchMask; // @[core.scala 389:51]
  wire [3:0] _divBranchMask_T_5 = divBranchMask ^ branchEvals_branchMask; // @[core.scala 391:40]
  wire  _GEN_80 = _T | _GEN_77; // @[core.scala 393:31 394:25]
  wire  _GEN_82 = branchEvals_valid & |_T_78 ? _GEN_80 : _GEN_77; // @[core.scala 389:73]
  wire  _GEN_84 = ~mExtensionReady ? _GEN_82 : _GEN_77; // @[core.scala 388:26]
  wire  _GEN_85 = extnMResponse_valid & extnResponseInstruction[14] | _GEN_84; // @[core.scala 398:{67,85}]
  wire [64:0] _division_remainder_T_2 = {division_remainder[63:0],division_quotient[64]}; // @[Cat.scala 33:92]
  wire [64:0] _division_remainder_T_6 = 65'h0 - division_divisor; // @[core.scala 400:134]
  wire [64:0] _division_remainder_T_7 = division_remainder[64] ? division_divisor : _division_remainder_T_6; // @[core.scala 400:84]
  wire [64:0] _division_remainder_T_9 = _division_remainder_T_2 + _division_remainder_T_7; // @[core.scala 400:79]
  wire  _division_quotient_T_12 = ~_division_remainder_T_9[64]; // @[core.scala 401:54]
  wire [64:0] _division_quotient_T_13 = {division_quotient[63:0],_division_quotient_T_12}; // @[Cat.scala 33:92]
  wire [6:0] _division_counter_T_1 = division_counter - 7'h1; // @[core.scala 402:40]
  wire [64:0] _division_divisor_T_1 = {33'h0,extnMRequest_rs2[31:0]}; // @[Cat.scala 33:92]
  wire [64:0] _division_quotient_T_15 = {33'h0,extnMRequest_rs1[31:0]}; // @[Cat.scala 33:92]
  wire [64:0] _GEN_86 = extnMRequest_instruction[3] ? _division_divisor_T_1 : {{1'd0}, extnMRequest_rs2}; // @[core.scala 406:22 408:46 409:24]
  wire [64:0] _GEN_87 = extnMRequest_instruction[3] ? _division_quotient_T_15 : {{1'd0}, extnMRequest_rs1}; // @[core.scala 407:23 408:46 410:25]
  wire [63:0] _division_quotient_T_17 = 64'h0 - extnMRequest_rs1; // @[core.scala 417:79]
  wire [64:0] _division_quotient_T_19 = {1'h0,_division_quotient_T_17}; // @[Cat.scala 33:92]
  wire [64:0] _GEN_88 = extnMRequest_rs1[63] ? _division_quotient_T_19 : _GEN_87; // @[core.scala 417:{41,61}]
  wire [63:0] _division_divisor_T_3 = 64'h0 - extnMRequest_rs2; // @[core.scala 418:78]
  wire [64:0] _division_divisor_T_5 = {1'h0,_division_divisor_T_3}; // @[Cat.scala 33:92]
  wire [64:0] _GEN_89 = extnMRequest_rs2[63] ? _division_divisor_T_5 : _GEN_86; // @[core.scala 418:{41,60}]
  wire [31:0] _division_quotient_T_22 = 32'h0 - extnMRequest_rs1[31:0]; // @[core.scala 420:82]
  wire [64:0] _division_quotient_T_24 = {33'h0,_division_quotient_T_22}; // @[Cat.scala 33:92]
  wire [31:0] _division_divisor_T_8 = 32'h0 - extnMRequest_rs2[31:0]; // @[core.scala 421:81]
  wire [64:0] _division_divisor_T_10 = {33'h0,_division_divisor_T_8}; // @[Cat.scala 33:92]
  wire  _GEN_101 = extnMRequest_valid & extnMRequest_instruction[14] ? extnMRequest_valid : division_request_valid; // @[core.scala 404:67 413:22 213:25]
  wire [3:0] _GEN_107 = extnMRequest_valid & extnMRequest_instruction[14] ? extnMRequest_branchMask :
    division_request_branchMask; // @[core.scala 404:67 413:22 213:25]
  wire  _extnMResponse_result_quotient32_T_6 = ~(division_quotient == 65'h1ffffffffffffffff); // @[core.scala 429:99]
  wire [64:0] _extnMResponse_result_quotient32_T_9 = 65'h0 - division_quotient; // @[core.scala 429:125]
  wire [31:0] extnMResponse_result_quotient32 = (division_request_rs1[31] ^ division_request_rs2[31]) & ~(
    division_quotient == 65'h1ffffffffffffffff) ? _extnMResponse_result_quotient32_T_9[31:0] : division_quotient[31:0]; // @[core.scala 429:27]
  wire [64:0] _extnMResponse_result_remainder64Unsigned_T_3 = division_remainder + division_divisor; // @[core.scala 430:87]
  wire [64:0] extnMResponse_result_remainder64Unsigned = division_remainder[64] ?
    _extnMResponse_result_remainder64Unsigned_T_3 : division_remainder; // @[core.scala 430:36]
  wire [64:0] _extnMResponse_result_remainder32Signed_T_3 = 65'h0 - extnMResponse_result_remainder64Unsigned; // @[core.scala 431:70]
  wire [64:0] extnMResponse_result_remainder32Signed = division_request_rs1[31] ?
    _extnMResponse_result_remainder32Signed_T_3 : extnMResponse_result_remainder64Unsigned; // @[core.scala 431:34]
  wire [64:0] _extnMResponse_result_T_47 = (division_request_rs1[63] ^ division_request_rs2[63]) &
    _extnMResponse_result_quotient32_T_6 ? _extnMResponse_result_quotient32_T_9 : division_quotient; // @[core.scala 434:10]
  wire [64:0] _extnMResponse_result_T_52 = division_request_rs1[63] ? _extnMResponse_result_remainder32Signed_T_3 :
    extnMResponse_result_remainder64Unsigned; // @[core.scala 436:10]
  wire [31:0] _extnMResponse_result_T_55 = extnMResponse_result_quotient32[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _extnMResponse_result_T_57 = {_extnMResponse_result_T_55,extnMResponse_result_quotient32}; // @[Cat.scala 33:92]
  wire [31:0] _extnMResponse_result_T_60 = division_quotient[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _extnMResponse_result_T_62 = {_extnMResponse_result_T_60,division_quotient[31:0]}; // @[Cat.scala 33:92]
  wire [31:0] _extnMResponse_result_T_65 = extnMResponse_result_remainder32Signed[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _extnMResponse_result_T_67 = {_extnMResponse_result_T_65,extnMResponse_result_remainder32Signed[31:0]}; // @[Cat.scala 33:92]
  wire [31:0] _extnMResponse_result_T_70 = extnMResponse_result_remainder64Unsigned[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _extnMResponse_result_T_72 = {_extnMResponse_result_T_70,extnMResponse_result_remainder64Unsigned[31:0]}; // @[Cat.scala 33:92]
  wire [2:0] _extnMResponse_result_T_75 = {division_request_instruction[3],division_request_instruction[13:12]}; // @[Cat.scala 33:92]
  wire [64:0] _GEN_110 = 3'h1 == _extnMResponse_result_T_75 ? division_quotient : _extnMResponse_result_T_47; // @[core.scala 428:{26,26}]
  wire [64:0] _GEN_111 = 3'h2 == _extnMResponse_result_T_75 ? _extnMResponse_result_T_52 : _GEN_110; // @[core.scala 428:{26,26}]
  wire [64:0] _GEN_112 = 3'h3 == _extnMResponse_result_T_75 ? extnMResponse_result_remainder64Unsigned : _GEN_111; // @[core.scala 428:{26,26}]
  wire [64:0] _extnMResponse_result_WIRE_1_4 = {{1'd0}, _extnMResponse_result_T_57}; // @[core.scala 433:{14,14}]
  wire [64:0] _GEN_113 = 3'h4 == _extnMResponse_result_T_75 ? _extnMResponse_result_WIRE_1_4 : _GEN_112; // @[core.scala 428:{26,26}]
  wire [64:0] _extnMResponse_result_WIRE_1_5 = {{1'd0}, _extnMResponse_result_T_62}; // @[core.scala 433:{14,14}]
  wire [64:0] _GEN_114 = 3'h5 == _extnMResponse_result_T_75 ? _extnMResponse_result_WIRE_1_5 : _GEN_113; // @[core.scala 428:{26,26}]
  wire [64:0] _extnMResponse_result_WIRE_1_6 = {{1'd0}, _extnMResponse_result_T_67}; // @[core.scala 433:{14,14}]
  wire [64:0] _GEN_115 = 3'h6 == _extnMResponse_result_T_75 ? _extnMResponse_result_WIRE_1_6 : _GEN_114; // @[core.scala 428:{26,26}]
  wire [64:0] _extnMResponse_result_WIRE_1_7 = {{1'd0}, _extnMResponse_result_T_72}; // @[core.scala 433:{14,14}]
  wire [64:0] _GEN_116 = 3'h7 == _extnMResponse_result_T_75 ? _extnMResponse_result_WIRE_1_7 : _GEN_115; // @[core.scala 428:{26,26}]
  wire [3:0] _T_106 = division_request_branchMask & branchEvals_branchMask; // @[core.scala 451:41]
  wire  _T_107 = |_T_106; // @[core.scala 451:65]
  wire [64:0] _GEN_120 = division_request_valid & ~(|division_counter) ? _GEN_116 : {{1'd0}, _GEN_61}; // @[core.scala 426:57 428:26]
  wire  _GEN_124 = division_request_valid & ~(|division_counter) ? 1'h0 : _GEN_101; // @[core.scala 426:57 449:28]
  wire  _GEN_126 = _T & _T_57 ? 1'h0 : _GEN_124; // @[core.scala 458:{112,87}]
  wire [3:0] _division_request_branchMask_T_1 = division_request_branchMask ^ branchEvals_branchMask; // @[core.scala 460:130]
  reg  branchPCs_0_valid; // @[core.scala 475:26]
  reg [63:0] branchPCs_0_pc; // @[core.scala 475:26]
  reg [3:0] branchPCs_0_branchMask; // @[core.scala 475:26]
  reg  branchPCs_1_valid; // @[core.scala 475:26]
  reg [63:0] branchPCs_1_pc; // @[core.scala 475:26]
  reg [3:0] branchPCs_1_branchMask; // @[core.scala 475:26]
  reg  branchPCs_2_valid; // @[core.scala 475:26]
  reg [63:0] branchPCs_2_pc; // @[core.scala 475:26]
  reg [3:0] branchPCs_2_branchMask; // @[core.scala 475:26]
  reg  branchPCs_3_valid; // @[core.scala 475:26]
  reg [63:0] branchPCs_3_pc; // @[core.scala 475:26]
  reg [3:0] branchPCs_3_branchMask; // @[core.scala 475:26]
  reg  predictedPCs_0_valid; // @[core.scala 482:29]
  reg [63:0] predictedPCs_0_pc; // @[core.scala 482:29]
  reg  predictedPCs_1_valid; // @[core.scala 482:29]
  reg [63:0] predictedPCs_1_pc; // @[core.scala 482:29]
  reg  predictedPCs_2_valid; // @[core.scala 482:29]
  reg [63:0] predictedPCs_2_pc; // @[core.scala 482:29]
  reg  predictedPCs_3_valid; // @[core.scala 482:29]
  reg [63:0] predictedPCs_3_pc; // @[core.scala 482:29]
  reg  branchInstruction_valid; // @[core.scala 487:34]
  reg [63:0] branchInstruction_rs1; // @[core.scala 487:34]
  reg [63:0] branchInstruction_rs2; // @[core.scala 487:34]
  reg [3:0] branchInstruction_robAddr; // @[core.scala 487:34]
  reg [31:0] branchInstruction_instruction; // @[core.scala 487:34]
  reg [63:0] branchInstruction_immediate; // @[core.scala 487:34]
  wire [63:0] _branchInstruction_immediate_T_6 = {_arithmeticImm_T_2,prf_toExec_instruction[7],prf_toExec_instruction[30
    :25],prf_toExec_instruction[11:8],1'h0}; // @[Cat.scala 33:92]
  wire [43:0] _branchInstruction_immediate_T_14 = prf_toExec_instruction[31] ? 44'hfffffffffff : 44'h0; // @[Bitwise.scala 77:12]
  wire [63:0] _branchInstruction_immediate_T_18 = {_branchInstruction_immediate_T_14,prf_toExec_instruction[19:12],
    prf_toExec_instruction[20],prf_toExec_instruction[30:21],1'h0}; // @[Cat.scala 33:92]
  reg [3:0] branchEvals_robAddr; // @[core.scala 509:28]
  reg [63:0] branchEvals_nextPC; // @[core.scala 509:28]
  wire [5:0] _GEN_140 = prf_toExec_valid & prf_toExec_instruction[6:5] == 2'h3 ? prf_toExec_robAddr : {{2'd0},
    branchInstruction_robAddr}; // @[core.scala 521:71 529:31 487:34]
  wire [3:0] _T_128 = branchEvals_branchMask & prf_toExec_branchmask; // @[core.scala 537:53]
  wire [63:0] branchTaken_rs1 = |branchInstruction_instruction[19:15] ? branchInstruction_rs1 : 64'h0; // @[core.scala 554:18]
  wire [63:0] branchTaken_rs2 = |branchInstruction_instruction[24:20] ? branchInstruction_rs2 : 64'h0; // @[core.scala 555:18]
  wire  branchTaken_conditionEval_0 = branchTaken_rs1 == branchTaken_rs2; // @[core.scala 559:41]
  wire [63:0] _branchTaken_conditionEval_T_2 = |branchInstruction_instruction[19:15] ? branchInstruction_rs1 : 64'h0; // @[core.scala 559:67]
  wire [63:0] _branchTaken_conditionEval_T_3 = |branchInstruction_instruction[24:20] ? branchInstruction_rs2 : 64'h0; // @[core.scala 559:80]
  wire  branchTaken_conditionEval_4 = $signed(_branchTaken_conditionEval_T_2) < $signed(_branchTaken_conditionEval_T_3); // @[core.scala 559:74]
  wire  branchTaken_conditionEval_6 = branchTaken_rs1 < branchTaken_rs2; // @[core.scala 559:92]
  wire  branchTaken_conditionEval_1 = ~branchTaken_conditionEval_0; // @[core.scala 559:125]
  wire  branchTaken_conditionEval_5 = ~branchTaken_conditionEval_4; // @[core.scala 559:125]
  wire  branchTaken_conditionEval_7 = ~branchTaken_conditionEval_6; // @[core.scala 559:125]
  wire  nextCorrectPC_conditionEval_0 = branchInstruction_rs1 == branchInstruction_rs2; // @[core.scala 579:11]
  wire  nextCorrectPC_conditionEval_1 = branchInstruction_rs1 != branchInstruction_rs2; // @[core.scala 580:11]
  wire  nextCorrectPC_conditionEval_4 = $signed(branchInstruction_rs1) < $signed(branchInstruction_rs2); // @[core.scala 583:18]
  wire  nextCorrectPC_conditionEval_5 = $signed(branchInstruction_rs1) >= $signed(branchInstruction_rs2); // @[core.scala 584:18]
  wire  nextCorrectPC_conditionEval_6 = branchInstruction_rs1 < branchInstruction_rs2; // @[core.scala 585:11]
  wire  nextCorrectPC_conditionEval_7 = branchInstruction_rs1 >= branchInstruction_rs2; // @[core.scala 586:11]
  wire [63:0] _nextCorrectPC_T_2 = branchPCs_0_pc + branchInstruction_immediate; // @[core.scala 590:50]
  wire [63:0] _nextCorrectPC_T_4 = branchPCs_0_pc + 64'h4; // @[core.scala 590:66]
  wire  _GEN_149 = 3'h1 == branchInstruction_instruction[14:12] ? nextCorrectPC_conditionEval_1 :
    nextCorrectPC_conditionEval_0; // @[core.scala 590:{10,10}]
  wire  _GEN_150 = 3'h2 == branchInstruction_instruction[14:12] ? 1'h0 : _GEN_149; // @[core.scala 590:{10,10}]
  wire  _GEN_151 = 3'h3 == branchInstruction_instruction[14:12] ? 1'h0 : _GEN_150; // @[core.scala 590:{10,10}]
  wire  _GEN_152 = 3'h4 == branchInstruction_instruction[14:12] ? nextCorrectPC_conditionEval_4 : _GEN_151; // @[core.scala 590:{10,10}]
  wire  _GEN_153 = 3'h5 == branchInstruction_instruction[14:12] ? nextCorrectPC_conditionEval_5 : _GEN_152; // @[core.scala 590:{10,10}]
  wire  _GEN_154 = 3'h6 == branchInstruction_instruction[14:12] ? nextCorrectPC_conditionEval_6 : _GEN_153; // @[core.scala 590:{10,10}]
  wire  _GEN_155 = 3'h7 == branchInstruction_instruction[14:12] ? nextCorrectPC_conditionEval_7 : _GEN_154; // @[core.scala 590:{10,10}]
  wire [63:0] _nextCorrectPC_T_5 = _GEN_155 ? _nextCorrectPC_T_2 : _nextCorrectPC_T_4; // @[core.scala 590:10]
  wire [63:0] _nextCorrectPC_T_7 = branchInstruction_rs1 + branchInstruction_immediate; // @[core.scala 591:11]
  wire [63:0] _GEN_157 = 2'h1 == branchInstruction_instruction[3:2] ? _nextCorrectPC_T_7 : _nextCorrectPC_T_5; // @[core.scala 596:{22,22}]
  wire [63:0] _GEN_158 = 2'h2 == branchInstruction_instruction[3:2] ? 64'h0 : _GEN_157; // @[core.scala 596:{22,22}]
  wire [63:0] _GEN_159 = 2'h3 == branchInstruction_instruction[3:2] ? _nextCorrectPC_T_2 : _GEN_158; // @[core.scala 596:{22,22}]
  wire  _T_133 = branchPCs_0_valid & branchPCs_1_valid; // @[core.scala 604:46]
  wire  _T_134 = branchPCs_0_valid & branchPCs_1_valid & branchPCs_2_valid; // @[core.scala 604:46]
  wire [63:0] _GEN_161 = ~branchPCs_0_valid ? decode_branchPCs_branchPC : branchPCs_0_pc; // @[core.scala 605:82 607:12 475:26]
  wire [3:0] _GEN_162 = ~branchPCs_0_valid ? decode_branchPCs_branchMask : branchPCs_0_branchMask; // @[core.scala 605:82 608:20 475:26]
  wire  _T_138 = ~branchPCs_1_valid; // @[core.scala 605:70]
  wire [63:0] _GEN_164 = branchPCs_0_valid & ~branchPCs_1_valid ? decode_branchPCs_branchPC : branchPCs_1_pc; // @[core.scala 605:82 607:12 475:26]
  wire [3:0] _GEN_165 = branchPCs_0_valid & ~branchPCs_1_valid ? decode_branchPCs_branchMask : branchPCs_1_branchMask; // @[core.scala 605:82 608:20 475:26]
  wire  _T_140 = ~branchPCs_2_valid; // @[core.scala 605:70]
  wire [63:0] _GEN_167 = _T_133 & ~branchPCs_2_valid ? decode_branchPCs_branchPC : branchPCs_2_pc; // @[core.scala 605:82 607:12 475:26]
  wire [3:0] _GEN_168 = _T_133 & ~branchPCs_2_valid ? decode_branchPCs_branchMask : branchPCs_2_branchMask; // @[core.scala 605:82 608:20 475:26]
  wire  _T_142 = ~branchPCs_3_valid; // @[core.scala 605:70]
  wire  _T_145 = branchEvals_valid & _T; // @[core.scala 610:24]
  wire  entry_1_valid = branchPCs_1_valid | decode_branchPCs_branchPCReady & (_T_138 & branchPCs_0_valid); // @[core.scala 616:32]
  wire  entry_2_valid = branchPCs_2_valid | decode_branchPCs_branchPCReady & (_T_140 & _T_133); // @[core.scala 616:32]
  wire  entry_3_valid = branchPCs_3_valid | decode_branchPCs_branchPCReady & (_T_142 & _T_134); // @[core.scala 616:32]
  wire  _T_151 = predictedPCs_0_valid & predictedPCs_1_valid; // @[core.scala 628:49]
  wire  _T_152 = predictedPCs_0_valid & predictedPCs_1_valid & predictedPCs_2_valid; // @[core.scala 628:49]
  wire [63:0] _GEN_193 = ~predictedPCs_0_valid ? decode_branchPCs_predictedPC : predictedPCs_0_pc; // @[core.scala 629:82 631:12 482:29]
  wire  _T_156 = ~predictedPCs_1_valid; // @[core.scala 629:70]
  wire [63:0] _GEN_195 = predictedPCs_0_valid & ~predictedPCs_1_valid ? decode_branchPCs_predictedPC : predictedPCs_1_pc
    ; // @[core.scala 629:82 631:12 482:29]
  wire  _T_158 = ~predictedPCs_2_valid; // @[core.scala 629:70]
  wire [63:0] _GEN_197 = _T_151 & ~predictedPCs_2_valid ? decode_branchPCs_predictedPC : predictedPCs_2_pc; // @[core.scala 629:82 631:12 482:29]
  wire  _T_160 = ~predictedPCs_3_valid; // @[core.scala 629:70]
  wire  entry_5_valid = predictedPCs_1_valid | decode_branchPCs_predictedPCReady & (_T_156 & predictedPCs_0_valid); // @[core.scala 639:32]
  wire  entry_6_valid = predictedPCs_2_valid | decode_branchPCs_predictedPCReady & (_T_158 & _T_151); // @[core.scala 639:32]
  wire  entry_7_valid = predictedPCs_3_valid | decode_branchPCs_predictedPCReady & (_T_160 & _T_152); // @[core.scala 639:32]
  reg  fetch_branchRes_branchTaken_REG; // @[core.scala 676:41]
  wire  _GEN_215 = 3'h1 == branchInstruction_instruction[14:12] ? branchTaken_conditionEval_1 :
    branchTaken_conditionEval_0; // @[core.scala 676:{41,41}]
  wire  _GEN_216 = 3'h2 == branchInstruction_instruction[14:12] ? branchTaken_conditionEval_0 : _GEN_215; // @[core.scala 676:{41,41}]
  wire  _GEN_217 = 3'h3 == branchInstruction_instruction[14:12] ? branchTaken_conditionEval_1 : _GEN_216; // @[core.scala 676:{41,41}]
  reg [63:0] fetch_branchRes_pc_REG; // @[core.scala 678:32]
  reg [63:0] rob_execPorts_0_mtval_REG; // @[core.scala 712:36]
  reg  REG; // @[core.scala 733:129]
  reg [5:0] prf_fromStore_rs2Addr_REG; // @[core.scala 769:43]
  reg [5:0] prf_fromStore_rs2Addr_REG_1; // @[core.scala 769:35]
  reg  prf_fromStore_valid_REG; // @[core.scala 770:41]
  reg  prf_fromStore_valid_REG_1; // @[core.scala 770:33]
  wire  _memAccess_initiateFence_T = rob_commit_fired & rob_commit_is_fence; // @[core.scala 812:47]
  reg [1:0] fenceState_state; // @[core.scala 816:27]
  reg [3:0] fenceState_branchMask; // @[core.scala 816:27]
  wire [19:0] _T_188 = fetch_toDecode_instruction[19:0] & 20'hfefff; // @[core.scala 825:72]
  wire [19:0] _T_195 = decode_toExec_instruction[19:0] & 20'hfefff; // @[core.scala 834:76]
  wire [1:0] _GEN_223 = decode_toExec_fired & _T_195 == 20'hf ? 2'h2 : fenceState_state; // @[core.scala 834:119 835:26 816:27]
  wire  _GEN_225 = _T_145 | rob_commit_fired & rob_commit_is_fence; // @[core.scala 812:27 830:54 832:33]
  wire [3:0] _T_199 = branchEvals_branchMask & fenceState_branchMask; // @[core.scala 840:57]
  wire  _T_201 = branchEvals_valid & |_T_199; // @[core.scala 840:30]
  wire [3:0] _fenceState_branchMask_T = fenceState_branchMask ^ branchEvals_branchMask; // @[core.scala 848:57]
  wire [3:0] _GEN_228 = _T_201 & branchEvals_passed ? _fenceState_branchMask_T : fenceState_branchMask; // @[core.scala 847:115 816:27 848:31]
  wire  _GEN_229 = rob_commit_fired & rob_commit_is_fence | rob_commit_fired & rob_commit_is_fence; // @[core.scala 812:27 844:59 845:33]
  wire [1:0] _GEN_230 = _memAccess_initiateFence_T ? 2'h0 : fenceState_state; // @[core.scala 844:59 846:26 816:27]
  wire [3:0] _GEN_231 = _memAccess_initiateFence_T ? fenceState_branchMask : _GEN_228; // @[core.scala 816:27 844:59]
  wire  _GEN_232 = branchEvals_valid & |_T_199 & _T | _GEN_229; // @[core.scala 840:110 842:33]
  wire [1:0] _GEN_233 = branchEvals_valid & |_T_199 & _T ? 2'h0 : _GEN_230; // @[core.scala 840:110 843:26]
  wire  _GEN_235 = 2'h2 == fenceState_state ? _GEN_232 : rob_commit_fired & rob_commit_is_fence; // @[core.scala 812:27 823:28]
  wire  _GEN_238 = 2'h1 == fenceState_state ? _GEN_225 : _GEN_235; // @[core.scala 823:28]
  wire  _GEN_242 = 2'h0 == fenceState_state ? rob_commit_fired & rob_commit_is_fence : _GEN_238; // @[core.scala 812:27 823:28]
  wire  _GEN_244 = _T_145 & fetch_cachelinesUpdatesResp_ready | _GEN_242; // @[core.scala 871:85 872:29]
  reg  REG_1; // @[core.scala 874:15]
  reg [2:0] branchCounter; // @[core.scala 987:30]
  wire  _branchCounter_T_2 = decode_fromFetch_fired & decode_fromFetch_instruction[6:4] == 3'h6; // @[core.scala 991:29]
  wire [2:0] _GEN_247 = {{2'd0}, _branchCounter_T_2}; // @[core.scala 988:34]
  wire [3:0] _branchCounter_T_3 = branchCounter + _GEN_247; // @[core.scala 988:34]
  wire [3:0] _GEN_248 = {{3'd0}, branchEvals_valid}; // @[core.scala 991:81]
  wire [4:0] _branchCounter_T_4 = _branchCounter_T_3 - _GEN_248; // @[core.scala 991:81]
  wire [4:0] _GEN_267 = _T_145 ? 5'h0 : _branchCounter_T_4; // @[core.scala 988:17 994:50 997:19]
  reg [3:0] lastBranchExecRob; // @[core.scala 1001:30]
  reg [63:0] lastBranchExecPC; // @[core.scala 1002:29]
  reg [63:0] lastBranchExecPC_REG; // @[core.scala 1005:32]
  reg  lastRetiredSystem; // @[core.scala 1021:34]
  reg [1:0] interruptInjectStatus; // @[core.scala 1024:38]
  wire  _T_231 = |branchCounter; // @[core.scala 1035:60]
  wire [1:0] _GEN_272 = branchInstruction_valid & branchInstruction_instruction[6:0] == 7'h63 ? 2'h2 :
    interruptInjectStatus; // @[core.scala 1036:135 1024:38 1037:79]
  wire  _GEN_273 = branchInstruction_valid & branchInstruction_instruction[6:0] == 7'h63 ? 1'h0 : predictedPCs_0_valid
     & _GEN_159 == predictedPCs_0_pc; // @[core.scala 1036:135 1040:76 598:22]
  wire [1:0] _GEN_274 = decode_fromFetch_fired ? 2'h0 : interruptInjectStatus; // @[core.scala 1050:110 1024:38 1050:86]
  wire [63:0] _GEN_275 = fetch_toDecode_instruction[6:0] != 7'hf & fetch_toDecode_instruction[6:0] != 7'h73 ? 64'h80000073
     : {{32'd0}, fetch_toDecode_instruction}; // @[core.scala 1043:162 1045:86 49:32]
  wire [1:0] _GEN_276 = fetch_toDecode_instruction[6:0] != 7'hf & fetch_toDecode_instruction[6:0] != 7'h73 ? _GEN_274 :
    interruptInjectStatus; // @[core.scala 1043:162 1024:38]
  wire [1:0] _GEN_277 = |branchCounter ? _GEN_272 : _GEN_276; // @[core.scala 1035:65]
  wire  _GEN_278 = |branchCounter ? _GEN_273 : predictedPCs_0_valid & _GEN_159 == predictedPCs_0_pc; // @[core.scala 1035:65 598:22]
  wire [63:0] _GEN_279 = |branchCounter ? {{32'd0}, fetch_toDecode_instruction} : _GEN_275; // @[core.scala 1035:65 49:32]
  wire [1:0] _GEN_280 = ~branchEvals_valid ? _GEN_277 : interruptInjectStatus; // @[core.scala 1024:38 1034:58]
  wire [63:0] _GEN_282 = ~branchEvals_valid ? _GEN_279 : {{32'd0}, fetch_toDecode_instruction}; // @[core.scala 1034:58 49:32]
  wire [63:0] _GEN_285 = decode_canTakeInterrupt ? _GEN_282 : {{32'd0}, fetch_toDecode_instruction}; // @[core.scala 1033:56 49:32]
  wire [1:0] _GEN_286 = decode_writeBackResult_fired ? 2'h0 : interruptInjectStatus; // @[core.scala 1024:38 1064:{44,68}]
  wire [63:0] _GEN_287 = rob_commit_robAddr == lastBranchExecRob ? 64'h80000073 : {{32'd0}, rob_commit_instruction}; // @[core.scala 1060:54 1062:44 683:38]
  wire [1:0] _GEN_288 = rob_commit_robAddr == lastBranchExecRob ? _GEN_286 : interruptInjectStatus; // @[core.scala 1024:38 1060:54]
  wire [63:0] _GEN_289 = 2'h3 == interruptInjectStatus ? _GEN_287 : {{32'd0}, rob_commit_instruction}; // @[core.scala 1025:33 683:38]
  wire [1:0] _GEN_290 = 2'h3 == interruptInjectStatus ? _GEN_288 : interruptInjectStatus; // @[core.scala 1025:33 1024:38]
  wire [63:0] _GEN_292 = 2'h2 == interruptInjectStatus ? {{32'd0}, rob_commit_instruction} : _GEN_289; // @[core.scala 1025:33 683:38]
  wire [63:0] _GEN_295 = 2'h1 == interruptInjectStatus ? _GEN_285 : {{32'd0}, fetch_toDecode_instruction}; // @[core.scala 1025:33 49:32]
  wire [63:0] _GEN_296 = 2'h1 == interruptInjectStatus ? {{32'd0}, rob_commit_instruction} : _GEN_292; // @[core.scala 1025:33 683:38]
  wire [63:0] _GEN_299 = 2'h0 == interruptInjectStatus ? {{32'd0}, fetch_toDecode_instruction} : _GEN_295; // @[core.scala 1025:33 49:32]
  wire [63:0] _GEN_300 = 2'h0 == interruptInjectStatus ? {{32'd0}, rob_commit_instruction} : _GEN_296; // @[core.scala 1025:33 683:38]
  wire [4:0] _GEN_249 = reset ? 5'h0 : _GEN_267; // @[core.scala 987:{30,30}]
  iCache icache ( // @[core.scala 19:22]
    .clock(icache_clock),
    .reset(icache_reset),
    .fromFetch_req_ready(icache_fromFetch_req_ready),
    .fromFetch_req_valid(icache_fromFetch_req_valid),
    .fromFetch_req_bits(icache_fromFetch_req_bits),
    .fromFetch_resp_ready(icache_fromFetch_resp_ready),
    .fromFetch_resp_valid(icache_fromFetch_resp_valid),
    .fromFetch_resp_bits(icache_fromFetch_resp_bits),
    .updateAllCachelines_ready(icache_updateAllCachelines_ready),
    .updateAllCachelines_fired(icache_updateAllCachelines_fired),
    .cachelinesUpdatesResp_ready(icache_cachelinesUpdatesResp_ready),
    .cachelinesUpdatesResp_fired(icache_cachelinesUpdatesResp_fired),
    .lowLevelMem_ARADDR(icache_lowLevelMem_ARADDR),
    .lowLevelMem_ARVALID(icache_lowLevelMem_ARVALID),
    .lowLevelMem_ARREADY(icache_lowLevelMem_ARREADY),
    .lowLevelMem_RDATA(icache_lowLevelMem_RDATA),
    .lowLevelMem_RLAST(icache_lowLevelMem_RLAST),
    .lowLevelMem_RVALID(icache_lowLevelMem_RVALID),
    .lowLevelMem_RREADY(icache_lowLevelMem_RREADY)
  );
  fetch fetch ( // @[core.scala 28:21]
    .clock(fetch_clock),
    .reset(fetch_reset),
    .cache_req_ready(fetch_cache_req_ready),
    .cache_req_valid(fetch_cache_req_valid),
    .cache_req_bits(fetch_cache_req_bits),
    .cache_resp_ready(fetch_cache_resp_ready),
    .cache_resp_valid(fetch_cache_resp_valid),
    .cache_resp_bits(fetch_cache_resp_bits),
    .toDecode_ready(fetch_toDecode_ready),
    .toDecode_fired(fetch_toDecode_fired),
    .toDecode_pc(fetch_toDecode_pc),
    .toDecode_instruction(fetch_toDecode_instruction),
    .toDecode_expected_valid(fetch_toDecode_expected_valid),
    .toDecode_expected_pc(fetch_toDecode_expected_pc),
    .branchRes_fired(fetch_branchRes_fired),
    .branchRes_branchTaken(fetch_branchRes_branchTaken),
    .branchRes_pc(fetch_branchRes_pc),
    .branchRes_pcAfterBrnach(fetch_branchRes_pcAfterBrnach),
    .carryOutFence_ready(fetch_carryOutFence_ready),
    .carryOutFence_fired(fetch_carryOutFence_fired),
    .updateAllCachelines_ready(fetch_updateAllCachelines_ready),
    .updateAllCachelines_fired(fetch_updateAllCachelines_fired),
    .cachelinesUpdatesResp_ready(fetch_cachelinesUpdatesResp_ready),
    .cachelinesUpdatesResp_fired(fetch_cachelinesUpdatesResp_fired)
  );
  core_Anon decode ( // @[core.scala 38:22]
    .clock(decode_clock),
    .reset(decode_reset),
    .fromFetch_ready(decode_fromFetch_ready),
    .fromFetch_fired(decode_fromFetch_fired),
    .fromFetch_pc(decode_fromFetch_pc),
    .fromFetch_instruction(decode_fromFetch_instruction),
    .fromFetch_expected_valid(decode_fromFetch_expected_valid),
    .fromFetch_expected_pc(decode_fromFetch_expected_pc),
    .toExec_ready(decode_toExec_ready),
    .toExec_fired(decode_toExec_fired),
    .toExec_instruction(decode_toExec_instruction),
    .toExec_pc(decode_toExec_pc),
    .toExec_PRFDest(decode_toExec_PRFDest),
    .toExec_rs1Addr(decode_toExec_rs1Addr),
    .toExec_rs1Ready(decode_toExec_rs1Ready),
    .toExec_rs2Addr(decode_toExec_rs2Addr),
    .toExec_rs2Ready(decode_toExec_rs2Ready),
    .toExec_branchMask(decode_toExec_branchMask),
    .writeBackResult_fired(decode_writeBackResult_fired),
    .writeBackResult_instruction(decode_writeBackResult_instruction),
    .writeBackResult_rdAddr(decode_writeBackResult_rdAddr),
    .writeBackResult_PRFDest(decode_writeBackResult_PRFDest),
    .writeBackResult_data(decode_writeBackResult_data),
    .writeAddrPRF_exec1Addr(decode_writeAddrPRF_exec1Addr),
    .writeAddrPRF_exec2Addr(decode_writeAddrPRF_exec2Addr),
    .writeAddrPRF_exec3Addr(decode_writeAddrPRF_exec3Addr),
    .writeAddrPRF_exec1Valid(decode_writeAddrPRF_exec1Valid),
    .writeAddrPRF_exec2Valid(decode_writeAddrPRF_exec2Valid),
    .writeAddrPRF_exec3Valid(decode_writeAddrPRF_exec3Valid),
    .jumpAddrWrite_ready(decode_jumpAddrWrite_ready),
    .jumpAddrWrite_fired(decode_jumpAddrWrite_fired),
    .jumpAddrWrite_PRFDest(decode_jumpAddrWrite_PRFDest),
    .jumpAddrWrite_linkAddr(decode_jumpAddrWrite_linkAddr),
    .branchPCs_branchPCReady(decode_branchPCs_branchPCReady),
    .branchPCs_branchPC(decode_branchPCs_branchPC),
    .branchPCs_predictedPCReady(decode_branchPCs_predictedPCReady),
    .branchPCs_predictedPC(decode_branchPCs_predictedPC),
    .branchPCs_branchMask(decode_branchPCs_branchMask),
    .branchEvalIn_fired(decode_branchEvalIn_fired),
    .branchEvalIn_passFail(decode_branchEvalIn_passFail),
    .branchEvalIn_branchMask(decode_branchEvalIn_branchMask),
    .branchEvalIn_targetPC(decode_branchEvalIn_targetPC),
    .interruptedPC(decode_interruptedPC),
    .canTakeInterrupt(decode_canTakeInterrupt)
  );
  storeDataIssue dataQueue ( // @[core.scala 52:25]
    .clock(dataQueue_clock),
    .reset(dataQueue_reset),
    .fromROB_readyNow(dataQueue_fromROB_readyNow),
    .fromBranch_passOrFail(dataQueue_fromBranch_passOrFail),
    .fromBranch_robAddr(dataQueue_fromBranch_robAddr),
    .fromBranch_valid(dataQueue_fromBranch_valid),
    .fromDecode_ready(dataQueue_fromDecode_ready),
    .fromDecode_valid(dataQueue_fromDecode_valid),
    .fromDecode_rs2Addr(dataQueue_fromDecode_rs2Addr),
    .fromDecode_branchMask(dataQueue_fromDecode_branchMask),
    .toPRF_valid(dataQueue_toPRF_valid),
    .toPRF_rs2Addr(dataQueue_toPRF_rs2Addr),
    .robMapUpdate_valid(dataQueue_robMapUpdate_valid),
    .robMapUpdate_robAddr(dataQueue_robMapUpdate_robAddr)
  );
  rob rob ( // @[core.scala 53:19]
    .clock(rob_clock),
    .reset(rob_reset),
    .allocate_ready(rob_allocate_ready),
    .allocate_fired(rob_allocate_fired),
    .allocate_pc(rob_allocate_pc),
    .allocate_instruction(rob_allocate_instruction),
    .allocate_prfDest(rob_allocate_prfDest),
    .allocate_robAddr(rob_allocate_robAddr),
    .allocate_isReady(rob_allocate_isReady),
    .commit_ready(rob_commit_ready),
    .commit_fired(rob_commit_fired),
    .commit_prfDest(rob_commit_prfDest),
    .commit_instruction(rob_commit_instruction),
    .commit_exceptionOccurred(rob_commit_exceptionOccurred),
    .commit_mtval(rob_commit_mtval),
    .commit_isStore(rob_commit_isStore),
    .commit_is_fence(rob_commit_is_fence),
    .commit_robAddr(rob_commit_robAddr),
    .branch_valid(rob_branch_valid),
    .branch_pass(rob_branch_pass),
    .branch_robAddr(rob_branch_robAddr),
    .execPorts_0_robAddr(rob_execPorts_0_robAddr),
    .execPorts_0_mtval(rob_execPorts_0_mtval),
    .execPorts_0_valid(rob_execPorts_0_valid),
    .execPorts_1_robAddr(rob_execPorts_1_robAddr),
    .execPorts_1_valid(rob_execPorts_1_valid),
    .execPorts_2_robAddr(rob_execPorts_2_robAddr),
    .execPorts_2_valid(rob_execPorts_2_valid),
    .execPorts_3_robAddr(rob_execPorts_3_robAddr),
    .execPorts_3_valid(rob_execPorts_3_valid)
  );
  scheduler scheduler ( // @[core.scala 54:25]
    .clock(scheduler_clock),
    .reset(scheduler_reset),
    .allocate_ready(scheduler_allocate_ready),
    .allocate_fired(scheduler_allocate_fired),
    .allocate_instruction(scheduler_allocate_instruction),
    .allocate_branchMask(scheduler_allocate_branchMask),
    .allocate_rs1_ready(scheduler_allocate_rs1_ready),
    .allocate_rs1_prfAddr(scheduler_allocate_rs1_prfAddr),
    .allocate_rs2_ready(scheduler_allocate_rs2_ready),
    .allocate_rs2_prfAddr(scheduler_allocate_rs2_prfAddr),
    .allocate_prfDest(scheduler_allocate_prfDest),
    .allocate_robAddr(scheduler_allocate_robAddr),
    .release_ready(scheduler_release_ready),
    .release_fired(scheduler_release_fired),
    .release_instruction(scheduler_release_instruction),
    .release_branchMask(scheduler_release_branchMask),
    .release_rs1prfAddr(scheduler_release_rs1prfAddr),
    .release_rs2prfAddr(scheduler_release_rs2prfAddr),
    .release_prfDest(scheduler_release_prfDest),
    .release_robAddr(scheduler_release_robAddr),
    .wakeUpExt_0_valid(scheduler_wakeUpExt_0_valid),
    .wakeUpExt_0_prfAddr(scheduler_wakeUpExt_0_prfAddr),
    .wakeUpExt_1_valid(scheduler_wakeUpExt_1_valid),
    .wakeUpExt_1_prfAddr(scheduler_wakeUpExt_1_prfAddr),
    .branchOps_valid(scheduler_branchOps_valid),
    .branchOps_branchMask(scheduler_branchOps_branchMask),
    .branchOps_passed(scheduler_branchOps_passed),
    .memoryReady(scheduler_memoryReady),
    .multuplyAndDivideReady(scheduler_multuplyAndDivideReady),
    .instrRetired_valid(scheduler_instrRetired_valid),
    .instrRetired_prfAddr(scheduler_instrRetired_prfAddr)
  );
  core_Anon_1 memAccess ( // @[core.scala 55:25]
    .clock(memAccess_clock),
    .reset(memAccess_reset),
    .peripheral_AWADDR(memAccess_peripheral_AWADDR),
    .peripheral_AWLEN(memAccess_peripheral_AWLEN),
    .peripheral_AWSIZE(memAccess_peripheral_AWSIZE),
    .peripheral_AWVALID(memAccess_peripheral_AWVALID),
    .peripheral_AWREADY(memAccess_peripheral_AWREADY),
    .peripheral_WDATA(memAccess_peripheral_WDATA),
    .peripheral_WSTRB(memAccess_peripheral_WSTRB),
    .peripheral_WLAST(memAccess_peripheral_WLAST),
    .peripheral_WVALID(memAccess_peripheral_WVALID),
    .peripheral_WREADY(memAccess_peripheral_WREADY),
    .peripheral_BVALID(memAccess_peripheral_BVALID),
    .peripheral_BREADY(memAccess_peripheral_BREADY),
    .peripheral_ARADDR(memAccess_peripheral_ARADDR),
    .peripheral_ARLEN(memAccess_peripheral_ARLEN),
    .peripheral_ARSIZE(memAccess_peripheral_ARSIZE),
    .peripheral_ARVALID(memAccess_peripheral_ARVALID),
    .peripheral_ARREADY(memAccess_peripheral_ARREADY),
    .peripheral_RDATA(memAccess_peripheral_RDATA),
    .peripheral_RLAST(memAccess_peripheral_RLAST),
    .peripheral_RVALID(memAccess_peripheral_RVALID),
    .peripheral_RREADY(memAccess_peripheral_RREADY),
    .branchOps_valid(memAccess_branchOps_valid),
    .branchOps_branchMask(memAccess_branchOps_branchMask),
    .branchOps_passed(memAccess_branchOps_passed),
    .writeDataIn_valid(memAccess_writeDataIn_valid),
    .writeDataIn_data(memAccess_writeDataIn_data),
    .responseOut_valid(memAccess_responseOut_valid),
    .responseOut_prfDest(memAccess_responseOut_prfDest),
    .responseOut_robAddr(memAccess_responseOut_robAddr),
    .responseOut_result(memAccess_responseOut_result),
    .responseOut_instruction(memAccess_responseOut_instruction),
    .request_valid(memAccess_request_valid),
    .request_address(memAccess_request_address),
    .request_instruction(memAccess_request_instruction),
    .request_branchMask(memAccess_request_branchMask),
    .request_robAddr(memAccess_request_robAddr),
    .request_prfDest(memAccess_request_prfDest),
    .dPort_AWADDR(memAccess_dPort_AWADDR),
    .dPort_AWLEN(memAccess_dPort_AWLEN),
    .dPort_AWSIZE(memAccess_dPort_AWSIZE),
    .dPort_AWVALID(memAccess_dPort_AWVALID),
    .dPort_AWREADY(memAccess_dPort_AWREADY),
    .dPort_WDATA(memAccess_dPort_WDATA),
    .dPort_WSTRB(memAccess_dPort_WSTRB),
    .dPort_WLAST(memAccess_dPort_WLAST),
    .dPort_WVALID(memAccess_dPort_WVALID),
    .dPort_WREADY(memAccess_dPort_WREADY),
    .dPort_BVALID(memAccess_dPort_BVALID),
    .dPort_BREADY(memAccess_dPort_BREADY),
    .dPort_ARADDR(memAccess_dPort_ARADDR),
    .dPort_ARVALID(memAccess_dPort_ARVALID),
    .dPort_ARREADY(memAccess_dPort_ARREADY),
    .dPort_RDATA(memAccess_dPort_RDATA),
    .dPort_RLAST(memAccess_dPort_RLAST),
    .dPort_RVALID(memAccess_dPort_RVALID),
    .dPort_RREADY(memAccess_dPort_RREADY),
    .writeCommit_ready(memAccess_writeCommit_ready),
    .writeCommit_fired(memAccess_writeCommit_fired),
    .canAllocate(memAccess_canAllocate),
    .initiateFence(memAccess_initiateFence),
    .fenceInstructions_ready(memAccess_fenceInstructions_ready),
    .fenceInstructions_fired(memAccess_fenceInstructions_fired)
  );
  PRF prf ( // @[core.scala 119:19]
    .clock(prf_clock),
    .reset(prf_reset),
    .w1_addr(prf_w1_addr),
    .w1_data(prf_w1_data),
    .w1_en(prf_w1_en),
    .w2_addr(prf_w2_addr),
    .w2_data(prf_w2_data),
    .w2_en(prf_w2_en),
    .w3_addr(prf_w3_addr),
    .w3_data(prf_w3_data),
    .w3_en(prf_w3_en),
    .w4_addr(prf_w4_addr),
    .w4_data(prf_w4_data),
    .w4_en(prf_w4_en),
    .execRead_valid(prf_execRead_valid),
    .execRead_instruction(prf_execRead_instruction),
    .execRead_branchmask(prf_execRead_branchmask),
    .execRead_rs1Addr(prf_execRead_rs1Addr),
    .execRead_rs2Addr(prf_execRead_rs2Addr),
    .execRead_robAddr(prf_execRead_robAddr),
    .execRead_prfDest(prf_execRead_prfDest),
    .toExec_valid(prf_toExec_valid),
    .toExec_instruction(prf_toExec_instruction),
    .toExec_branchmask(prf_toExec_branchmask),
    .toExec_rs1Addr(prf_toExec_rs1Addr),
    .toExec_rs1Data(prf_toExec_rs1Data),
    .toExec_rs2Addr(prf_toExec_rs2Addr),
    .toExec_rs2Data(prf_toExec_rs2Data),
    .toExec_robAddr(prf_toExec_robAddr),
    .toExec_prfDest(prf_toExec_prfDest),
    .fromStore_valid(prf_fromStore_valid),
    .fromStore_rs2Addr(prf_fromStore_rs2Addr),
    .toStore_valid(prf_toStore_valid),
    .toStore_rs2Data(prf_toStore_rs2Data),
    .branchCheck_pass(prf_branchCheck_pass),
    .branchCheck_branchmask(prf_branchCheck_branchmask),
    .branchCheck_valid(prf_branchCheck_valid)
  );
  assign iPort_AWID = 1'h0; // @[core.scala 22:9]
  assign iPort_AWADDR = 32'h0; // @[core.scala 22:9]
  assign iPort_AWLEN = 8'h0; // @[core.scala 22:9]
  assign iPort_AWSIZE = 3'h0; // @[core.scala 22:9]
  assign iPort_AWBURST = 2'h1; // @[core.scala 22:9]
  assign iPort_AWLOCK = 1'h0; // @[core.scala 22:9]
  assign iPort_AWCACHE = 4'h2; // @[core.scala 22:9]
  assign iPort_AWPROT = 3'h0; // @[core.scala 22:9]
  assign iPort_AWQOS = 4'h0; // @[core.scala 22:9]
  assign iPort_AWVALID = 1'h0; // @[core.scala 22:9]
  assign iPort_WDATA = 32'h0; // @[core.scala 22:9]
  assign iPort_WSTRB = 4'h0; // @[core.scala 22:9]
  assign iPort_WLAST = 1'h0; // @[core.scala 22:9]
  assign iPort_WVALID = 1'h0; // @[core.scala 22:9]
  assign iPort_BREADY = 1'h0; // @[core.scala 22:9]
  assign iPort_ARID = 1'h0; // @[core.scala 22:9]
  assign iPort_ARADDR = icache_lowLevelMem_ARADDR; // @[core.scala 22:9]
  assign iPort_ARLEN = 8'h3; // @[core.scala 22:9]
  assign iPort_ARSIZE = 3'h2; // @[core.scala 22:9]
  assign iPort_ARBURST = 2'h1; // @[core.scala 22:9]
  assign iPort_ARLOCK = 1'h0; // @[core.scala 22:9]
  assign iPort_ARCACHE = 4'h2; // @[core.scala 22:9]
  assign iPort_ARPROT = 3'h0; // @[core.scala 22:9]
  assign iPort_ARQOS = 4'h0; // @[core.scala 22:9]
  assign iPort_ARVALID = icache_lowLevelMem_ARVALID; // @[core.scala 22:9]
  assign iPort_RREADY = icache_lowLevelMem_RREADY; // @[core.scala 22:9]
  assign dPort_AWID = 1'h0; // @[core.scala 800:9]
  assign dPort_AWADDR = memAccess_dPort_AWADDR; // @[core.scala 800:9]
  assign dPort_AWLEN = memAccess_dPort_AWLEN; // @[core.scala 800:9]
  assign dPort_AWSIZE = memAccess_dPort_AWSIZE; // @[core.scala 800:9]
  assign dPort_AWBURST = 2'h1; // @[core.scala 800:9]
  assign dPort_AWLOCK = 1'h0; // @[core.scala 800:9]
  assign dPort_AWCACHE = 4'h2; // @[core.scala 800:9]
  assign dPort_AWPROT = 3'h0; // @[core.scala 800:9]
  assign dPort_AWQOS = 4'h0; // @[core.scala 800:9]
  assign dPort_AWVALID = memAccess_dPort_AWVALID; // @[core.scala 800:9]
  assign dPort_WDATA = memAccess_dPort_WDATA; // @[core.scala 800:9]
  assign dPort_WSTRB = memAccess_dPort_WSTRB; // @[core.scala 800:9]
  assign dPort_WLAST = memAccess_dPort_WLAST; // @[core.scala 800:9]
  assign dPort_WVALID = memAccess_dPort_WVALID; // @[core.scala 800:9]
  assign dPort_BREADY = memAccess_dPort_BREADY; // @[core.scala 800:9]
  assign dPort_ARID = 1'h0; // @[core.scala 800:9]
  assign dPort_ARADDR = memAccess_dPort_ARADDR; // @[core.scala 800:9]
  assign dPort_ARLEN = 8'hf; // @[core.scala 800:9]
  assign dPort_ARSIZE = 3'h2; // @[core.scala 800:9]
  assign dPort_ARBURST = 2'h1; // @[core.scala 800:9]
  assign dPort_ARLOCK = 1'h0; // @[core.scala 800:9]
  assign dPort_ARCACHE = 4'h2; // @[core.scala 800:9]
  assign dPort_ARPROT = 3'h0; // @[core.scala 800:9]
  assign dPort_ARQOS = 4'h0; // @[core.scala 800:9]
  assign dPort_ARVALID = memAccess_dPort_ARVALID; // @[core.scala 800:9]
  assign dPort_RREADY = memAccess_dPort_RREADY; // @[core.scala 800:9]
  assign peripheral_AWID = 1'h0; // @[core.scala 801:14]
  assign peripheral_AWADDR = memAccess_peripheral_AWADDR; // @[core.scala 801:14]
  assign peripheral_AWLEN = memAccess_peripheral_AWLEN; // @[core.scala 801:14]
  assign peripheral_AWSIZE = memAccess_peripheral_AWSIZE; // @[core.scala 801:14]
  assign peripheral_AWBURST = 2'h1; // @[core.scala 801:14]
  assign peripheral_AWLOCK = 1'h0; // @[core.scala 801:14]
  assign peripheral_AWCACHE = 4'h2; // @[core.scala 801:14]
  assign peripheral_AWPROT = 3'h0; // @[core.scala 801:14]
  assign peripheral_AWQOS = 4'h0; // @[core.scala 801:14]
  assign peripheral_AWVALID = memAccess_peripheral_AWVALID; // @[core.scala 801:14]
  assign peripheral_WDATA = memAccess_peripheral_WDATA; // @[core.scala 801:14]
  assign peripheral_WSTRB = memAccess_peripheral_WSTRB; // @[core.scala 801:14]
  assign peripheral_WLAST = memAccess_peripheral_WLAST; // @[core.scala 801:14]
  assign peripheral_WVALID = memAccess_peripheral_WVALID; // @[core.scala 801:14]
  assign peripheral_BREADY = memAccess_peripheral_BREADY; // @[core.scala 801:14]
  assign peripheral_ARID = 1'h0; // @[core.scala 801:14]
  assign peripheral_ARADDR = memAccess_peripheral_ARADDR; // @[core.scala 801:14]
  assign peripheral_ARLEN = memAccess_peripheral_ARLEN; // @[core.scala 801:14]
  assign peripheral_ARSIZE = memAccess_peripheral_ARSIZE; // @[core.scala 801:14]
  assign peripheral_ARBURST = 2'h1; // @[core.scala 801:14]
  assign peripheral_ARLOCK = 1'h0; // @[core.scala 801:14]
  assign peripheral_ARCACHE = 4'h2; // @[core.scala 801:14]
  assign peripheral_ARPROT = 3'h0; // @[core.scala 801:14]
  assign peripheral_ARQOS = 4'h0; // @[core.scala 801:14]
  assign peripheral_ARVALID = memAccess_peripheral_ARVALID; // @[core.scala 801:14]
  assign peripheral_RREADY = memAccess_peripheral_RREADY; // @[core.scala 801:14]
  assign core_sample0 = decode_fromFetch_expected_valid; // @[core.scala 949:16]
  assign core_sample1 = decode_fromFetch_expected_pc[30]; // @[core.scala 950:47]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_fromFetch_req_valid = fetch_cache_req_valid; // @[core.scala 30:24]
  assign icache_fromFetch_req_bits = {32'h0,fetch_cache_req_bits[31:0]}; // @[Cat.scala 33:92]
  assign icache_fromFetch_resp_ready = fetch_cache_resp_ready; // @[core.scala 32:20]
  assign icache_updateAllCachelines_fired = memAccess_fenceInstructions_ready & icache_updateAllCachelines_ready; // @[core.scala 855:45]
  assign icache_cachelinesUpdatesResp_fired = icache_cachelinesUpdatesResp_ready & fetch_cachelinesUpdatesResp_ready; // @[core.scala 865:46]
  assign icache_lowLevelMem_ARREADY = iPort_ARREADY; // @[core.scala 22:9]
  assign icache_lowLevelMem_RDATA = iPort_RDATA; // @[core.scala 22:9]
  assign icache_lowLevelMem_RLAST = iPort_RLAST; // @[core.scala 22:9]
  assign icache_lowLevelMem_RVALID = iPort_RVALID; // @[core.scala 22:9]
  assign fetch_clock = clock;
  assign fetch_reset = reset;
  assign fetch_cache_req_ready = icache_fromFetch_req_ready; // @[core.scala 30:24]
  assign fetch_cache_resp_valid = icache_fromFetch_resp_valid; // @[core.scala 32:20]
  assign fetch_cache_resp_bits = icache_fromFetch_resp_bits; // @[core.scala 32:20]
  assign fetch_toDecode_fired = ~(interruptInjectStatus == 2'h0 | interruptInjectStatus == 2'h1 & ~_T_231) ? 1'h0 :
    decode_fromFetch_ready & fetch_toDecode_ready & _fetch_toDecode_fired_T_3; // @[core.scala 1068:126 1070:26 44:7]
  assign fetch_toDecode_expected_valid = decode_fromFetch_expected_valid; // @[core.scala 48:27]
  assign fetch_toDecode_expected_pc = decode_fromFetch_expected_pc; // @[core.scala 48:27]
  assign fetch_branchRes_fired = branchEvals_valid; // @[core.scala 680:50]
  assign fetch_branchRes_branchTaken = fetch_branchRes_branchTaken_REG; // @[core.scala 676:31]
  assign fetch_branchRes_pc = fetch_branchRes_pc_REG; // @[core.scala 678:22]
  assign fetch_branchRes_pcAfterBrnach = branchEvals_nextPC; // @[core.scala 679:33]
  assign fetch_carryOutFence_fired = fetch_carryOutFence_ready; // @[core.scala 857:29]
  assign fetch_updateAllCachelines_fired = fetch_updateAllCachelines_ready; // @[core.scala 862:35]
  assign fetch_cachelinesUpdatesResp_fired = icache_cachelinesUpdatesResp_ready & fetch_cachelinesUpdatesResp_ready; // @[core.scala 865:46]
  assign decode_clock = clock;
  assign decode_reset = reset;
  assign decode_fromFetch_fired = ~(interruptInjectStatus == 2'h0 | interruptInjectStatus == 2'h1 & ~_T_231) ? 1'h0 :
    decode_fromFetch_ready & fetch_toDecode_ready & _fetch_toDecode_fired_T_3; // @[core.scala 1068:126 1071:28 44:7]
  assign decode_fromFetch_pc = fetch_toDecode_pc; // @[core.scala 50:23]
  assign decode_fromFetch_instruction = _GEN_299[31:0];
  assign decode_toExec_fired = decode_toExec_ready & rob_allocate_ready & scheduler_allocate_ready & (
    decode_toExec_instruction[6:4] != 3'h2 | dataQueue_fromDecode_ready); // @[core.scala 79:81]
  assign decode_writeBackResult_fired = rob_commit_ready & (memAccess_writeCommit_ready | rob_commit_instruction[6:4]
     != 3'h2); // @[core.scala 687:60]
  assign decode_writeBackResult_instruction = _GEN_300[31:0];
  assign decode_writeBackResult_rdAddr = rob_commit_instruction[11:7]; // @[core.scala 685:58]
  assign decode_writeBackResult_PRFDest = rob_commit_prfDest; // @[core.scala 682:34]
  assign decode_writeBackResult_data = rob_commit_mtval; // @[core.scala 869:31]
  assign decode_writeAddrPRF_exec1Addr = scheduler_instrRetired_prfAddr; // @[core.scala 690:33]
  assign decode_writeAddrPRF_exec2Addr = memAccess_responseOut_prfDest; // @[core.scala 692:33]
  assign decode_writeAddrPRF_exec3Addr = extnMResponse_prfDest; // @[core.scala 693:33]
  assign decode_writeAddrPRF_exec1Valid = scheduler_instrRetired_valid; // @[core.scala 691:34]
  assign decode_writeAddrPRF_exec2Valid = memAccess_responseOut_valid & _T_181; // @[core.scala 694:65]
  assign decode_writeAddrPRF_exec3Valid = extnMResponse_valid & _T_184; // @[core.scala 695:57]
  assign decode_jumpAddrWrite_fired = decode_jumpAddrWrite_ready; // @[core.scala 761:30]
  assign decode_branchEvalIn_fired = branchEvals_valid; // @[core.scala 700:58]
  assign decode_branchEvalIn_passFail = branchEvals_passed; // @[core.scala 698:32]
  assign decode_branchEvalIn_branchMask = branchEvals_branchMask; // @[core.scala 697:34]
  assign decode_branchEvalIn_targetPC = branchEvals_nextPC; // @[core.scala 699:32]
  assign decode_interruptedPC = lastBranchExecPC; // @[core.scala 1007:24]
  assign dataQueue_clock = clock;
  assign dataQueue_reset = reset;
  assign dataQueue_fromROB_readyNow = memAccess_writeCommit_fired; // @[core.scala 780:30]
  assign dataQueue_fromBranch_passOrFail = branchEvals_passed; // @[core.scala 517:20 65:23]
  assign dataQueue_fromBranch_robAddr = branchEvals_robAddr; // @[core.scala 773:32]
  assign dataQueue_fromBranch_valid = branchEvals_valid; // @[core.scala 516:19 65:23]
  assign dataQueue_fromDecode_valid = branchEvals_valid ? _GEN_3 : scheduler_allocate_fired & decode_toExec_instruction[
    6:4] == 3'h2; // @[core.scala 100:25 98:30]
  assign dataQueue_fromDecode_rs2Addr = decode_toExec_rs2Addr; // @[core.scala 96:32]
  assign dataQueue_fromDecode_branchMask = branchEvals_valid ? _scheduler_allocate_branchMask_T :
    decode_toExec_branchMask; // @[core.scala 100:25 102:36 94:35]
  assign dataQueue_robMapUpdate_valid = rob_allocate_fired; // @[core.scala 778:32]
  assign dataQueue_robMapUpdate_robAddr = rob_allocate_robAddr; // @[core.scala 777:34]
  assign rob_clock = clock;
  assign rob_reset = reset;
  assign rob_allocate_fired = branchEvals_valid ? _GEN_2 : decode_toExec_ready & rob_allocate_ready &
    scheduler_allocate_ready & (decode_toExec_instruction[6:4] != 3'h2 | dataQueue_fromDecode_ready); // @[core.scala 100:25 79:7]
  assign rob_allocate_pc = decode_toExec_pc; // @[core.scala 82:19]
  assign rob_allocate_instruction = decode_toExec_instruction; // @[core.scala 83:28]
  assign rob_allocate_prfDest = decode_toExec_PRFDest; // @[core.scala 84:24]
  assign rob_allocate_isReady = 5'h3 == decode_toExec_instruction[6:2] | 5'h5 == decode_toExec_instruction[6:2] | 5'hd
     == decode_toExec_instruction[6:2]; // @[core.scala 77:125]
  assign rob_commit_fired = rob_commit_ready & (memAccess_writeCommit_ready | rob_commit_instruction[6:4] != 3'h2); // @[core.scala 687:60]
  assign rob_branch_valid = branchEvals_valid; // @[core.scala 704:20]
  assign rob_branch_pass = branchEvals_passed; // @[core.scala 702:19]
  assign rob_branch_robAddr = branchEvals_robAddr; // @[core.scala 703:22]
  assign rob_execPorts_0_robAddr = singleCycleArithmeticResponse_robAddr; // @[core.scala 728:22]
  assign rob_execPorts_0_mtval = rob_execPorts_0_mtval_REG; // @[core.scala 712:26]
  assign rob_execPorts_0_valid = singleCycleArithmeticResponse_valid; // @[core.scala 729:20]
  assign rob_execPorts_1_robAddr = branchEvals_robAddr; // @[core.scala 728:22]
  assign rob_execPorts_1_valid = branchEvals_valid; // @[core.scala 729:20]
  assign rob_execPorts_2_robAddr = memAccess_responseOut_robAddr; // @[core.scala 728:22]
  assign rob_execPorts_2_valid = memAccess_responseOut_valid; // @[core.scala 729:20]
  assign rob_execPorts_3_robAddr = extnMResponse_robAddr; // @[core.scala 728:22]
  assign rob_execPorts_3_valid = extnMResponse_valid; // @[core.scala 729:20]
  assign scheduler_clock = clock;
  assign scheduler_reset = reset;
  assign scheduler_allocate_fired = branchEvals_valid ? _GEN_1 : _GEN_0; // @[core.scala 100:25]
  assign scheduler_allocate_instruction = decode_toExec_instruction; // @[core.scala 86:34]
  assign scheduler_allocate_branchMask = branchEvals_valid ? _scheduler_allocate_branchMask_T : decode_toExec_branchMask
    ; // @[core.scala 100:25 101:34 87:33]
  assign scheduler_allocate_rs1_ready = wakeUps_2_valid ? _GEN_17 : _GEN_15; // @[core.scala 111:24]
  assign scheduler_allocate_rs1_prfAddr = decode_toExec_rs1Addr; // @[core.scala 89:34]
  assign scheduler_allocate_rs2_ready = wakeUps_2_valid ? _GEN_18 : _GEN_16; // @[core.scala 111:24]
  assign scheduler_allocate_rs2_prfAddr = decode_toExec_rs2Addr; // @[core.scala 91:34]
  assign scheduler_allocate_prfDest = decode_toExec_PRFDest; // @[core.scala 92:30]
  assign scheduler_allocate_robAddr = rob_allocate_robAddr; // @[core.scala 93:30]
  assign scheduler_release_fired = scheduler_release_ready & _scheduler_release_fired_T_5; // @[core.scala 121:29]
  assign scheduler_wakeUpExt_0_valid = memAccess_responseOut_valid & |memAccess_responseOut_instruction[11:7]; // @[core.scala 752:33]
  assign scheduler_wakeUpExt_0_prfAddr = memAccess_responseOut_prfDest; // @[core.scala 71:21 757:20]
  assign scheduler_wakeUpExt_1_valid = extnMResponse_valid & |extnResponseInstruction[11:7]; // @[core.scala 753:25]
  assign scheduler_wakeUpExt_1_prfAddr = extnMResponse_prfDest; // @[core.scala 71:21 757:20]
  assign scheduler_branchOps_valid = branchEvals_valid; // @[core.scala 516:19 65:23]
  assign scheduler_branchOps_branchMask = branchEvals_branchMask; // @[core.scala 65:23 518:24]
  assign scheduler_branchOps_passed = branchEvals_passed; // @[core.scala 517:20 65:23]
  assign scheduler_memoryReady = memAccess_canAllocate; // @[core.scala 706:25]
  assign scheduler_multuplyAndDivideReady = mExtensionReady; // @[core.scala 707:36]
  assign memAccess_clock = clock;
  assign memAccess_reset = reset;
  assign memAccess_peripheral_AWREADY = peripheral_AWREADY; // @[core.scala 801:14]
  assign memAccess_peripheral_WREADY = peripheral_WREADY; // @[core.scala 801:14]
  assign memAccess_peripheral_BVALID = peripheral_BVALID; // @[core.scala 801:14]
  assign memAccess_peripheral_ARREADY = peripheral_ARREADY; // @[core.scala 801:14]
  assign memAccess_peripheral_RDATA = peripheral_RDATA; // @[core.scala 801:14]
  assign memAccess_peripheral_RLAST = peripheral_RLAST; // @[core.scala 801:14]
  assign memAccess_peripheral_RVALID = peripheral_RVALID; // @[core.scala 801:14]
  assign memAccess_branchOps_valid = branchEvals_valid; // @[core.scala 516:19 65:23]
  assign memAccess_branchOps_branchMask = branchEvals_branchMask; // @[core.scala 65:23 518:24]
  assign memAccess_branchOps_passed = branchEvals_passed; // @[core.scala 517:20 65:23]
  assign memAccess_writeDataIn_valid = prf_toStore_valid; // @[core.scala 783:31]
  assign memAccess_writeDataIn_data = prf_toStore_rs2Data; // @[core.scala 782:30]
  assign memAccess_request_valid = memoryRequest_valid; // @[core.scala 182:21]
  assign memAccess_request_address = memoryRequest_address; // @[core.scala 182:21]
  assign memAccess_request_instruction = memoryRequest_instruction; // @[core.scala 182:21]
  assign memAccess_request_branchMask = memoryRequest_branchMask; // @[core.scala 182:21]
  assign memAccess_request_robAddr = memoryRequest_robAddr; // @[core.scala 182:21]
  assign memAccess_request_prfDest = memoryRequest_prfDest; // @[core.scala 182:21]
  assign memAccess_dPort_AWREADY = dPort_AWREADY; // @[core.scala 800:9]
  assign memAccess_dPort_WREADY = dPort_WREADY; // @[core.scala 800:9]
  assign memAccess_dPort_BVALID = dPort_BVALID; // @[core.scala 800:9]
  assign memAccess_dPort_ARREADY = dPort_ARREADY; // @[core.scala 800:9]
  assign memAccess_dPort_RDATA = dPort_RDATA; // @[core.scala 800:9]
  assign memAccess_dPort_RLAST = dPort_RLAST; // @[core.scala 800:9]
  assign memAccess_dPort_RVALID = dPort_RVALID; // @[core.scala 800:9]
  assign memAccess_writeCommit_fired = memAccess_writeCommit_ready & rob_commit_instruction[6:4] == 3'h2 &
    rob_commit_fired; // @[core.scala 785:109]
  assign memAccess_initiateFence = REG_1 | _GEN_244; // @[core.scala 874:131 875:29]
  assign memAccess_fenceInstructions_fired = memAccess_fenceInstructions_ready & icache_updateAllCachelines_ready; // @[core.scala 855:45]
  assign prf_clock = clock;
  assign prf_reset = reset;
  assign prf_w1_addr = singleCycleArithmeticResponse_prfDest; // @[core.scala 740:20]
  assign prf_w1_data = singleCycleArithmeticResponse_result; // @[core.scala 741:20]
  assign prf_w1_en = singleCycleArithmeticResponse_valid & REG; // @[core.scala 733:119]
  assign prf_w2_addr = decode_jumpAddrWrite_PRFDest; // @[core.scala 740:20]
  assign prf_w2_data = decode_jumpAddrWrite_linkAddr; // @[core.scala 741:20]
  assign prf_w2_en = decode_jumpAddrWrite_ready; // @[core.scala 742:18]
  assign prf_w3_addr = memAccess_responseOut_prfDest; // @[core.scala 740:20]
  assign prf_w3_data = memAccess_responseOut_result; // @[core.scala 741:20]
  assign prf_w3_en = memAccess_responseOut_valid & _T_181; // @[core.scala 735:95]
  assign prf_w4_addr = extnMResponse_prfDest; // @[core.scala 740:20]
  assign prf_w4_data = extnMResponse_result; // @[core.scala 741:20]
  assign prf_w4_en = extnMResponse_valid & _T_184; // @[core.scala 736:71]
  assign prf_execRead_valid = scheduler_release_instruction[4:2] == 3'h2 ? 1'h0 : _GEN_21; // @[core.scala 880:{63,84}]
  assign prf_execRead_instruction = scheduler_release_instruction; // @[core.scala 125:28]
  assign prf_execRead_branchmask = scheduler_release_branchMask; // @[core.scala 126:27]
  assign prf_execRead_rs1Addr = scheduler_release_rs1prfAddr; // @[core.scala 127:24]
  assign prf_execRead_rs2Addr = scheduler_release_rs2prfAddr; // @[core.scala 128:24]
  assign prf_execRead_robAddr = {{2'd0}, scheduler_release_robAddr}; // @[core.scala 129:24]
  assign prf_execRead_prfDest = scheduler_release_prfDest; // @[core.scala 131:24]
  assign prf_fromStore_valid = prf_fromStore_valid_REG_1; // @[core.scala 770:23]
  assign prf_fromStore_rs2Addr = prf_fromStore_rs2Addr_REG_1; // @[core.scala 769:25]
  assign prf_branchCheck_pass = branchEvals_passed; // @[core.scala 517:20 65:23]
  assign prf_branchCheck_branchmask = branchEvals_branchMask; // @[core.scala 65:23 518:24]
  assign prf_branchCheck_valid = branchEvals_valid; // @[core.scala 516:19 65:23]
  always @(posedge clock) begin
    branchEvals_branchMask <= branchPCs_0_branchMask; // @[core.scala 544:26]
    if (2'h0 == interruptInjectStatus) begin // @[core.scala 1025:33]
      branchEvals_passed <= predictedPCs_0_valid & _GEN_159 == predictedPCs_0_pc; // @[core.scala 598:22]
    end else if (2'h1 == interruptInjectStatus) begin // @[core.scala 1025:33]
      if (decode_canTakeInterrupt) begin // @[core.scala 1033:56]
        if (~branchEvals_valid) begin // @[core.scala 1034:58]
          branchEvals_passed <= _GEN_278;
        end else begin
          branchEvals_passed <= predictedPCs_0_valid & _GEN_159 == predictedPCs_0_pc; // @[core.scala 598:22]
        end
      end else begin
        branchEvals_passed <= predictedPCs_0_valid & _GEN_159 == predictedPCs_0_pc; // @[core.scala 598:22]
      end
    end else begin
      branchEvals_passed <= predictedPCs_0_valid & _GEN_159 == predictedPCs_0_pc; // @[core.scala 598:22]
    end
    if (reset) begin // @[core.scala 509:28]
      branchEvals_valid <= 1'h0; // @[core.scala 509:28]
    end else if (branchEvals_valid) begin // @[core.scala 546:25]
      if (_T) begin // @[core.scala 548:29]
        branchEvals_valid <= 1'h0; // @[core.scala 549:25]
      end else begin
        branchEvals_valid <= branchInstruction_valid; // @[core.scala 542:21]
      end
    end else begin
      branchEvals_valid <= branchInstruction_valid; // @[core.scala 542:21]
    end
    if (division_request_valid & ~(|division_counter)) begin // @[core.scala 426:57]
      extnMResponse_prfDest <= division_request_prfDest; // @[core.scala 427:27]
    end else begin
      extnMResponse_prfDest <= extnMServicing_prfDest; // @[core.scala 352:25]
    end
    if (reset) begin // @[core.scala 211:30]
      extnMResponse_valid <= 1'h0; // @[core.scala 211:30]
    end else if (division_request_valid & ~(|division_counter)) begin // @[core.scala 426:57]
      if (branchEvals_valid) begin // @[core.scala 450:27]
        if (|_T_106 & _T) begin // @[core.scala 451:91]
          extnMResponse_valid <= 1'h0; // @[core.scala 451:113]
        end else begin
          extnMResponse_valid <= division_request_valid; // @[core.scala 447:25]
        end
      end else begin
        extnMResponse_valid <= division_request_valid; // @[core.scala 447:25]
      end
    end else if (branchEvals_valid) begin // @[core.scala 367:25]
      if (_T) begin // @[core.scala 373:29]
        extnMResponse_valid <= _GEN_67;
      end else begin
        extnMResponse_valid <= extnMServicing_valid; // @[core.scala 364:23]
      end
    end else begin
      extnMResponse_valid <= extnMServicing_valid; // @[core.scala 364:23]
    end
    if (division_request_valid & ~(|division_counter)) begin // @[core.scala 426:57]
      extnResponseInstruction <= division_request_instruction; // @[core.scala 448:29]
    end else begin
      extnResponseInstruction <= extnMServicing_instruction; // @[core.scala 365:27]
    end
    mExtensionReady <= reset | _GEN_85; // @[core.scala 117:{32,32}]
    if (reset) begin // @[core.scala 140:39]
      addressGenerationInput_valid <= 1'h0; // @[core.scala 140:39]
    end else if (branchEvals_valid) begin // @[core.scala 156:25]
      if (_T & _T_10) begin // @[core.scala 160:83]
        addressGenerationInput_valid <= 1'h0; // @[core.scala 160:114]
      end else begin
        addressGenerationInput_valid <= prf_toExec_valid & ~(prf_toExec_instruction[6] | prf_toExec_instruction[4]); // @[core.scala 149:32]
      end
    end else begin
      addressGenerationInput_valid <= prf_toExec_valid & ~(prf_toExec_instruction[6] | prf_toExec_instruction[4]); // @[core.scala 149:32]
    end
    if (|prf_toExec_instruction[19:15]) begin // @[core.scala 235:36]
      if (_addressGenerationInput_rs1_T_3) begin // @[Mux.scala 101:16]
        addressGenerationInput_rs1 <= fwdFrom_0_result;
      end else if (_addressGenerationInput_rs1_T_5) begin // @[Mux.scala 101:16]
        addressGenerationInput_rs1 <= fwdBuffers_0_result;
      end else if (_addressGenerationInput_rs1_T_7) begin // @[Mux.scala 101:16]
        addressGenerationInput_rs1 <= fwdBuffers_1_result;
      end else begin
        addressGenerationInput_rs1 <= prf_toExec_rs1Data;
      end
    end else begin
      addressGenerationInput_rs1 <= 64'h0;
    end
    addressGenerationInput_instruction <= prf_toExec_instruction; // @[core.scala 151:38]
    addressGenerationInput_prfDest <= prf_toExec_prfDest; // @[core.scala 152:34]
    addressGenerationInput_robAddr <= prf_toExec_robAddr[3:0]; // @[core.scala 153:34]
    if (branchEvals_valid) begin // @[core.scala 156:25]
      if (|_T_9) begin // @[core.scala 157:62]
        addressGenerationInput_branchMask <= _addressGenerationInput_branchMask_T; // @[core.scala 158:41]
      end else begin
        addressGenerationInput_branchMask <= prf_toExec_branchmask; // @[core.scala 154:37]
      end
    end else begin
      addressGenerationInput_branchMask <= prf_toExec_branchmask; // @[core.scala 154:37]
    end
    if (reset) begin // @[core.scala 163:30]
      memoryRequest_valid <= 1'h0; // @[core.scala 163:30]
    end else if (branchEvals_valid) begin // @[core.scala 175:25]
      if (_T & _T_16) begin // @[core.scala 179:95]
        memoryRequest_valid <= 1'h0; // @[core.scala 179:117]
      end else begin
        memoryRequest_valid <= addressGenerationInput_valid; // @[core.scala 173:23]
      end
    end else begin
      memoryRequest_valid <= addressGenerationInput_valid; // @[core.scala 173:23]
    end
    memoryRequest_address <= _memoryRequest_address_T_15[31:0]; // @[core.scala 164:25]
    memoryRequest_instruction <= addressGenerationInput_instruction; // @[core.scala 170:29]
    if (branchEvals_valid) begin // @[core.scala 175:25]
      if (|_T_15) begin // @[core.scala 176:74]
        memoryRequest_branchMask <= _memoryRequest_branchMask_T; // @[core.scala 177:32]
      end else begin
        memoryRequest_branchMask <= addressGenerationInput_branchMask; // @[core.scala 169:28]
      end
    end else begin
      memoryRequest_branchMask <= addressGenerationInput_branchMask; // @[core.scala 169:28]
    end
    memoryRequest_robAddr <= addressGenerationInput_robAddr; // @[core.scala 172:25]
    memoryRequest_prfDest <= addressGenerationInput_prfDest; // @[core.scala 171:25]
    if (reset) begin // @[core.scala 185:45]
      singleCycleArithmeticRequest_valid <= 1'h0; // @[core.scala 185:45]
    end else if (branchEvals_valid) begin // @[core.scala 286:25]
      if (_T_14) begin // @[core.scala 290:83]
        singleCycleArithmeticRequest_valid <= 1'h0; // @[core.scala 291:42]
      end else begin
        singleCycleArithmeticRequest_valid <= prf_toExec_valid & 3'h4 == _singleCycleArithmeticRequest_valid_T_1 & (
          prf_toExec_instruction[6] | ~prf_toExec_instruction[5] | ~prf_toExec_instruction[25]); // @[core.scala 274:38]
      end
    end else begin
      singleCycleArithmeticRequest_valid <= prf_toExec_valid & 3'h4 == _singleCycleArithmeticRequest_valid_T_1 & (
        prf_toExec_instruction[6] | ~prf_toExec_instruction[5] | ~prf_toExec_instruction[25]); // @[core.scala 274:38]
    end
    if (_addressGenerationInput_rs1_T_1) begin // @[core.scala 279:42]
      if (_addressGenerationInput_rs1_T_3) begin // @[Mux.scala 101:16]
        singleCycleArithmeticRequest_rs1 <= fwdFrom_0_result;
      end else if (_addressGenerationInput_rs1_T_5) begin // @[Mux.scala 101:16]
        singleCycleArithmeticRequest_rs1 <= fwdBuffers_0_result;
      end else if (_addressGenerationInput_rs1_T_7) begin // @[Mux.scala 101:16]
        singleCycleArithmeticRequest_rs1 <= fwdBuffers_1_result;
      end else begin
        singleCycleArithmeticRequest_rs1 <= prf_toExec_rs1Data;
      end
    end else begin
      singleCycleArithmeticRequest_rs1 <= 64'h0;
    end
    if (prf_toExec_instruction[5]) begin // @[core.scala 282:42]
      if (|prf_toExec_instruction[24:20]) begin // @[core.scala 282:80]
        if (_singleCycleArithmeticRequest_rs2_T_5) begin // @[Mux.scala 101:16]
          singleCycleArithmeticRequest_rs2 <= fwdFrom_0_result;
        end else if (_singleCycleArithmeticRequest_rs2_T_7) begin // @[Mux.scala 101:16]
          singleCycleArithmeticRequest_rs2 <= fwdBuffers_0_result;
        end else begin
          singleCycleArithmeticRequest_rs2 <= _singleCycleArithmeticRequest_rs2_T_10;
        end
      end else begin
        singleCycleArithmeticRequest_rs2 <= 64'h0;
      end
    end else begin
      singleCycleArithmeticRequest_rs2 <= arithmeticImm;
    end
    singleCycleArithmeticRequest_instruction <= prf_toExec_instruction; // @[core.scala 276:44]
    singleCycleArithmeticRequest_prfDest <= prf_toExec_prfDest; // @[core.scala 277:40]
    singleCycleArithmeticRequest_robAddr <= prf_toExec_robAddr[3:0]; // @[core.scala 278:40]
    if (branchEvals_valid) begin // @[core.scala 286:25]
      if (|_T_9) begin // @[core.scala 157:62]
        singleCycleArithmeticRequest_branchMask <= _addressGenerationInput_branchMask_T; // @[core.scala 158:41]
      end else begin
        singleCycleArithmeticRequest_branchMask <= prf_toExec_branchmask; // @[core.scala 154:37]
      end
    end else begin
      singleCycleArithmeticRequest_branchMask <= prf_toExec_branchmask; // @[core.scala 275:43]
    end
    if (reset) begin // @[core.scala 195:46]
      singleCycleArithmeticResponse_valid <= 1'h0; // @[core.scala 195:46]
    end else if (branchEvals_valid) begin // @[core.scala 301:25]
      if (_T & |_T_30) begin // @[core.scala 302:101]
        singleCycleArithmeticResponse_valid <= 1'h0; // @[core.scala 303:43]
      end else begin
        singleCycleArithmeticResponse_valid <= singleCycleArithmeticRequest_valid; // @[core.scala 299:39]
      end
    end else begin
      singleCycleArithmeticResponse_valid <= singleCycleArithmeticRequest_valid; // @[core.scala 299:39]
    end
    singleCycleArithmeticResponse_result <= arithmeticResult[63:0]; // @[core.scala 297:40]
    singleCycleArithmeticResponse_prfDest <= singleCycleArithmeticRequest_prfDest; // @[core.scala 296:41]
    singleCycleArithmeticResponse_robAddr <= singleCycleArithmeticRequest_robAddr; // @[core.scala 298:41]
    if (reset) begin // @[core.scala 202:29]
      extnMRequest_valid <= 1'h0; // @[core.scala 202:29]
    end else if (branchEvals_valid) begin // @[core.scala 367:25]
      if (_T) begin // @[core.scala 373:29]
        if (_T_10 & prf_toExec_valid) begin // @[core.scala 376:101]
          extnMRequest_valid <= 1'h0; // @[core.scala 376:107]
        end else begin
          extnMRequest_valid <= _GEN_56;
        end
      end else begin
        extnMRequest_valid <= _GEN_56;
      end
    end else begin
      extnMRequest_valid <= _GEN_56;
    end
    if (_addressGenerationInput_rs1_T_3) begin // @[Mux.scala 101:16]
      extnMRequest_rs1 <= fwdFrom_0_result;
    end else if (_addressGenerationInput_rs1_T_5) begin // @[Mux.scala 101:16]
      extnMRequest_rs1 <= fwdBuffers_0_result;
    end else if (_addressGenerationInput_rs1_T_7) begin // @[Mux.scala 101:16]
      extnMRequest_rs1 <= fwdBuffers_1_result;
    end else begin
      extnMRequest_rs1 <= prf_toExec_rs1Data;
    end
    if (_singleCycleArithmeticRequest_rs2_T_5) begin // @[Mux.scala 101:16]
      extnMRequest_rs2 <= fwdFrom_0_result;
    end else if (_singleCycleArithmeticRequest_rs2_T_7) begin // @[Mux.scala 101:16]
      extnMRequest_rs2 <= fwdBuffers_0_result;
    end else if (_singleCycleArithmeticRequest_rs2_T_9) begin // @[Mux.scala 101:16]
      extnMRequest_rs2 <= fwdBuffers_1_result;
    end else begin
      extnMRequest_rs2 <= prf_toExec_rs2Data;
    end
    extnMRequest_instruction <= prf_toExec_instruction; // @[core.scala 310:28]
    extnMRequest_prfDest <= prf_toExec_prfDest; // @[core.scala 319:24]
    extnMRequest_robAddr <= prf_toExec_robAddr[3:0]; // @[core.scala 320:24]
    if (branchEvals_valid) begin // @[core.scala 367:25]
      if (_T_10) begin // @[core.scala 370:73]
        extnMRequest_branchMask <= _addressGenerationInput_branchMask_T; // @[core.scala 371:11]
      end else begin
        extnMRequest_branchMask <= _GEN_24;
      end
    end else begin
      extnMRequest_branchMask <= _GEN_24;
    end
    if (reset) begin // @[core.scala 204:31]
      extnMServicing_valid <= 1'h0; // @[core.scala 204:31]
    end else if (branchEvals_valid) begin // @[core.scala 367:25]
      if (_T) begin // @[core.scala 373:29]
        if (_T_57 & extnMRequest_valid) begin // @[core.scala 376:101]
          extnMServicing_valid <= 1'h0; // @[core.scala 376:107]
        end else begin
          extnMServicing_valid <= extnMPartialServicing_valid; // @[core.scala 208:18]
        end
      end else begin
        extnMServicing_valid <= extnMPartialServicing_valid; // @[core.scala 208:18]
      end
    end else begin
      extnMServicing_valid <= extnMPartialServicing_valid; // @[core.scala 208:18]
    end
    extnMServicing_instruction <= extnMPartialServicing_instruction; // @[core.scala 208:18]
    extnMServicing_prfDest <= extnMPartialServicing_prfDest; // @[core.scala 208:18]
    extnMServicing_robAddr <= extnMPartialServicing_robAddr; // @[core.scala 208:18]
    if (branchEvals_valid) begin // @[core.scala 367:25]
      if (_T_60) begin // @[core.scala 370:73]
        extnMServicing_branchMask <= _T_58; // @[core.scala 371:11]
      end else begin
        extnMServicing_branchMask <= extnMPartialServicing_branchMask; // @[core.scala 208:18]
      end
    end else begin
      extnMServicing_branchMask <= extnMPartialServicing_branchMask; // @[core.scala 208:18]
    end
    if (reset) begin // @[core.scala 205:38]
      extnMPartialServicing_valid <= 1'h0; // @[core.scala 205:38]
    end else if (extnMRequest_instruction[14]) begin // @[core.scala 209:45]
      extnMPartialServicing_valid <= 1'h0; // @[core.scala 209:75]
    end else begin
      extnMPartialServicing_valid <= extnMRequest_valid; // @[core.scala 207:25]
    end
    extnMPartialServicing_instruction <= extnMRequest_instruction; // @[core.scala 207:25]
    extnMPartialServicing_prfDest <= extnMRequest_prfDest; // @[core.scala 207:25]
    extnMPartialServicing_robAddr <= extnMRequest_robAddr; // @[core.scala 207:25]
    if (branchEvals_valid) begin // @[core.scala 367:25]
      if (_T_57) begin // @[core.scala 370:73]
        extnMPartialServicing_branchMask <= _T_55; // @[core.scala 371:11]
      end else begin
        extnMPartialServicing_branchMask <= extnMRequest_branchMask; // @[core.scala 207:25]
      end
    end else begin
      extnMPartialServicing_branchMask <= extnMRequest_branchMask; // @[core.scala 207:25]
    end
    muls_0 <= _GEN_94 + _muls_0_T; // @[core.scala 343:29]
    muls_1 <= _GEN_108 + _muls_1_T; // @[core.scala 344:28]
    muls_2 <= _GEN_108 + _muls_2_T; // @[core.scala 345:28]
    muls_3 <= _muls_3_T_3 + _muls_3_T_4; // @[core.scala 346:62]
    muls_4 <= _GEN_94 + _muls_4_T; // @[core.scala 347:28]
    muls_5 <= {{32'd0}, narrowMuls_8}; // @[core.scala 348:11]
    extnMResponse_result <= _GEN_120[63:0];
    if (division_request_valid & ~(|division_counter)) begin // @[core.scala 426:57]
      extnMResponse_robAddr <= division_request_robAddr; // @[core.scala 446:27]
    end else begin
      extnMResponse_robAddr <= extnMServicing_robAddr; // @[core.scala 363:25]
    end
    if (reset) begin // @[core.scala 213:25]
      division_request_valid <= 1'h0; // @[core.scala 213:25]
    end else if (branchEvals_valid) begin // @[core.scala 455:25]
      if (_T & _T_107) begin // @[core.scala 461:89]
        division_request_valid <= 1'h0; // @[core.scala 461:114]
      end else if (extnMRequest_valid) begin // @[core.scala 456:30]
        division_request_valid <= _GEN_126;
      end else begin
        division_request_valid <= _GEN_124;
      end
    end else begin
      division_request_valid <= _GEN_124;
    end
    if (extnMRequest_valid & extnMRequest_instruction[14]) begin // @[core.scala 404:67]
      division_request_rs1 <= extnMRequest_rs1; // @[core.scala 413:22]
    end
    if (extnMRequest_valid & extnMRequest_instruction[14]) begin // @[core.scala 404:67]
      division_request_rs2 <= extnMRequest_rs2; // @[core.scala 413:22]
    end
    if (extnMRequest_valid & extnMRequest_instruction[14]) begin // @[core.scala 404:67]
      division_request_instruction <= extnMRequest_instruction; // @[core.scala 413:22]
    end
    if (extnMRequest_valid & extnMRequest_instruction[14]) begin // @[core.scala 404:67]
      division_request_prfDest <= extnMRequest_prfDest; // @[core.scala 413:22]
    end
    if (extnMRequest_valid & extnMRequest_instruction[14]) begin // @[core.scala 404:67]
      division_request_robAddr <= extnMRequest_robAddr; // @[core.scala 413:22]
    end
    if (branchEvals_valid) begin // @[core.scala 455:25]
      if (_T_107) begin // @[core.scala 460:69]
        division_request_branchMask <= _division_request_branchMask_T_1; // @[core.scala 460:99]
      end else if (extnMRequest_valid) begin // @[core.scala 456:30]
        if (_T_57) begin // @[core.scala 457:67]
          division_request_branchMask <= _T_55; // @[core.scala 457:97]
        end else begin
          division_request_branchMask <= _GEN_107;
        end
      end else begin
        division_request_branchMask <= _GEN_107;
      end
    end else begin
      division_request_branchMask <= _GEN_107;
    end
    if (extnMRequest_valid & extnMRequest_instruction[14]) begin // @[core.scala 404:67]
      if (~extnMRequest_instruction[12]) begin // @[core.scala 415:47]
        if (extnMRequest_instruction[3]) begin // @[core.scala 419:48]
          if (extnMRequest_rs1[31]) begin // @[core.scala 420:43]
            division_quotient <= _division_quotient_T_24; // @[core.scala 420:63]
          end else begin
            division_quotient <= _GEN_88;
          end
        end else begin
          division_quotient <= _GEN_88;
        end
      end else begin
        division_quotient <= _GEN_87;
      end
    end else begin
      division_quotient <= _division_quotient_T_13; // @[core.scala 401:21]
    end
    if (extnMRequest_valid & extnMRequest_instruction[14]) begin // @[core.scala 404:67]
      division_remainder <= 65'h0; // @[core.scala 412:24]
    end else begin
      division_remainder <= _division_remainder_T_9; // @[core.scala 400:22]
    end
    if (extnMRequest_valid & extnMRequest_instruction[14]) begin // @[core.scala 404:67]
      if (~extnMRequest_instruction[12]) begin // @[core.scala 415:47]
        if (extnMRequest_instruction[3]) begin // @[core.scala 419:48]
          if (extnMRequest_rs2[31]) begin // @[core.scala 421:43]
            division_divisor <= _division_divisor_T_10; // @[core.scala 421:62]
          end else begin
            division_divisor <= _GEN_89;
          end
        end else begin
          division_divisor <= _GEN_89;
        end
      end else begin
        division_divisor <= _GEN_86;
      end
    end
    if (extnMRequest_valid & extnMRequest_instruction[14]) begin // @[core.scala 404:67]
      division_counter <= 7'h41; // @[core.scala 405:22]
    end else begin
      division_counter <= _division_counter_T_1; // @[core.scala 402:20]
    end
    if (reset) begin // @[core.scala 222:27]
      fwdBuffers_0_valid <= 1'h0; // @[core.scala 222:27]
    end else begin
      fwdBuffers_0_valid <= fwdFrom_0_valid; // @[core.scala 466:64]
    end
    fwdBuffers_0_prfDest <= singleCycleArithmeticRequest_prfDest; // @[core.scala 228:33 232:22]
    fwdBuffers_0_result <= arithmeticResult[63:0]; // @[core.scala 228:33 269:21]
    if (reset) begin // @[core.scala 222:27]
      fwdBuffers_1_valid <= 1'h0; // @[core.scala 222:27]
    end else begin
      fwdBuffers_1_valid <= fwdBuffers_0_valid; // @[core.scala 466:64]
    end
    fwdBuffers_1_prfDest <= fwdBuffers_0_prfDest; // @[core.scala 228:33 229:14]
    fwdBuffers_1_result <= fwdBuffers_0_result; // @[core.scala 228:33 229:14]
    narrowMuls_0 <= extnMRequest_rs1[31:0] * extnMRequest_rs2[31:0]; // @[core.scala 329:29]
    narrowMuls_1 <= extnMRequest_rs1[63:32] * extnMRequest_rs2[31:0]; // @[core.scala 330:30]
    narrowMuls_2 <= _T_39[63:0]; // @[core.scala 340:80]
    narrowMuls_3 <= extnMRequest_rs1[31:0] * extnMRequest_rs2[63:32]; // @[core.scala 332:29]
    narrowMuls_4 <= _T_40[63:0]; // @[core.scala 340:80]
    narrowMuls_5 <= extnMRequest_rs1[63:32] * extnMRequest_rs2[63:32]; // @[core.scala 334:30]
    narrowMuls_6 <= _T_41[63:0]; // @[core.scala 340:80]
    narrowMuls_7 <= $signed(_partialMuls32x32_T_30) * $signed(_partialMuls32x32_T_32); // @[core.scala 340:41]
    narrowMuls_8 <= $signed(_partialMuls32x32_T_34) * $signed(_partialMuls32x32_T_36); // @[core.scala 340:41]
    if (~mExtensionReady) begin // @[core.scala 388:26]
      if (branchEvals_valid & |_T_78) begin // @[core.scala 389:73]
        if (branchEvals_passed) begin // @[core.scala 390:30]
          divBranchMask <= _divBranchMask_T_5; // @[core.scala 391:23]
        end else begin
          divBranchMask <= _GEN_78;
        end
      end else begin
        divBranchMask <= _GEN_78;
      end
    end else begin
      divBranchMask <= _GEN_78;
    end
    if (reset) begin // @[core.scala 475:26]
      branchPCs_0_valid <= 1'h0; // @[core.scala 475:26]
    end else if (branchEvals_valid & _T) begin // @[core.scala 610:46]
      branchPCs_0_valid <= 1'h0; // @[core.scala 611:32]
    end else if (branchInstruction_valid) begin // @[core.scala 612:39]
      branchPCs_0_valid <= entry_1_valid; // @[core.scala 623:40]
    end else if (~branchPCs_0_valid) begin // @[core.scala 605:82]
      branchPCs_0_valid <= decode_branchPCs_branchPCReady; // @[core.scala 606:15]
    end
    if (branchEvals_valid & _T) begin // @[core.scala 610:46]
      branchPCs_0_pc <= _GEN_161;
    end else if (branchInstruction_valid) begin // @[core.scala 612:39]
      if (branchPCs_1_valid) begin // @[core.scala 617:22]
        branchPCs_0_pc <= branchPCs_1_pc;
      end else begin
        branchPCs_0_pc <= decode_branchPCs_branchPC;
      end
    end else begin
      branchPCs_0_pc <= _GEN_161;
    end
    if (branchEvals_valid & _T) begin // @[core.scala 610:46]
      branchPCs_0_branchMask <= _GEN_162;
    end else if (branchInstruction_valid) begin // @[core.scala 612:39]
      if (branchPCs_1_valid) begin // @[core.scala 618:30]
        branchPCs_0_branchMask <= branchPCs_1_branchMask;
      end else begin
        branchPCs_0_branchMask <= decode_branchPCs_branchMask;
      end
    end else begin
      branchPCs_0_branchMask <= _GEN_162;
    end
    if (reset) begin // @[core.scala 475:26]
      branchPCs_1_valid <= 1'h0; // @[core.scala 475:26]
    end else if (branchEvals_valid & _T) begin // @[core.scala 610:46]
      branchPCs_1_valid <= 1'h0; // @[core.scala 611:32]
    end else if (branchInstruction_valid) begin // @[core.scala 612:39]
      branchPCs_1_valid <= entry_2_valid; // @[core.scala 623:40]
    end else if (branchPCs_0_valid & ~branchPCs_1_valid) begin // @[core.scala 605:82]
      branchPCs_1_valid <= decode_branchPCs_branchPCReady; // @[core.scala 606:15]
    end
    if (branchEvals_valid & _T) begin // @[core.scala 610:46]
      branchPCs_1_pc <= _GEN_164;
    end else if (branchInstruction_valid) begin // @[core.scala 612:39]
      if (branchPCs_2_valid) begin // @[core.scala 617:22]
        branchPCs_1_pc <= branchPCs_2_pc;
      end else begin
        branchPCs_1_pc <= decode_branchPCs_branchPC;
      end
    end else begin
      branchPCs_1_pc <= _GEN_164;
    end
    if (branchEvals_valid & _T) begin // @[core.scala 610:46]
      branchPCs_1_branchMask <= _GEN_165;
    end else if (branchInstruction_valid) begin // @[core.scala 612:39]
      if (branchPCs_2_valid) begin // @[core.scala 618:30]
        branchPCs_1_branchMask <= branchPCs_2_branchMask;
      end else begin
        branchPCs_1_branchMask <= decode_branchPCs_branchMask;
      end
    end else begin
      branchPCs_1_branchMask <= _GEN_165;
    end
    if (reset) begin // @[core.scala 475:26]
      branchPCs_2_valid <= 1'h0; // @[core.scala 475:26]
    end else if (branchEvals_valid & _T) begin // @[core.scala 610:46]
      branchPCs_2_valid <= 1'h0; // @[core.scala 611:32]
    end else if (branchInstruction_valid) begin // @[core.scala 612:39]
      branchPCs_2_valid <= entry_3_valid; // @[core.scala 623:40]
    end else if (_T_133 & ~branchPCs_2_valid) begin // @[core.scala 605:82]
      branchPCs_2_valid <= decode_branchPCs_branchPCReady; // @[core.scala 606:15]
    end
    if (branchEvals_valid & _T) begin // @[core.scala 610:46]
      branchPCs_2_pc <= _GEN_167;
    end else if (branchInstruction_valid) begin // @[core.scala 612:39]
      if (branchPCs_3_valid) begin // @[core.scala 617:22]
        branchPCs_2_pc <= branchPCs_3_pc;
      end else begin
        branchPCs_2_pc <= decode_branchPCs_branchPC;
      end
    end else begin
      branchPCs_2_pc <= _GEN_167;
    end
    if (branchEvals_valid & _T) begin // @[core.scala 610:46]
      branchPCs_2_branchMask <= _GEN_168;
    end else if (branchInstruction_valid) begin // @[core.scala 612:39]
      if (branchPCs_3_valid) begin // @[core.scala 618:30]
        branchPCs_2_branchMask <= branchPCs_3_branchMask;
      end else begin
        branchPCs_2_branchMask <= decode_branchPCs_branchMask;
      end
    end else begin
      branchPCs_2_branchMask <= _GEN_168;
    end
    if (reset) begin // @[core.scala 475:26]
      branchPCs_3_valid <= 1'h0; // @[core.scala 475:26]
    end else if (branchEvals_valid & _T) begin // @[core.scala 610:46]
      branchPCs_3_valid <= 1'h0; // @[core.scala 611:32]
    end else if (branchInstruction_valid) begin // @[core.scala 612:39]
      branchPCs_3_valid <= 1'h0; // @[core.scala 624:41]
    end else if (_T_134 & ~branchPCs_3_valid) begin // @[core.scala 605:82]
      branchPCs_3_valid <= decode_branchPCs_branchPCReady; // @[core.scala 606:15]
    end
    if (_T_134 & ~branchPCs_3_valid) begin // @[core.scala 605:82]
      branchPCs_3_pc <= decode_branchPCs_branchPC; // @[core.scala 607:12]
    end
    if (_T_134 & ~branchPCs_3_valid) begin // @[core.scala 605:82]
      branchPCs_3_branchMask <= decode_branchPCs_branchMask; // @[core.scala 608:20]
    end
    if (reset) begin // @[core.scala 482:29]
      predictedPCs_0_valid <= 1'h0; // @[core.scala 482:29]
    end else if (_T_145) begin // @[core.scala 633:46]
      predictedPCs_0_valid <= 1'h0; // @[core.scala 634:35]
    end else if (branchInstruction_valid) begin // @[core.scala 635:39]
      predictedPCs_0_valid <= entry_5_valid; // @[core.scala 645:40]
    end else if (~predictedPCs_0_valid) begin // @[core.scala 629:82]
      predictedPCs_0_valid <= decode_branchPCs_predictedPCReady; // @[core.scala 630:15]
    end
    if (_T_145) begin // @[core.scala 633:46]
      predictedPCs_0_pc <= _GEN_193;
    end else if (branchInstruction_valid) begin // @[core.scala 635:39]
      if (predictedPCs_1_valid) begin // @[core.scala 640:22]
        predictedPCs_0_pc <= predictedPCs_1_pc;
      end else begin
        predictedPCs_0_pc <= decode_branchPCs_predictedPC;
      end
    end else begin
      predictedPCs_0_pc <= _GEN_193;
    end
    if (reset) begin // @[core.scala 482:29]
      predictedPCs_1_valid <= 1'h0; // @[core.scala 482:29]
    end else if (_T_145) begin // @[core.scala 633:46]
      predictedPCs_1_valid <= 1'h0; // @[core.scala 634:35]
    end else if (branchInstruction_valid) begin // @[core.scala 635:39]
      predictedPCs_1_valid <= entry_6_valid; // @[core.scala 645:40]
    end else if (predictedPCs_0_valid & ~predictedPCs_1_valid) begin // @[core.scala 629:82]
      predictedPCs_1_valid <= decode_branchPCs_predictedPCReady; // @[core.scala 630:15]
    end
    if (_T_145) begin // @[core.scala 633:46]
      predictedPCs_1_pc <= _GEN_195;
    end else if (branchInstruction_valid) begin // @[core.scala 635:39]
      if (predictedPCs_2_valid) begin // @[core.scala 640:22]
        predictedPCs_1_pc <= predictedPCs_2_pc;
      end else begin
        predictedPCs_1_pc <= decode_branchPCs_predictedPC;
      end
    end else begin
      predictedPCs_1_pc <= _GEN_195;
    end
    if (reset) begin // @[core.scala 482:29]
      predictedPCs_2_valid <= 1'h0; // @[core.scala 482:29]
    end else if (_T_145) begin // @[core.scala 633:46]
      predictedPCs_2_valid <= 1'h0; // @[core.scala 634:35]
    end else if (branchInstruction_valid) begin // @[core.scala 635:39]
      predictedPCs_2_valid <= entry_7_valid; // @[core.scala 645:40]
    end else if (_T_151 & ~predictedPCs_2_valid) begin // @[core.scala 629:82]
      predictedPCs_2_valid <= decode_branchPCs_predictedPCReady; // @[core.scala 630:15]
    end
    if (_T_145) begin // @[core.scala 633:46]
      predictedPCs_2_pc <= _GEN_197;
    end else if (branchInstruction_valid) begin // @[core.scala 635:39]
      if (predictedPCs_3_valid) begin // @[core.scala 640:22]
        predictedPCs_2_pc <= predictedPCs_3_pc;
      end else begin
        predictedPCs_2_pc <= decode_branchPCs_predictedPC;
      end
    end else begin
      predictedPCs_2_pc <= _GEN_197;
    end
    if (reset) begin // @[core.scala 482:29]
      predictedPCs_3_valid <= 1'h0; // @[core.scala 482:29]
    end else if (_T_145) begin // @[core.scala 633:46]
      predictedPCs_3_valid <= 1'h0; // @[core.scala 634:35]
    end else if (branchInstruction_valid) begin // @[core.scala 635:39]
      predictedPCs_3_valid <= 1'h0; // @[core.scala 646:44]
    end else if (_T_152 & ~predictedPCs_3_valid) begin // @[core.scala 629:82]
      predictedPCs_3_valid <= decode_branchPCs_predictedPCReady; // @[core.scala 630:15]
    end
    if (_T_152 & ~predictedPCs_3_valid) begin // @[core.scala 629:82]
      predictedPCs_3_pc <= decode_branchPCs_predictedPC; // @[core.scala 631:12]
    end
    if (reset) begin // @[core.scala 487:34]
      branchInstruction_valid <= 1'h0; // @[core.scala 487:34]
    end else if (branchEvals_valid) begin // @[core.scala 533:25]
      if (_T & |_T_128) begin // @[core.scala 537:83]
        branchInstruction_valid <= 1'h0; // @[core.scala 538:31]
      end else begin
        branchInstruction_valid <= prf_toExec_valid & prf_toExec_instruction[6:4] == 3'h6; // @[core.scala 520:27]
      end
    end else begin
      branchInstruction_valid <= prf_toExec_valid & prf_toExec_instruction[6:4] == 3'h6; // @[core.scala 520:27]
    end
    if (prf_toExec_valid & prf_toExec_instruction[6:5] == 2'h3) begin // @[core.scala 521:71]
      if (_addressGenerationInput_rs1_T_3) begin // @[Mux.scala 101:16]
        branchInstruction_rs1 <= fwdFrom_0_result;
      end else if (_addressGenerationInput_rs1_T_5) begin // @[Mux.scala 101:16]
        branchInstruction_rs1 <= fwdBuffers_0_result;
      end else if (_addressGenerationInput_rs1_T_7) begin // @[Mux.scala 101:16]
        branchInstruction_rs1 <= fwdBuffers_1_result;
      end else begin
        branchInstruction_rs1 <= prf_toExec_rs1Data;
      end
    end
    if (prf_toExec_valid & prf_toExec_instruction[6:5] == 2'h3) begin // @[core.scala 521:71]
      if (_singleCycleArithmeticRequest_rs2_T_5) begin // @[Mux.scala 101:16]
        branchInstruction_rs2 <= fwdFrom_0_result;
      end else if (_singleCycleArithmeticRequest_rs2_T_7) begin // @[Mux.scala 101:16]
        branchInstruction_rs2 <= fwdBuffers_0_result;
      end else if (_singleCycleArithmeticRequest_rs2_T_9) begin // @[Mux.scala 101:16]
        branchInstruction_rs2 <= fwdBuffers_1_result;
      end else begin
        branchInstruction_rs2 <= prf_toExec_rs2Data;
      end
    end
    branchInstruction_robAddr <= _GEN_140[3:0];
    if (prf_toExec_valid & prf_toExec_instruction[6:5] == 2'h3) begin // @[core.scala 521:71]
      branchInstruction_instruction <= prf_toExec_instruction; // @[core.scala 530:35]
    end
    if (2'h3 == prf_toExec_instruction[3:2]) begin // @[core.scala 498:31]
      branchInstruction_immediate <= _branchInstruction_immediate_T_18; // @[core.scala 498:31]
    end else if (2'h2 == prf_toExec_instruction[3:2]) begin // @[core.scala 498:31]
      branchInstruction_immediate <= 64'h0; // @[core.scala 498:31]
    end else if (2'h1 == prf_toExec_instruction[3:2]) begin // @[core.scala 498:31]
      branchInstruction_immediate <= arithmeticImm; // @[core.scala 498:31]
    end else begin
      branchInstruction_immediate <= _branchInstruction_immediate_T_6;
    end
    branchEvals_robAddr <= branchInstruction_robAddr; // @[core.scala 543:23]
    if (2'h3 == branchInstruction_instruction[3:2]) begin // @[core.scala 596:22]
      branchEvals_nextPC <= _nextCorrectPC_T_2; // @[core.scala 596:22]
    end else if (2'h2 == branchInstruction_instruction[3:2]) begin // @[core.scala 596:22]
      branchEvals_nextPC <= 64'h0; // @[core.scala 596:22]
    end else if (2'h1 == branchInstruction_instruction[3:2]) begin // @[core.scala 596:22]
      branchEvals_nextPC <= _nextCorrectPC_T_7; // @[core.scala 596:22]
    end else if (_GEN_155) begin // @[core.scala 590:10]
      branchEvals_nextPC <= _nextCorrectPC_T_2;
    end else begin
      branchEvals_nextPC <= _nextCorrectPC_T_4;
    end
    if (3'h7 == branchInstruction_instruction[14:12]) begin // @[core.scala 676:41]
      fetch_branchRes_branchTaken_REG <= branchTaken_conditionEval_7; // @[core.scala 676:41]
    end else if (3'h6 == branchInstruction_instruction[14:12]) begin // @[core.scala 676:41]
      fetch_branchRes_branchTaken_REG <= branchTaken_conditionEval_6; // @[core.scala 676:41]
    end else if (3'h5 == branchInstruction_instruction[14:12]) begin // @[core.scala 676:41]
      fetch_branchRes_branchTaken_REG <= branchTaken_conditionEval_5; // @[core.scala 676:41]
    end else if (3'h4 == branchInstruction_instruction[14:12]) begin // @[core.scala 676:41]
      fetch_branchRes_branchTaken_REG <= branchTaken_conditionEval_4; // @[core.scala 676:41]
    end else begin
      fetch_branchRes_branchTaken_REG <= _GEN_217;
    end
    fetch_branchRes_pc_REG <= branchPCs_0_pc; // @[core.scala 678:32]
    rob_execPorts_0_mtval_REG <= singleCycleArithmeticRequest_rs1; // @[core.scala 712:36]
    if (reset) begin // @[core.scala 733:129]
      REG <= 1'h0; // @[core.scala 733:129]
    end else begin
      REG <= _fwdFrom_0_valid_T_1 & singleCycleArithmeticRequest_instruction[6:2] != 5'h1c; // @[core.scala 733:129]
    end
    prf_fromStore_rs2Addr_REG <= dataQueue_toPRF_rs2Addr; // @[core.scala 769:43]
    prf_fromStore_rs2Addr_REG_1 <= prf_fromStore_rs2Addr_REG; // @[core.scala 769:35]
    if (reset) begin // @[core.scala 770:41]
      prf_fromStore_valid_REG <= 1'h0; // @[core.scala 770:41]
    end else begin
      prf_fromStore_valid_REG <= dataQueue_toPRF_valid & dataQueue_fromROB_readyNow; // @[core.scala 770:41]
    end
    if (reset) begin // @[core.scala 770:33]
      prf_fromStore_valid_REG_1 <= 1'h0; // @[core.scala 770:33]
    end else begin
      prf_fromStore_valid_REG_1 <= prf_fromStore_valid_REG; // @[core.scala 770:33]
    end
    if (reset) begin // @[core.scala 816:27]
      fenceState_state <= 2'h0; // @[core.scala 816:27]
    end else if (2'h0 == fenceState_state) begin // @[core.scala 823:28]
      if (fetch_toDecode_fired & _T_188 == 20'hf) begin // @[core.scala 825:115]
        fenceState_state <= 2'h1; // @[core.scala 826:26]
      end
    end else if (2'h1 == fenceState_state) begin // @[core.scala 823:28]
      if (_T_145) begin // @[core.scala 830:54]
        fenceState_state <= 2'h0; // @[core.scala 833:26]
      end else begin
        fenceState_state <= _GEN_223;
      end
    end else if (2'h2 == fenceState_state) begin // @[core.scala 823:28]
      fenceState_state <= _GEN_233;
    end
    if (!(2'h0 == fenceState_state)) begin // @[core.scala 823:28]
      if (2'h1 == fenceState_state) begin // @[core.scala 823:28]
        if (!(_T_145)) begin // @[core.scala 830:54]
          if (decode_toExec_fired & _T_195 == 20'hf) begin // @[core.scala 834:119]
            fenceState_branchMask <= decode_toExec_branchMask; // @[core.scala 836:31]
          end
        end
      end else if (2'h2 == fenceState_state) begin // @[core.scala 823:28]
        if (!(branchEvals_valid & |_T_199 & _T)) begin // @[core.scala 840:110]
          fenceState_branchMask <= _GEN_231;
        end
      end
    end
    REG_1 <= _T_145 & (fetch_toDecode_instruction == 32'hff0000f & fetch_toDecode_fired); // @[core.scala 874:53]
    branchCounter <= _GEN_249[2:0]; // @[core.scala 987:{30,30}]
    if (branchEvals_valid) begin // @[core.scala 1003:27]
      lastBranchExecRob <= branchEvals_robAddr; // @[core.scala 1004:23]
    end
    if (branchEvals_valid) begin // @[core.scala 1003:27]
      lastBranchExecPC <= lastBranchExecPC_REG; // @[core.scala 1005:22]
    end
    lastBranchExecPC_REG <= branchPCs_0_pc; // @[core.scala 1005:32]
    if (reset) begin // @[core.scala 1021:34]
      lastRetiredSystem <= 1'h0; // @[core.scala 1021:34]
    end else if (decode_fromFetch_fired) begin // @[core.scala 1022:32]
      lastRetiredSystem <= fetch_toDecode_instruction[6:0] == 7'h73; // @[core.scala 1022:52]
    end
    if (reset) begin // @[core.scala 1024:38]
      interruptInjectStatus <= 2'h0; // @[core.scala 1024:38]
    end else if (2'h0 == interruptInjectStatus) begin // @[core.scala 1025:33]
      if (decode_canTakeInterrupt & MTIP & ~lastRetiredSystem) begin // @[core.scala 1029:67]
        interruptInjectStatus <= 2'h1; // @[core.scala 1029:91]
      end
    end else if (2'h1 == interruptInjectStatus) begin // @[core.scala 1025:33]
      if (decode_canTakeInterrupt) begin // @[core.scala 1033:56]
        interruptInjectStatus <= _GEN_280;
      end
    end else if (2'h2 == interruptInjectStatus) begin // @[core.scala 1025:33]
      interruptInjectStatus <= 2'h3; // @[core.scala 1057:29]
    end else begin
      interruptInjectStatus <= _GEN_290;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  branchEvals_branchMask = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  branchEvals_passed = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  branchEvals_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  extnMResponse_prfDest = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  extnMResponse_valid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  extnResponseInstruction = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  mExtensionReady = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  addressGenerationInput_valid = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  addressGenerationInput_rs1 = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  addressGenerationInput_instruction = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  addressGenerationInput_prfDest = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  addressGenerationInput_robAddr = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  addressGenerationInput_branchMask = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  memoryRequest_valid = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  memoryRequest_address = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  memoryRequest_instruction = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  memoryRequest_branchMask = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  memoryRequest_robAddr = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  memoryRequest_prfDest = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  singleCycleArithmeticRequest_valid = _RAND_19[0:0];
  _RAND_20 = {2{`RANDOM}};
  singleCycleArithmeticRequest_rs1 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  singleCycleArithmeticRequest_rs2 = _RAND_21[63:0];
  _RAND_22 = {1{`RANDOM}};
  singleCycleArithmeticRequest_instruction = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  singleCycleArithmeticRequest_prfDest = _RAND_23[5:0];
  _RAND_24 = {1{`RANDOM}};
  singleCycleArithmeticRequest_robAddr = _RAND_24[3:0];
  _RAND_25 = {1{`RANDOM}};
  singleCycleArithmeticRequest_branchMask = _RAND_25[3:0];
  _RAND_26 = {1{`RANDOM}};
  singleCycleArithmeticResponse_valid = _RAND_26[0:0];
  _RAND_27 = {2{`RANDOM}};
  singleCycleArithmeticResponse_result = _RAND_27[63:0];
  _RAND_28 = {1{`RANDOM}};
  singleCycleArithmeticResponse_prfDest = _RAND_28[5:0];
  _RAND_29 = {1{`RANDOM}};
  singleCycleArithmeticResponse_robAddr = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  extnMRequest_valid = _RAND_30[0:0];
  _RAND_31 = {2{`RANDOM}};
  extnMRequest_rs1 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  extnMRequest_rs2 = _RAND_32[63:0];
  _RAND_33 = {1{`RANDOM}};
  extnMRequest_instruction = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  extnMRequest_prfDest = _RAND_34[5:0];
  _RAND_35 = {1{`RANDOM}};
  extnMRequest_robAddr = _RAND_35[3:0];
  _RAND_36 = {1{`RANDOM}};
  extnMRequest_branchMask = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  extnMServicing_valid = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  extnMServicing_instruction = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  extnMServicing_prfDest = _RAND_39[5:0];
  _RAND_40 = {1{`RANDOM}};
  extnMServicing_robAddr = _RAND_40[3:0];
  _RAND_41 = {1{`RANDOM}};
  extnMServicing_branchMask = _RAND_41[3:0];
  _RAND_42 = {1{`RANDOM}};
  extnMPartialServicing_valid = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  extnMPartialServicing_instruction = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  extnMPartialServicing_prfDest = _RAND_44[5:0];
  _RAND_45 = {1{`RANDOM}};
  extnMPartialServicing_robAddr = _RAND_45[3:0];
  _RAND_46 = {1{`RANDOM}};
  extnMPartialServicing_branchMask = _RAND_46[3:0];
  _RAND_47 = {3{`RANDOM}};
  muls_0 = _RAND_47[95:0];
  _RAND_48 = {3{`RANDOM}};
  muls_1 = _RAND_48[95:0];
  _RAND_49 = {3{`RANDOM}};
  muls_2 = _RAND_49[95:0];
  _RAND_50 = {3{`RANDOM}};
  muls_3 = _RAND_50[95:0];
  _RAND_51 = {3{`RANDOM}};
  muls_4 = _RAND_51[95:0];
  _RAND_52 = {3{`RANDOM}};
  muls_5 = _RAND_52[95:0];
  _RAND_53 = {2{`RANDOM}};
  extnMResponse_result = _RAND_53[63:0];
  _RAND_54 = {1{`RANDOM}};
  extnMResponse_robAddr = _RAND_54[3:0];
  _RAND_55 = {1{`RANDOM}};
  division_request_valid = _RAND_55[0:0];
  _RAND_56 = {2{`RANDOM}};
  division_request_rs1 = _RAND_56[63:0];
  _RAND_57 = {2{`RANDOM}};
  division_request_rs2 = _RAND_57[63:0];
  _RAND_58 = {1{`RANDOM}};
  division_request_instruction = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  division_request_prfDest = _RAND_59[5:0];
  _RAND_60 = {1{`RANDOM}};
  division_request_robAddr = _RAND_60[3:0];
  _RAND_61 = {1{`RANDOM}};
  division_request_branchMask = _RAND_61[3:0];
  _RAND_62 = {3{`RANDOM}};
  division_quotient = _RAND_62[64:0];
  _RAND_63 = {3{`RANDOM}};
  division_remainder = _RAND_63[64:0];
  _RAND_64 = {3{`RANDOM}};
  division_divisor = _RAND_64[64:0];
  _RAND_65 = {1{`RANDOM}};
  division_counter = _RAND_65[6:0];
  _RAND_66 = {1{`RANDOM}};
  fwdBuffers_0_valid = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  fwdBuffers_0_prfDest = _RAND_67[5:0];
  _RAND_68 = {2{`RANDOM}};
  fwdBuffers_0_result = _RAND_68[63:0];
  _RAND_69 = {1{`RANDOM}};
  fwdBuffers_1_valid = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  fwdBuffers_1_prfDest = _RAND_70[5:0];
  _RAND_71 = {2{`RANDOM}};
  fwdBuffers_1_result = _RAND_71[63:0];
  _RAND_72 = {2{`RANDOM}};
  narrowMuls_0 = _RAND_72[63:0];
  _RAND_73 = {2{`RANDOM}};
  narrowMuls_1 = _RAND_73[63:0];
  _RAND_74 = {2{`RANDOM}};
  narrowMuls_2 = _RAND_74[63:0];
  _RAND_75 = {2{`RANDOM}};
  narrowMuls_3 = _RAND_75[63:0];
  _RAND_76 = {2{`RANDOM}};
  narrowMuls_4 = _RAND_76[63:0];
  _RAND_77 = {2{`RANDOM}};
  narrowMuls_5 = _RAND_77[63:0];
  _RAND_78 = {2{`RANDOM}};
  narrowMuls_6 = _RAND_78[63:0];
  _RAND_79 = {2{`RANDOM}};
  narrowMuls_7 = _RAND_79[63:0];
  _RAND_80 = {2{`RANDOM}};
  narrowMuls_8 = _RAND_80[63:0];
  _RAND_81 = {1{`RANDOM}};
  divBranchMask = _RAND_81[3:0];
  _RAND_82 = {1{`RANDOM}};
  branchPCs_0_valid = _RAND_82[0:0];
  _RAND_83 = {2{`RANDOM}};
  branchPCs_0_pc = _RAND_83[63:0];
  _RAND_84 = {1{`RANDOM}};
  branchPCs_0_branchMask = _RAND_84[3:0];
  _RAND_85 = {1{`RANDOM}};
  branchPCs_1_valid = _RAND_85[0:0];
  _RAND_86 = {2{`RANDOM}};
  branchPCs_1_pc = _RAND_86[63:0];
  _RAND_87 = {1{`RANDOM}};
  branchPCs_1_branchMask = _RAND_87[3:0];
  _RAND_88 = {1{`RANDOM}};
  branchPCs_2_valid = _RAND_88[0:0];
  _RAND_89 = {2{`RANDOM}};
  branchPCs_2_pc = _RAND_89[63:0];
  _RAND_90 = {1{`RANDOM}};
  branchPCs_2_branchMask = _RAND_90[3:0];
  _RAND_91 = {1{`RANDOM}};
  branchPCs_3_valid = _RAND_91[0:0];
  _RAND_92 = {2{`RANDOM}};
  branchPCs_3_pc = _RAND_92[63:0];
  _RAND_93 = {1{`RANDOM}};
  branchPCs_3_branchMask = _RAND_93[3:0];
  _RAND_94 = {1{`RANDOM}};
  predictedPCs_0_valid = _RAND_94[0:0];
  _RAND_95 = {2{`RANDOM}};
  predictedPCs_0_pc = _RAND_95[63:0];
  _RAND_96 = {1{`RANDOM}};
  predictedPCs_1_valid = _RAND_96[0:0];
  _RAND_97 = {2{`RANDOM}};
  predictedPCs_1_pc = _RAND_97[63:0];
  _RAND_98 = {1{`RANDOM}};
  predictedPCs_2_valid = _RAND_98[0:0];
  _RAND_99 = {2{`RANDOM}};
  predictedPCs_2_pc = _RAND_99[63:0];
  _RAND_100 = {1{`RANDOM}};
  predictedPCs_3_valid = _RAND_100[0:0];
  _RAND_101 = {2{`RANDOM}};
  predictedPCs_3_pc = _RAND_101[63:0];
  _RAND_102 = {1{`RANDOM}};
  branchInstruction_valid = _RAND_102[0:0];
  _RAND_103 = {2{`RANDOM}};
  branchInstruction_rs1 = _RAND_103[63:0];
  _RAND_104 = {2{`RANDOM}};
  branchInstruction_rs2 = _RAND_104[63:0];
  _RAND_105 = {1{`RANDOM}};
  branchInstruction_robAddr = _RAND_105[3:0];
  _RAND_106 = {1{`RANDOM}};
  branchInstruction_instruction = _RAND_106[31:0];
  _RAND_107 = {2{`RANDOM}};
  branchInstruction_immediate = _RAND_107[63:0];
  _RAND_108 = {1{`RANDOM}};
  branchEvals_robAddr = _RAND_108[3:0];
  _RAND_109 = {2{`RANDOM}};
  branchEvals_nextPC = _RAND_109[63:0];
  _RAND_110 = {1{`RANDOM}};
  fetch_branchRes_branchTaken_REG = _RAND_110[0:0];
  _RAND_111 = {2{`RANDOM}};
  fetch_branchRes_pc_REG = _RAND_111[63:0];
  _RAND_112 = {2{`RANDOM}};
  rob_execPorts_0_mtval_REG = _RAND_112[63:0];
  _RAND_113 = {1{`RANDOM}};
  REG = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  prf_fromStore_rs2Addr_REG = _RAND_114[5:0];
  _RAND_115 = {1{`RANDOM}};
  prf_fromStore_rs2Addr_REG_1 = _RAND_115[5:0];
  _RAND_116 = {1{`RANDOM}};
  prf_fromStore_valid_REG = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  prf_fromStore_valid_REG_1 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  fenceState_state = _RAND_118[1:0];
  _RAND_119 = {1{`RANDOM}};
  fenceState_branchMask = _RAND_119[3:0];
  _RAND_120 = {1{`RANDOM}};
  REG_1 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  branchCounter = _RAND_121[2:0];
  _RAND_122 = {1{`RANDOM}};
  lastBranchExecRob = _RAND_122[3:0];
  _RAND_123 = {2{`RANDOM}};
  lastBranchExecPC = _RAND_123[63:0];
  _RAND_124 = {2{`RANDOM}};
  lastBranchExecPC_REG = _RAND_124[63:0];
  _RAND_125 = {1{`RANDOM}};
  lastRetiredSystem = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  interruptInjectStatus = _RAND_126[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
